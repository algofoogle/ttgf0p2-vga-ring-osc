* NGSPICE file created from tt_um_algofoogle_vgaringosc_parax.ext - technology: gf180mcuD

.subckt tt_um_algofoogle_vgaringosc_parax VGND VPWR clk ena rst_n ui_in[0] ui_in[1]
+ ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2]
+ uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2]
+ uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2]
+ uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2]
+ uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
X0 VPWR.t1209 a_66204_5863# a_66116_5960# VPWR.t1208 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_33948_16839# a_33860_16936# VGND.t1133 VGND.t1132 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 VPWR.t319 a_42236_2727# a_42148_2824# VPWR.t318 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3 VPWR.t236 a_44296_24393.t14 clkbuf_1_0__f_clk.I.t15 VPWR.t235 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4 a_43600_22504# _304_.ZN.t10 VGND.t235 VGND.t234 nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VPWR.t321 a_9635_30644# uio_oe[5].t0 VPWR.t320 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6 a_35224_23705# a_33376_23659# a_34939_23705# VPWR.t1913 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X7 VPWR.t552 a_59484_9432# a_59396_9476# VPWR.t551 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X8 VPWR.t5245 a_66204_2727# a_66116_2824# VPWR.t5244 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X9 a_44812_19369# _325_.ZN a_43888_19204# VGND.t326 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X10 a_55228_20408# a_55140_20452# VGND.t5390 VGND.t5389 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X11 a_2364_27815# a_2276_27912# VGND.t5767 VGND.t4204 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X12 _332_.Z a_40244_18180# VPWR.t899 VPWR.t898 pfet_06v0 ad=0.5346p pd=3.31u as=0.4268p ps=2.175u w=1.215u l=0.5u
X13 _324_.C.t7 a_65072_29860# VGND.t1063 VGND.t1059 nfet_06v0 ad=0.1183p pd=0.975u as=0.23432p ps=1.94u w=0.455u l=0.6u
X14 VPWR.t1018 a_41564_1592# a_41476_1636# VPWR.t1017 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 VPWR.t351 a_3260_30951# a_3172_31048# VPWR.t350 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X16 VPWR.t5161 _473_.Q a_47860_21640# VPWR.t5160 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X17 a_28054_30196# _359_.B.t2 VGND.t6465 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.2911p ps=1.53u w=0.82u l=0.6u
X18 a_27328_25227# a_26916_25640.t2 VPWR.t6740 VPWR.t6739 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X19 uo_out[6].t11 _287_.A1.t8 VGND.t6478 VGND.t6477 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X20 VPWR.t840 a_65532_1592# a_65444_1636# VPWR.t839 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X21 VPWR.t1100 a_16028_1592# a_15940_1636# VPWR.t1099 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X22 _416_.ZN _416_.A2 VGND.t6026 VGND.t6025 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X23 VPWR.t6734 _268_.A1.t2 a_53212_29816# VPWR.t6733 pfet_06v0 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X24 a_66540_19975# a_66452_20072# VGND.t876 VGND.t875 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X25 VPWR.t6743 _474_.CLK.t32 a_48384_26724# VPWR.t6742 pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X26 a_15244_28248# a_15156_28292# VGND.t1380 VGND.t1379 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X27 VPWR.t976 a_47164_13703# a_47076_13800# VPWR.t975 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X28 a_48529_22460# _473_.Q VGND.t4998 VGND.t4997 nfet_06v0 ad=93.59999f pd=0.88u as=0.2288p ps=1.58u w=0.36u l=0.6u
X29 a_1916_2727# a_1828_2824# VGND.t4702 VGND.t1224 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X30 VPWR.t364 a_48956_18407# a_48868_18504# VPWR.t363 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X31 a_55340_19975# a_55252_20072# VGND.t773 VGND.t772 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X32 a_63516_19975# a_63428_20072# VGND.t2843 VGND.t2842 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X33 VPWR.t3638 _346_.A2 a_21268_27912# VPWR.t3637 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X34 a_48956_2727# a_48868_2824# VGND.t1355 VGND.t1354 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X35 a_49764_26724# _402_.A1.t4 VGND.t6427 VGND.t6426 nfet_06v0 ad=0.14p pd=1.1u as=0.104p ps=0.92u w=0.4u l=0.6u
X36 _421_.A1 _324_.B.t20 VPWR.t6707 VPWR.t6706 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X37 VGND.t951 _435_.A3 _435_.ZN VGND.t950 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X38 a_1020_24679# a_932_24776# VGND.t767 VGND.t766 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X39 VGND.t828 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN VGND.t827 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X40 a_48308_23588# _279_.Z a_49764_23588# VPWR.t5589 pfet_06v0 ad=0.5016p pd=3.16u as=0.3534p ps=1.76u w=1.14u l=0.5u
X41 VPWR.t905 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN VPWR.t904 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X42 a_44252_30951# a_44164_31048# VGND.t1385 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X43 a_2812_29383# a_2724_29480# VGND.t459 VGND.t458 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X44 VGND.t5051 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN VGND.t5050 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X45 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I VPWR.t1127 VPWR.t1126 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X46 VPWR.t1433 a_67996_2727# a_67908_2824# VPWR.t1432 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X47 VPWR.t5045 a_59372_14136# a_59284_14180# VPWR.t4307 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X48 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN VPWR.t3000 VPWR.t2999 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X49 VGND.t1191 _399_.ZN a_50940_24072# VGND.t1190 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X50 VPWR.t2996 a_49628_15704# a_49540_15748# VPWR.t2995 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X51 a_1020_21543# a_932_21640# VGND.t4976 VGND.t3839 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X52 VPWR.t313 a_62732_16839# a_62644_16936# VPWR.t312 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X53 VGND.t6479 _287_.A1.t9 uo_out[2].t7 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X54 a_67100_9432# a_67012_9476# VGND.t4475 VGND.t4474 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X55 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I VPWR.t6005 VPWR.t6004 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X56 a_66428_14136# a_66340_14180# VGND.t5024 VGND.t5023 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X57 VPWR.t5979 a_56348_14136# a_56260_14180# VPWR.t5978 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X58 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I VGND.t4975 VGND.t4974 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X59 VGND.t5786 a_35008_22461# a_34960_22505# VGND.t5785 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X60 VPWR.t3639 a_1020_6296# a_932_6340# VPWR.t2610 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X61 VGND.t1078 _237_.A1 a_60401_30300# VGND.t1077 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X62 a_67100_6296# a_67012_6340# VGND.t1117 VGND.t1116 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X63 a_41048_29816.t3 vgaringosc.workerclkbuff_notouch_.I.t4 VPWR.t6699 VPWR.t6698 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X64 a_66428_11000# a_66340_11044# VGND.t1357 VGND.t1356 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X65 VPWR.t5995 a_56348_11000# a_56260_11044# VPWR.t5994 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X66 VPWR.t1460 a_1468_4295# a_1380_4392# VPWR.t1459 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X67 a_32476_29167# _461_.D a_32308_29167# VGND.t835 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X68 VGND.t6382 _355_.C.t4 _346_.B VGND.t6381 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X69 VPWR.t4287 a_1020_3160# a_932_3204# VPWR.t3076 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X70 VPWR.t1392 a_47612_12135# a_47524_12232# VPWR.t1391 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X71 _252_.ZN _251_.ZN VGND.t1115 VGND.t1114 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X72 VGND.t5728 a_52415_31220# a_52891_30644# VGND.t45 nfet_06v0 ad=0.28262p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X73 VPWR.t1470 a_1468_1159# a_1380_1256# VPWR.t1364 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X74 VPWR.t894 a_16588_21543# a_16500_21640# VPWR.t893 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X75 a_39985_24372# _260_.A2 a_39781_24372# VGND.t6024 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X76 a_45148_2727# a_45060_2824# VGND.t3518 VGND.t3517 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X77 VPWR.t1164 a_35292_30951# a_35204_31048# VPWR.t1163 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X78 VPWR.t5145 _337_.ZN a_31964_28292# VPWR.t5144 pfet_06v0 ad=0.3766p pd=1.815u as=0.4599p ps=1.935u w=1.095u l=0.5u
X79 a_43192_25640# _284_.B a_42168_25640.t8 VGND.t5394 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X80 a_49628_9432# a_49540_9476# VGND.t500 VGND.t499 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X81 VPWR.t984 a_62172_17272# a_62084_17316# VPWR.t983 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X82 VGND.t6344 _230_.I.t2 a_60059_28776# VGND.t6343 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X83 VPWR.t1600 a_19948_27815# a_19860_27912# VPWR.t1599 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X84 VPWR.t846 a_64188_2727# a_64100_2824# VPWR.t845 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X85 a_43192_22504# _302_.Z a_42168_22504# VGND.t4847 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X86 a_65308_15704# a_65220_15748# VGND.t4141 VGND.t4140 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X87 a_37386_31048# _350_.A1.t2 _296_.ZN VPWR.t6621 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X88 VGND.t6354 _452_.CLK.t32 a_36548_27591.t1 VGND.t6353 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X89 VGND.t1106 _373_.A2 _373_.ZN VGND.t1105 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X90 VPWR.t787 a_50412_18407# a_50324_18504# VPWR.t786 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X91 a_55452_21543# a_55364_21640# VGND.t5987 VGND.t5986 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X92 a_33500_17272# a_33412_17316# VGND.t977 VGND.t976 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X93 a_50940_24072# _324_.C.t8 _424_.B1.t4 VGND.t6497 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X94 a_38529_22804# _304_.A1.t2 a_38325_22804# VGND.t6314 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X95 VPWR.t1594 a_20956_24679# a_20868_24776# VPWR.t1593 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X96 a_57020_23111# a_56932_23208# VGND.t5509 VGND.t5508 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X97 a_41048_29816.t6 vgaringosc.workerclkbuff_notouch_.I.t5 VGND.t6410 VGND.t6409 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X98 a_54864_22461.t0 _474_.CLK.t33 VPWR.t6745 VPWR.t6744 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X99 VPWR.t503 a_53996_25112# a_53908_25156# VPWR.t502 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X100 a_43254_21236# a_42778_21812# a_42982_21730# VGND.t4895 nfet_06v0 ad=43.2f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X101 VGND.t5388 _279_.Z _399_.A2 VGND.t5387 nfet_06v0 ad=0.2266p pd=1.91u as=0.1339p ps=1.035u w=0.515u l=0.6u
X102 _300_.ZN _447_.Q.t2 a_39333_20936# VGND.t6300 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X103 VPWR.t5635 a_4828_30951# a_4740_31048# VPWR.t5634 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X104 a_22344_26399# a_20496_26344# a_22059_26399# VPWR.t4818 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X105 a_2364_7864# a_2276_7908# VGND.t608 VGND.t607 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X106 a_45372_13703# a_45284_13800# VGND.t614 VGND.t613 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X107 a_37888_27555# a_37516_27599# VPWR.t911 VPWR.t910 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X108 VPWR.t961 _300_.A2 a_38576_22504# VPWR.t960 pfet_06v0 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X109 a_52884_18884# _424_.A1 _424_.ZN VPWR.t305 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X110 a_12444_29383# a_12356_29480# VGND.t4107 VGND.t4106 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X111 _350_.A2.t7 _337_.ZN a_30388_28776# VGND.t4980 nfet_06v0 ad=0.30965p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X112 a_2364_4728# a_2276_4772# VGND.t449 VGND.t448 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X113 a_66316_12135# a_66228_12232# VGND.t1175 VGND.t1174 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X114 VPWR.t3755 _267_.A2 _258_.I VPWR.t3754 pfet_06v0 ad=0.2561p pd=1.505u as=0.44325p ps=2.87u w=0.985u l=0.5u
X115 VGND.t306 _424_.A1 a_51240_20452# VGND.t305 nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X116 VPWR.t2498 a_59260_23111# a_59172_23208# VPWR.t2497 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X117 a_56516_26344# a_55956_25940# a_56388_25940# VGND.t2374 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X118 a_18380_23544# a_18292_23588# VGND.t3390 VGND.t3389 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X119 a_55116_12135# a_55028_12232# VGND.t4892 VGND.t4891 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X120 VPWR.t1115 a_30812_1159# a_30724_1256# VPWR.t1114 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X121 VGND.t1256 _397_.A4 a_46171_27508# VGND.t1255 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X122 VPWR.t6543 a_48272_25156.t14 _474_.CLK.t0 VPWR.t6542 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X123 VGND.t2870 a_48384_26724# clkload0.Z VGND.t2869 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X124 a_65756_4295# a_65668_4392# VGND.t465 VGND.t464 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X125 a_60276_29032# _252_.ZN VGND.t6009 VGND.t6008 nfet_06v0 ad=0.14p pd=1.1u as=0.224p ps=1.52u w=0.4u l=0.6u
X126 VPWR.t331 a_23532_23544# a_23444_23588# VPWR.t330 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X127 a_38340_21327# _301_.A1 VPWR.t3352 VPWR.t3351 pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X128 a_35140_26680# _362_.B.t4 VPWR.t6526 VPWR.t6525 pfet_06v0 ad=0.2354p pd=1.95u as=0.1391p ps=1.055u w=0.535u l=0.5u
X129 a_32916_29860# _359_.B.t3 _461_.D VPWR.t6768 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X130 VPWR.t317 a_2364_20408# a_2276_20452# VPWR.t316 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X131 VPWR.t5837 a_64412_7431# a_64324_7528# VPWR.t2340 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X132 VPWR.t692 a_63740_9432# a_63652_9476# VPWR.t691 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X133 VPWR.t3080 a_49180_15271# a_49092_15368# VPWR.t1806 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X134 a_43620_29167# a_42820_29159.t2 VGND.t6727 VGND.t6726 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X135 VPWR.t909 _395_.A1 a_49044_28292# VPWR.t908 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X136 a_3708_13703# a_3620_13800# VGND.t783 VGND.t782 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X137 _355_.C.t3 a_28054_30196# VGND.t868 VGND.t71 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X138 VGND.t6330 _424_.B1.t6 a_50068_27508# VGND.t6329 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X139 a_20284_1592# a_20196_1636# VGND.t3083 VGND.t3082 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X140 a_46624_19715# a_46252_19759# VGND.t1821 VGND.t1820 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X141 _371_.ZN _371_.A1.t8 VGND.t6230 VGND.t6229 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X142 a_44252_1592# a_44164_1636# VGND.t1177 VGND.t1176 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X143 a_47636_25940# _397_.A2.t4 _284_.B VGND.t6716 nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X144 uo_out[0].t4 _284_.ZN.t20 a_40196_31048# VPWR.t6514 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X145 a_16588_27815# a_16500_27912# VGND.t451 VGND.t450 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X146 a_50532_24072# _399_.ZN VGND.t1189 VGND.t1188 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X147 a_42996_18840# a_43440_19325.t2 a_43392_19369# VGND.t6188 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X148 VPWR.t327 a_44364_17272# a_44276_17316# VPWR.t326 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X149 _459_.CLK.t15 a_41048_29816.t7 VGND.t6401 VGND.t6400 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X150 VPWR.t785 a_22748_2727# a_22660_2824# VPWR.t784 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X151 _459_.CLK.t7 a_41048_29816.t8 VPWR.t6683 VPWR.t6682 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X152 VPWR.t1327 _397_.A4 a_47636_23588# VPWR.t1326 pfet_06v0 ad=0.389p pd=2.02u as=0.1736p ps=1.18u w=0.56u l=0.5u
X153 VPWR.t461 a_36544_24419# a_36516_24831# VPWR.t460 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X154 a_59955_30600# a_60285_30600# a_60405_30644# VGND.t45 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X155 VPWR.t5130 a_46716_2727# a_46628_2824# VPWR.t5129 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X156 a_1916_26680# a_1828_26724# VGND.t1261 VGND.t1260 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X157 VPWR.t6642 _452_.CLK.t33 a_45284_19751.t0 VPWR.t6641 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X158 VPWR.t6465 _459_.CLK.t16 a_23668_25640.t0 VPWR.t6464 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X159 a_3708_1592# a_3620_1636# VGND.t5768 VGND.t2952 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X160 a_61052_26247# a_60964_26344# VGND.t478 VGND.t477 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X161 VPWR.t694 a_2364_14136# a_2276_14180# VPWR.t693 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X162 VPWR.t1254 a_32604_18407# a_32516_18504# VPWR.t1253 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X163 a_48396_16839# a_48308_16936# VGND.t1581 VGND.t1580 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X164 VGND.t1810 a_47776_20893# a_47728_20937# VGND.t1809 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X165 VPWR.t1353 a_2364_11000# a_2276_11044# VPWR.t1352 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X166 a_15244_24679# a_15156_24776# VGND.t1250 VGND.t1249 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X167 a_62844_27815# a_62756_27912# VGND.t2372 VGND.t2371 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X168 VPWR.t753 vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I VPWR.t752 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X169 a_15244_21543# a_15156_21640# VGND.t5729 VGND.t1041 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X170 a_15692_28248# a_15604_28292# VGND.t300 VGND.t299 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X171 VPWR.t5830 a_52764_1159# a_52676_1256# VPWR.t5829 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X172 a_62172_15271# a_62084_15368# VGND.t704 VGND.t703 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X173 a_29680_26724# _371_.A3 VPWR.t982 VPWR.t981 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X174 VPWR.t792 a_2364_7864# a_2276_7908# VPWR.t791 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X175 a_62763_28776# _251_.A1.t8 _250_.ZN VGND.t6685 nfet_06v0 ad=85.2f pd=0.95u as=0.21175p ps=1.41u w=0.71u l=0.6u
X176 a_63964_19975# a_63876_20072# VGND.t1067 VGND.t49 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X177 vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN VGND.t1071 VGND.t1070 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X178 a_35140_26680# _358_.A3 VPWR.t481 VPWR.t480 pfet_06v0 ad=0.1391p pd=1.055u as=0.4268p ps=2.175u w=0.535u l=0.5u
X179 VGND.t4966 _438_.A2 _435_.ZN VGND.t4965 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X180 a_48508_12135# a_48420_12232# VGND.t1815 VGND.t1814 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X181 a_37308_15271# a_37220_15368# VGND.t308 VGND.t307 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X182 VPWR.t2503 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN VPWR.t2502 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X183 VPWR.t5999 _421_.A1 _400_.ZN VPWR.t5998 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X184 a_64860_3160# a_64772_3204# VGND.t5611 VGND.t2960 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X185 VPWR.t615 a_23920_27555# a_23912_27967# VPWR.t614 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X186 a_47612_9432# a_47524_9476# VGND.t1288 VGND.t1287 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X187 a_67100_2727# a_67012_2824# VGND.t685 VGND.t684 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X188 a_59572_29076# _257_.B a_59348_29076# VGND.t317 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X189 _247_.ZN _252_.B a_59380_27508# VGND.t771 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X190 VPWR.t892 a_66204_4728# a_66116_4772# VPWR.t891 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X191 a_66876_14136# a_66788_14180# VGND.t880 VGND.t879 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X192 VPWR.t497 a_56796_14136# a_56708_14180# VPWR.t496 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X193 VGND.t4860 _475_.Q a_48529_22460# VGND.t4859 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X194 VPWR.t4995 a_27228_26247# a_27140_26344# VPWR.t4994 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X195 a_36076_18407# a_35988_18504# VGND.t765 VGND.t764 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X196 a_28891_25273# a_26916_25640.t3 a_28256_25597# VPWR.t6741 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X197 VGND.t6194 _459_.CLK.t17 a_20084_26023.t1 VGND.t6193 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X198 a_10204_29816# a_10116_29860# VGND.t2373 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X199 a_66876_11000# a_66788_11044# VGND.t1467 VGND.t1466 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X200 VPWR.t1248 a_56796_11000# a_56708_11044# VPWR.t1247 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X201 a_49988_21236# _424_.B1.t7 VGND.t6332 VGND.t6331 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X202 VGND.t872 _397_.Z a_48908_24080# VGND.t871 nfet_06v0 ad=0.23325p pd=1.48u as=93.59999f ps=1.02u w=0.78u l=0.6u
X203 a_40644_29480# _284_.ZN.t21 uo_out[1].t1 VPWR.t6515 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X204 a_39212_16839# a_39124_16936# VGND.t1393 VGND.t1392 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X205 a_41996_28777# _265_.ZN a_41872_28409# VPWR.t299 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X206 VGND.t1506 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I a_60524_25640# VGND.t1505 nfet_06v0 ad=0.2132p pd=1.34u as=98.39999f ps=1.06u w=0.82u l=0.6u
X207 VPWR.t800 _223_.ZN _350_.A2.t3 VPWR.t799 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X208 VPWR.t1336 a_47164_12568# a_47076_12612# VPWR.t1335 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X209 a_38971_18559# a_37408_18504# a_38336_18147# VGND.t1755 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X210 VPWR.t238 a_44296_24393.t15 clkbuf_1_0__f_clk.I.t14 VPWR.t237 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X211 a_30388_28776# _335_.ZN.t20 a_33720_28776# VGND.t6677 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X212 VGND.t5708 _285_.Z _296_.ZN VGND.t102 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X213 a_19388_2727# a_19300_2824# VGND.t5709 VGND.t1943 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X214 _371_.A3 _336_.Z VPWR.t4562 VPWR.t4561 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X215 VPWR.t3643 a_67996_4728# a_67908_4772# VPWR.t3642 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X216 a_65756_15704# a_65668_15748# VGND.t398 VGND.t397 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X217 VPWR.t2994 a_50860_18407# a_50772_18504# VPWR.t2993 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X218 _248_.B1 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I VGND.t4224 VGND.t4223 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X219 a_47636_25940# _381_.A2.t2 _284_.B VGND.t6648 nfet_06v0 ad=0.3608p pd=2.52u as=0.30965p ps=1.685u w=0.82u l=0.6u
X220 a_51868_9432# a_51780_9476# VGND.t4503 VGND.t4502 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X221 a_27172_24328# _352_.A2.t16 a_27552_24397# VGND.t6665 nfet_06v0 ad=0.1584p pd=1.6u as=57.59999f ps=0.68u w=0.36u l=0.6u
X222 VPWR.t1045 a_47612_14136# a_47524_14180# VPWR.t1044 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X223 VPWR.t4777 a_9084_2727# a_8996_2824# VPWR.t4776 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X224 a_32156_15704# a_32068_15748# VGND.t2878 VGND.t2877 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X225 a_30932_26020# _459_.Q.t2 a_30724_26020# VGND.t6649 nfet_06v0 ad=60.8f pd=0.7u as=0.1672p ps=1.64u w=0.38u l=0.6u
X226 a_67548_3160# a_67460_3204# VGND.t3524 VGND.t3523 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X227 VPWR.t1053 a_47612_11000# a_47524_11044# VPWR.t1052 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X228 VPWR.t5013 a_41048_17341# a_42404_17433# VPWR.t5012 pfet_06v0 ad=0.4554p pd=3.25u as=54f ps=0.66u w=0.36u l=0.5u
X229 a_12892_29383# a_12804_29480# VGND.t1149 VGND.t1148 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X230 a_26668_20408# a_26580_20452# VGND.t2872 VGND.t2871 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X231 VPWR.t4339 a_16588_20408# a_16500_20452# VPWR.t4338 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X232 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I VPWR.t5623 VPWR.t5622 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X233 a_66764_12135# a_66676_12232# VGND.t979 VGND.t978 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X234 a_65084_2727# a_64996_2824# VGND.t565 VGND.t564 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X235 VPWR.t5508 a_52988_26680# a_52900_26724# VPWR.t5507 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X236 VGND.t6636 _452_.Q.t4 a_42084_24072# VGND.t6635 nfet_06v0 ad=0.226p pd=1.515u as=88.2f ps=0.84u w=0.42u l=0.6u
X237 a_24512_25273# a_24080_25227# VPWR.t4423 VPWR.t4422 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X238 a_55564_12135# a_55476_12232# VGND.t5247 VGND.t5246 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X239 a_46848_20893# a_46476_20937# VPWR.t1047 VPWR.t1046 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X240 VPWR.t343 a_19948_26680# a_19860_26724# VPWR.t342 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X241 VPWR.t5495 a_42908_30951# a_42820_31048# VPWR.t5494 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X242 VPWR.t1010 a_64188_1592# a_64100_1636# VPWR.t1009 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X243 a_16796_27209# _467_.D a_16628_27209# VGND.t990 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X244 VPWR.t6545 a_48272_25156.t15 _474_.CLK.t1 VPWR.t6544 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X245 _287_.A1.t7 a_38472_30169# VGND.t4816 VGND.t1059 nfet_06v0 ad=0.1183p pd=0.975u as=0.2002p ps=1.79u w=0.455u l=0.6u
X246 VPWR.t4486 a_23980_23544# a_23892_23588# VPWR.t4485 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X247 a_28903_24776# _355_.B a_28679_24776# VPWR.t2990 pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X248 a_49496_30345# a_49152_30301.t2 a_48708_29816# VPWR.t6945 pfet_06v0 ad=0.1791p pd=1.355u as=0.1665p ps=1.285u w=0.36u l=0.5u
X249 VPWR.t3015 a_23084_29383# a_22996_29480# VPWR.t3014 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X250 VPWR.t1051 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I VPWR.t1050 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X251 VPWR.t1150 a_55228_27815# a_55140_27912# VPWR.t1149 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X252 a_51084_10567# a_50996_10664# VGND.t5731 VGND.t5730 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X253 a_37796_18191# a_36996_18183.t2 VGND.t6629 VGND.t6628 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X254 VGND.t5410 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN VGND.t537 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X255 VPWR.t5954 a_26668_21976# a_26580_22020# VPWR.t5953 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X256 a_40357_24776# _433_.ZN _436_.ZN VPWR.t568 pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X257 VPWR.t5706 a_44028_27815# a_43940_27912# VPWR.t5705 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X258 a_26160_27165# a_25867_26841# VGND.t3510 VGND.t3509 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X259 VPWR.t5008 a_66540_19975# a_66452_20072# VPWR.t5007 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X260 VPWR.t501 a_44700_2727# a_44612_2824# VPWR.t500 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X261 VGND.t781 _223_.ZN a_33312_28776# VGND.t780 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X262 a_54444_16839# a_54356_16936# VGND.t992 VGND.t991 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X263 VPWR.t5236 a_55340_19975# a_55252_20072# VPWR.t5235 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X264 VPWR.t1576 a_63516_19975# a_63428_20072# VPWR.t1575 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X265 VPWR.t436 a_33520_25597# a_33492_25273# VPWR.t435 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X266 VPWR.t865 a_18604_20408# a_18516_20452# VPWR.t864 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X267 VPWR.t5453 a_62396_12568# a_62308_12612# VPWR.t5452 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X268 a_38336_18147# a_37964_18191# VPWR.t4384 VPWR.t4383 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X269 a_18492_1592# a_18404_1636# VGND.t1121 VGND.t1120 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X270 VPWR.t5633 a_45036_28248# a_44948_28292# VPWR.t5632 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X271 a_38523_27967# a_36548_27591.t2 a_37888_27555# VPWR.t6612 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X272 VPWR.t6192 a_51196_12568# a_51108_12612# VPWR.t6191 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X273 a_43232_29480# a_42820_29159.t3 VGND.t6729 VGND.t6728 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X274 a_45360_29977# a_44632_30206# VPWR.t838 VPWR.t837 pfet_06v0 ad=50.4f pd=0.64u as=0.23p ps=1.54u w=0.36u l=0.5u
X275 a_42392_22825.t13 clkbuf_1_0__f_clk.I.t32 VGND.t245 VGND.t244 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X276 VPWR.t4354 a_50636_13703# a_50548_13800# VPWR.t4353 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X277 a_64300_10567# a_64212_10664# VGND.t463 VGND.t462 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X278 VPWR.t5646 a_64412_9432# a_64324_9476# VPWR.t5077 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X279 VPWR.t6685 a_41048_29816.t9 _459_.CLK.t6 VPWR.t6684 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X280 a_17860_28777# a_17060_28776.t2 VGND.t6592 VGND.t6591 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X281 VPWR.t5697 a_25212_1159# a_25124_1256# VPWR.t5696 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X282 VPWR.t408 a_18096_27165# a_18088_26841# VPWR.t407 pfet_06v0 ad=0.2619p pd=1.685u as=50.4f ps=0.64u w=0.36u l=0.5u
X283 a_1468_18407# a_1380_18504# VGND.t3508 VGND.t3507 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X284 VPWR.t5137 a_10204_29816# a_10116_29860# VPWR.t5136 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X285 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN VGND.t4566 VGND.t4565 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X286 _441_.B _430_.ZN a_38759_24072# VGND.t4673 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X287 VPWR.t1193 a_58252_18407# a_58164_18504# VPWR.t1192 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X288 VPWR.t3641 a_44924_15704# a_44836_15748# VPWR.t3640 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X289 VPWR.t5700 a_62844_14136# a_62756_14180# VPWR.t5699 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X290 a_15692_24679# a_15604_24776# VGND.t4606 VGND.t2743 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X291 VPWR.t4860 a_58140_9432# a_58052_9476# VPWR.t4859 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X292 a_36636_26247# a_36548_26344# VGND.t5241 VGND.t5240 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X293 VGND.t5797 a_19328_28733# uio_out[6].t7 VGND.t5796 nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X294 VPWR.t3025 a_40220_1592# a_40132_1636# VPWR.t3024 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X295 VGND.t6402 a_41048_29816.t10 _459_.CLK.t14 VGND.t6400 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X296 VPWR.t1195 a_62844_11000# a_62756_11044# VPWR.t1194 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X297 VPWR.t5710 a_51644_14136# a_51556_14180# VPWR.t5709 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X298 a_15692_21543# a_15604_21640# VGND.t3166 VGND.t3165 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X299 VPWR.t5606 a_51644_11000# a_51556_11044# VPWR.t5605 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X300 a_25436_23111# a_25348_23208# VGND.t4513 VGND.t4512 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X301 a_6396_29816# a_6308_29860# VGND.t4443 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X302 a_52988_1592# a_52900_1636# VGND.t4635 VGND.t4634 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X303 VPWR.t1466 a_53212_12568# a_53124_12612# VPWR.t1465 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X304 a_37756_15271# a_37668_15368# VGND.t4755 VGND.t4754 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X305 a_55208_22505# a_54864_22461.t2 a_54420_21976# VPWR.t6595 pfet_06v0 ad=0.1791p pd=1.355u as=0.1665p ps=1.285u w=0.36u l=0.5u
X306 VPWR.t5619 a_37084_21543# a_36996_21640# VPWR.t5618 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X307 a_18760_29032# uio_out[7].t8 VGND.t6583 VGND.t6582 nfet_06v0 ad=93.59999f pd=0.88u as=0.218p ps=1.52u w=0.36u l=0.6u
X308 a_47612_2727# a_47524_2824# VGND.t1135 VGND.t1134 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X309 VPWR.t6020 a_66652_5863# a_66564_5960# VPWR.t5505 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X310 VPWR.t5023 a_20672_30301# uio_out[5].t3 VPWR.t5022 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X311 VGND.t6572 _448_.Q.t2 _323_.A3 VGND.t6571 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X312 VGND.t6718 _397_.A2.t5 a_46984_23588# VGND.t6717 nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X313 VPWR.t3013 a_66652_2727# a_66564_2824# VPWR.t2509 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X314 VPWR.t362 a_27676_26247# a_27588_26344# VPWR.t361 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X315 a_63524_29098# _229_.I.t2 VGND.t6561 VGND.t6560 nfet_06v0 ad=85.2f pd=0.95u as=0.3124p ps=2.3u w=0.71u l=0.6u
X316 VPWR.t1199 a_17148_2727# a_17060_2824# VPWR.t1198 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X317 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I VPWR.t5604 VPWR.t5603 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X318 a_10652_29816# a_10564_29860# VGND.t1104 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X319 VPWR.t2484 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I VPWR.t2483 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X320 VPWR.t4765 a_32604_17272# a_32516_17316# VPWR.t4764 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X321 VPWR.t5968 a_65980_1592# a_65892_1636# VPWR.t5967 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X322 _352_.A2.t13 _350_.A1.t3 a_30520_27508# VGND.t6352 nfet_06v0 ad=0.2132p pd=1.34u as=98.39999f ps=1.06u w=0.82u l=0.6u
X323 a_29808_29167# a_27588_29159.t2 a_29563_29535# VGND.t6555 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X324 a_39660_16839# a_39572_16936# VGND.t4613 VGND.t4612 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X325 a_43328_18559# a_42896_18504# VPWR.t5976 VPWR.t5975 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X326 VPWR.t5532 a_19612_24679# a_19524_24776# VPWR.t5531 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X327 a_31516_28292# _337_.ZN VPWR.t5143 VPWR.t5142 pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X328 a_41696_24072# _304_.A1.t3 a_41488_24072# VGND.t6315 nfet_06v0 ad=67.2f pd=0.74u as=0.1848p ps=1.72u w=0.42u l=0.6u
X329 VGND.t6542 _437_.A1.t2 a_39480_28776# VGND.t6541 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X330 VPWR.t1578 a_62396_9432# a_62308_9476# VPWR.t1577 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X331 VPWR.t240 a_44296_24393.t16 clkbuf_1_0__f_clk.I.t13 VPWR.t239 pfet_06v0 ad=0.428p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
X332 a_45088_29123# a_44795_29535# VPWR.t5480 VPWR.t5479 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X333 VPWR.t957 a_23196_1159# a_23108_1256# VPWR.t956 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X334 a_32716_20408# a_32628_20452# VGND.t5398 VGND.t5397 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X335 VPWR.t1070 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN _245_.I1 VPWR.t1069 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X336 VPWR.t4753 a_47164_1159# a_47076_1256# VPWR.t4752 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X337 a_51240_23340# _384_.A1 VGND.t918 VGND.t917 nfet_06v0 ad=0.126p pd=1.06u as=0.1584p ps=1.6u w=0.36u l=0.6u
X338 VGND.t396 a_18096_27165# a_18048_27209# VGND.t395 nfet_06v0 ad=0.2333p pd=1.555u as=43.2f ps=0.6u w=0.36u l=0.6u
X339 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[1\].I VPWR.t1431 VPWR.t1430 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X340 a_61612_12135# a_61524_12232# VGND.t2366 VGND.t2365 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X341 a_52512_19715# a_52024_20083# a_52944_19759# VGND.t428 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X342 _304_.B a_54432_31128# VGND.t4518 VGND.t4514 nfet_06v0 ad=0.1183p pd=0.975u as=0.2002p ps=1.79u w=0.455u l=0.6u
X343 a_21868_27208# _455_.Q.t2 _455_.D VGND.t6534 nfet_06v0 ad=0.1312p pd=1.14u as=0.2569p ps=1.56u w=0.82u l=0.6u
X344 a_51868_2727# a_51780_2824# VGND.t5406 VGND.t5405 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X345 VPWR.t3655 a_62172_1592# a_62084_1636# VPWR.t3654 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X346 VPWR.t1072 a_58028_13703# a_57940_13800# VPWR.t1071 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X347 VPWR.t5698 a_2812_24679# a_2724_24776# VPWR.t1358 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X348 a_46716_18407# a_46628_18504# VGND.t3490 VGND.t3489 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X349 uo_out[5].t3 _290_.ZN VGND.t1142 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X350 a_32904_28776# _223_.ZN VGND.t779 VGND.t778 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X351 a_39216_18191# a_36996_18183.t3 a_38971_18559# VGND.t6630 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X352 VPWR.t6138 a_63404_23544# a_63316_23588# VPWR.t5291 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X353 VPWR.t5956 a_62060_10567# a_61972_10664# VPWR.t5955 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X354 uo_out[6].t4 _287_.A1.t10 a_32132_27912# VPWR.t6777 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X355 _312_.ZN _304_.A1.t4 VGND.t6317 VGND.t6316 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X356 _324_.B.t3 _305_.A2 a_42168_22504# VGND.t2876 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X357 a_21740_30951# a_21652_31048# VGND.t5130 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X358 _448_.Q.t0 a_37360_19325# VPWR.t5704 VPWR.t5703 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X359 a_44296_24393.t0 clk.t0 VPWR.t6831 VPWR.t6830 pfet_06v0 ad=0.2542p pd=1.44u as=0.428p ps=2.02u w=0.82u l=0.5u
X360 VPWR.t5597 _284_.B _284_.ZN.t19 VPWR.t5596 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X361 a_45596_2727# a_45508_2824# VGND.t5430 VGND.t5429 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X362 VPWR.t5946 a_21516_21976# a_21428_22020# VPWR.t5945 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X363 a_40668_26247# a_40580_26344# VGND.t480 VGND.t479 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X364 a_10540_30951# a_10452_31048# VGND.t1111 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X365 a_1020_7864# a_932_7908# VGND.t476 VGND.t475 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X366 VPWR.t1041 a_65420_16839# a_65332_16936# VPWR.t1040 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X367 VGND.t606 vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN VGND.t605 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X368 _432_.ZN _325_.A1.t4 a_40880_23588# VPWR.t224 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X369 VGND.t820 a_44632_30206# _388_.B VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X370 VPWR.t5712 a_2364_16839# a_2276_16936# VPWR.t5711 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X371 a_56348_12568# a_56260_12612# VGND.t5438 VGND.t5437 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X372 a_20508_1159# a_20420_1256# VGND.t411 VGND.t410 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X373 a_1020_4728# a_932_4772# VGND.t1407 VGND.t1406 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X374 VGND.t6356 _452_.CLK.t34 a_39124_27208.t1 VGND.t6355 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X375 a_52988_15271# a_52900_15368# VGND.t2856 VGND.t2855 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X376 a_47271_21640# _419_.Z _475_.D VPWR.t4464 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X377 VPWR.t4807 a_59036_11000# a_58948_11044# VPWR.t4806 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X378 _325_.A1.t1 a_42392_19243# VPWR.t589 VPWR.t588 pfet_06v0 ad=0.3172p pd=1.74u as=0.854p ps=3.84u w=1.22u l=0.5u
X379 a_17120_27209# a_16240_26795# a_16796_27209# VGND.t5416 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X380 VPWR.t3012 a_43020_16839# a_42932_16936# VPWR.t3011 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X381 vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN VPWR.t4414 VPWR.t4413 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X382 a_62172_18840# a_62084_18884# VGND.t5151 VGND.t5150 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X383 a_19280_28777# a_17060_28776.t3 a_19035_28409# VGND.t6593 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X384 VPWR.t5598 a_55676_27815# a_55588_27912# VPWR.t2521 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X385 a_64412_4295# a_64324_4392# VGND.t4549 VGND.t4548 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X386 VGND.t207 _330_.A1.t4 _316_.ZN VGND.t206 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X387 a_45820_15704# a_45732_15748# VGND.t5434 VGND.t5433 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X388 VPWR.t5398 a_44476_27815# a_44388_27912# VPWR.t5397 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X389 a_3708_17272# a_3620_17316# VGND.t5499 VGND.t5498 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X390 _285_.Z a_38584_28292# VGND.t3895 VGND.t3894 nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X391 a_14796_25112# a_14708_25156# VGND.t2218 VGND.t2217 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X392 VPWR.t3595 a_1020_10567# a_932_10664# VPWR.t3594 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X393 a_54892_16839# a_54804_16936# VGND.t1832 VGND.t1831 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X394 a_18044_29816# a_17956_29860# VGND.t3966 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X395 a_46268_9432# a_46180_9476# VGND.t3898 VGND.t3897 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X396 a_29916_1159# a_29828_1256# VGND.t1735 VGND.t1734 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X397 VPWR.t2302 a_2812_15271# a_2724_15368# VPWR.t1567 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X398 a_14796_21976# a_14708_22020# VGND.t3978 VGND.t3977 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X399 VPWR.t2619 a_34844_24679# a_34756_24776# VPWR.t2618 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X400 VPWR.t1793 a_53100_18407# a_53012_18504# VPWR.t1792 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X401 VPWR.t471 a_63964_19975# a_63876_20072# VPWR.t470 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X402 VPWR.t3606 a_18940_2727# a_18852_2824# VPWR.t3605 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X403 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN VPWR.t5322 VPWR.t5321 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X404 _355_.ZN _336_.Z a_28903_24776# VPWR.t4560 pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X405 VPWR.t1996 a_23644_24679# a_23556_24776# VPWR.t1995 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X406 VPWR.t1197 a_6396_29816# a_6308_29860# VPWR.t1196 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X407 VPWR.t2583 a_4156_6296# a_4068_6340# VPWR.t2582 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X408 a_17932_20408# a_17844_20452# VGND.t3374 VGND.t369 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X409 hold1.Z a_44038_21236# VPWR.t6240 VPWR.t6239 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X410 VPWR.t4229 a_45484_28248# a_45396_28292# VPWR.t4228 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X411 VPWR.t4131 a_4156_3160# a_4068_3204# VPWR.t4130 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X412 VPWR.t6281 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN VPWR.t6280 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X413 a_33028_27912# _287_.A2 VPWR.t2034 VPWR.t2033 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X414 _474_.CLK.t2 a_48272_25156.t16 VGND.t6262 VGND.t6261 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X415 a_58228_27912# _241_.Z VPWR.t3565 VPWR.t3564 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X416 a_31708_1592# a_31620_1636# VGND.t1119 VGND.t1118 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X417 _416_.A1.t3 _324_.C.t9 VGND.t6499 VGND.t6498 nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X418 VPWR.t6238 a_64860_7431# a_64772_7528# VPWR.t3432 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X419 a_48060_13703# a_47972_13800# VGND.t3572 VGND.t3571 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X420 VPWR.t5240 a_7068_29383# a_6980_29480# VPWR.t5239 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X421 VGND.t4122 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I VGND.t4121 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X422 a_15132_29383# a_15044_29480# VGND.t3883 VGND.t3882 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X423 VPWR.t3867 a_21404_2727# a_21316_2824# VPWR.t3866 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X424 VPWR.t1231 a_10652_29816# a_10564_29860# VPWR.t1230 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X425 a_62284_23544# a_62196_23588# VGND.t1320 VGND.t1319 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X426 VPWR.t6321 a_23084_28248# a_22996_28292# VPWR.t6320 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X427 a_32604_15271# a_32516_15368# VGND.t3805 VGND.t3804 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X428 a_47483_20569# a_45508_20936.t2 a_46848_20893# VPWR.t197 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X429 a_35088_20893# a_34716_20937# VPWR.t4013 VPWR.t4012 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X430 VPWR.t3268 hold2.Z _265_.ZN VPWR.t3267 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X431 a_25436_1592# a_25348_1636# VGND.t5727 VGND.t5726 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X432 VPWR.t6267 a_20732_1592# a_20644_1636# VPWR.t6266 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X433 a_51912_20452# _419_.Z _424_.B2 VPWR.t4463 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X434 VPWR.t1261 a_67548_18840# a_67460_18884# VPWR.t1260 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X435 VPWR.t4053 a_23084_25112# a_22996_25156# VPWR.t4052 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X436 a_30847_27208# _336_.Z VGND.t4415 VGND.t4414 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X437 VPWR.t3562 a_17932_21976# a_17844_22020# VPWR.t381 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X438 a_49404_1592# a_49316_1636# VGND.t3815 VGND.t1867 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X439 VPWR.t4248 a_49600_30180# a_49496_30345# VPWR.t4247 pfet_06v0 ad=0.1044p pd=0.94u as=0.1791p ps=1.355u w=0.36u l=0.5u
X440 VPWR.t3408 a_44700_1592# a_44612_1636# VPWR.t924 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X441 VPWR.t3135 a_15132_2727# a_15044_2824# VPWR.t3134 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X442 VPWR.t1458 a_11324_29383# a_11236_29480# VPWR.t1457 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X443 VPWR.t5559 a_48172_18840# a_48084_18884# VPWR.t5558 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X444 VGND.t6544 _437_.A1.t3 _437_.ZN VGND.t6543 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X445 VPWR.t3092 a_33724_23111# a_33636_23208# VPWR.t3091 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X446 VPWR.t6870 _229_.I.t3 _243_.A1 VPWR.t6869 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X447 a_48508_30951# a_48420_31048# VGND.t2455 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X448 VPWR.t5900 a_67548_15704# a_67460_15748# VPWR.t5899 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X449 VPWR.t1456 a_40644_17272# a_40040_17675# VPWR.t1455 pfet_06v0 ad=0.23p pd=1.54u as=0.352p ps=2.48u w=0.8u l=0.5u
X450 VPWR.t5447 _323_.A3 a_36836_20072# VPWR.t5446 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X451 VPWR.t3783 a_52428_10567# a_52340_10664# VPWR.t3782 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X452 VPWR.t1776 a_39100_2727# a_39012_2824# VPWR.t1775 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X453 a_35816_21192# _447_.Q.t3 a_36204_21327# VGND.t6301 nfet_06v0 ad=0.1606p pd=1.61u as=58.39999f ps=0.685u w=0.365u l=0.6u
X454 VPWR.t3272 a_26220_23544# a_26132_23588# VPWR.t3271 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X455 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I VGND.t2362 VGND.t2361 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X456 VPWR.t4114 a_5052_20408# a_4964_20452# VPWR.t4113 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X457 a_46198_27060# _424_.A2.t6 VPWR.t188 VPWR.t187 pfet_06v0 ad=0.5368p pd=3.32u as=0.4941p ps=2.03u w=1.22u l=0.5u
X458 a_33776_29123# a_33483_29535# VGND.t3376 VGND.t3375 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X459 a_25884_23111# a_25796_23208# VGND.t3764 VGND.t3763 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X460 a_39300_29480# _293_.A2 VPWR.t5926 VPWR.t5925 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X461 VGND.t6467 _359_.B.t4 _359_.ZN VGND.t6466 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X462 a_54444_26680# a_54356_26724# VGND.t6058 VGND.t6057 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X463 VGND.t6429 _402_.A1.t5 a_38584_28292# VGND.t6428 nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X464 VPWR.t483 a_1020_7864# a_932_7908# VPWR.t482 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X465 VPWR.t3875 a_51420_1159# a_51332_1256# VPWR.t3874 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X466 uo_out[1].t5 _284_.ZN.t22 VGND.t6238 VGND.t6237 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X467 VPWR.t4025 a_53660_12568# a_53572_12612# VPWR.t4024 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X468 a_26108_30951# a_26020_31048# VGND.t3255 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X469 a_28556_29167# _373_.ZN a_28388_29167# VGND.t1345 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X470 _335_.ZN.t3 _334_.A1 VPWR.t2362 VPWR.t2361 pfet_06v0 ad=0.2197p pd=1.365u as=0.4056p ps=1.805u w=0.845u l=0.5u
X471 _402_.B _402_.A1.t6 a_46356_24072# VGND.t6430 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X472 a_38971_18559# a_36996_18183.t4 a_38336_18147# VPWR.t6941 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X473 VGND.t1254 _397_.A4 a_46984_23588# VGND.t1253 nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X474 VPWR.t4805 _474_.Q _384_.A3.t7 VPWR.t4804 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X475 VPWR.t3365 a_62508_12135# a_62420_12232# VPWR.t3364 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X476 a_64300_23544# a_64212_23588# VGND.t4253 VGND.t4252 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X477 VPWR.t7009 _251_.A1.t9 a_55956_25940# VPWR.t7008 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X478 a_62620_17272# a_62532_17316# VGND.t5712 VGND.t3718 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X479 a_1020_19975# a_932_20072# VGND.t5066 VGND.t622 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X480 VPWR.t3143 a_40038_28720# uo_out[7].t2 VPWR.t3142 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X481 _399_.A1 _218_.ZN VPWR.t3773 VPWR.t3772 pfet_06v0 ad=0.4012p pd=1.85u as=0.4972p ps=3.14u w=1.13u l=0.5u
X482 _336_.A1 a_29184_25597# VGND.t4052 VGND.t4051 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X483 a_31964_28292# _371_.A1.t9 _350_.A2.t8 VPWR.t6508 pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X484 a_24316_1159# a_24228_1256# VGND.t6030 VGND.t6029 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X485 a_32828_1159# a_32740_1256# VGND.t3087 VGND.t3086 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X486 VPWR.t1402 a_67548_7431# a_67460_7528# VPWR.t1401 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X487 a_51420_17272# a_51332_17316# VGND.t3561 VGND.t3560 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X488 VPWR.t4188 a_41160_29083# uo_out[3].t3 VPWR.t4187 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X489 a_4604_26680# a_4516_26724# VGND.t3415 VGND.t3414 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X490 a_24316_2727# a_24228_2824# VGND.t3293 VGND.t3292 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X491 VPWR.t5973 a_27676_1159# a_27588_1256# VPWR.t5972 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X492 a_2364_12568# a_2276_12612# VGND.t3722 VGND.t1839 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X493 a_27900_23111# a_27812_23208# VGND.t4091 VGND.t4090 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X494 a_29136_25641# a_26916_25640.t4 a_28891_25273# VGND.t6472 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X495 VPWR.t3465 a_5052_14136# a_4964_14180# VPWR.t3464 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X496 a_8860_29816# a_8772_29860# VGND.t3085 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X497 VPWR.t5578 a_43356_2727# a_43268_2824# VPWR.t5577 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X498 VGND.t176 uio_in[0].t0 a_51791_30644# VGND.t45 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X499 VPWR.t6719 _402_.A1.t7 a_38772_28292# VPWR.t6718 pfet_06v0 ad=0.4005p pd=2.12u as=0.1456p ps=1.08u w=0.56u l=0.5u
X500 a_4940_8999# a_4852_9096# VGND.t3965 VGND.t3964 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X501 a_44571_26841# a_43008_26795# a_43936_27165# VGND.t5760 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X502 VPWR.t3261 a_5052_11000# a_4964_11044# VPWR.t3260 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X503 VPWR.t921 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN VPWR.t920 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X504 a_18044_2727# a_17956_2824# VGND.t5212 VGND.t1128 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X505 VPWR.t3437 a_66652_4728# a_66564_4772# VPWR.t3436 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X506 a_47388_1592# a_47300_1636# VGND.t3089 VGND.t3088 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X507 a_42996_18840# a_43400_18909# a_43344_19001# VPWR.t3898 pfet_06v0 ad=0.1665p pd=1.285u as=50.4f ps=0.64u w=0.36u l=0.5u
X508 a_4940_5863# a_4852_5960# VGND.t3580 VGND.t3579 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X509 VGND.t1830 a_47552_19715# a_47504_19759# VGND.t1829 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X510 a_44784_25987.t1 _474_.CLK.t34 VGND.t6447 VGND.t6446 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X511 VPWR.t4029 a_37084_2727# a_36996_2824# VPWR.t4028 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X512 VPWR.t6039 a_58476_13703# a_58388_13800# VPWR.t6038 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X513 VPWR.t1020 a_55312_22340# a_55208_22505# VPWR.t1019 pfet_06v0 ad=0.1044p pd=0.94u as=0.1791p ps=1.355u w=0.36u l=0.5u
X514 VPWR.t166 _336_.A2.t2 a_28820_24072# VPWR.t165 pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X515 _470_.Q a_44864_27165# VPWR.t3374 VPWR.t3373 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X516 a_60268_13703# a_60180_13800# VGND.t590 VGND.t589 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X517 a_41088_17757.t0 _452_.CLK.t35 VPWR.t6644 VPWR.t6643 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X518 VPWR.t4193 a_62284_26680# a_62196_26724# VPWR.t4192 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X519 VPWR.t5576 a_17148_1592# a_17060_1636# VPWR.t952 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X520 VPWR.t3969 a_63852_23544# a_63764_23588# VPWR.t1036 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X521 VGND.t6589 uio_out[6].t8 a_20003_29611# VGND.t6588 nfet_06v0 ad=0.2288p pd=1.58u as=93.59999f ps=0.88u w=0.36u l=0.6u
X522 a_43132_27815# a_43044_27912# VGND.t2987 VGND.t2986 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X523 VPWR.t2032 _287_.A2 a_32580_27912# VPWR.t2031 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X524 VPWR.t4118 a_18044_29816# a_17956_29860# VPWR.t4117 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X525 a_50524_9432# a_50436_9476# VGND.t3143 VGND.t3142 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X526 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I VPWR.t1586 VPWR.t1585 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X527 a_25764_29977# a_24452_30344.t2 a_25420_30345# VPWR.t157 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X528 _436_.B a_41392_27165# VGND.t804 VGND.t803 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X529 VPWR.t1716 a_21964_21976# a_21876_22020# VPWR.t1715 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X530 a_33376_23659# a_32964_24072.t2 VGND.t152 VGND.t151 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X531 a_66204_3160# a_66116_3204# VGND.t5812 VGND.t2640 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X532 a_56796_12568# a_56708_12612# VGND.t3474 VGND.t3473 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X533 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I VGND.t3568 VGND.t3567 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X534 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN VGND.t2250 VGND.t2249 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X535 a_29664_29977# a_29232_29931# VPWR.t1032 VPWR.t1031 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X536 a_33052_19975# a_32964_20072# VGND.t3354 VGND.t3353 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X537 VGND.t6480 _287_.A1.t11 uo_out[5].t9 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X538 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t1195 VGND.t1194 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X539 VPWR.t3467 a_59484_11000# a_59396_11044# VPWR.t3466 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X540 VGND.t1513 a_41536_17636# a_41432_17801# VGND.t1512 nfet_06v0 ad=0.2637p pd=1.825u as=93.59999f ps=0.88u w=0.36u l=0.6u
X541 a_36636_26680# a_36548_26724# VGND.t5017 VGND.t5016 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X542 a_43788_29167# _480_.Q a_43620_29167# VGND.t4929 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X543 VPWR.t2057 a_58924_12135# a_58836_12232# VPWR.t2056 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X544 a_47164_14136# a_47076_14180# VGND.t5168 VGND.t5167 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X545 VPWR.t146 _294_.ZN.t3 a_35156_29860# VPWR.t145 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X546 a_40038_28720# _234_.ZN VGND.t3447 VGND.t3446 nfet_06v0 ad=0.3608p pd=2.52u as=0.2911p ps=1.53u w=0.82u l=0.6u
X547 a_46820_20569# a_45508_20936.t3 a_46476_20937# VPWR.t198 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X548 a_47164_11000# a_47076_11044# VGND.t3896 VGND.t2927 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X549 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN VPWR.t3891 VPWR.t3890 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X550 VPWR.t3558 a_2812_23544# a_2724_23588# VPWR.t3099 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X551 a_3708_9432# a_3620_9476# VGND.t3874 VGND.t997 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X552 a_5724_30951# a_5636_31048# VGND.t3625 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X553 a_19140_29612# uio_out[7].t9 VPWR.t6895 VPWR.t6894 pfet_06v0 ad=0.1456p pd=1.08u as=0.4005p ps=2.12u w=0.56u l=0.5u
X554 a_67996_3160# a_67908_3204# VGND.t3702 VGND.t3701 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X555 VGND.t6292 _350_.A2.t20 a_30912_27508# VGND.t6291 nfet_06v0 ad=0.3608p pd=2.52u as=98.39999f ps=1.06u w=0.82u l=0.6u
X556 a_43396_27209# a_42596_27208.t2 VGND.t142 VGND.t141 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X557 VGND.t6195 _459_.CLK.t18 a_18404_30344.t1 VGND.t139 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X558 a_3708_6296# a_3620_6340# VGND.t5750 VGND.t4080 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X559 VPWR.t4003 a_2364_18840# a_2276_18884# VPWR.t2513 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X560 VPWR.t5966 a_61724_18407# a_61636_18504# VPWR.t5965 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X561 a_50280_19369# a_49896_18909# a_49492_18840# VGND.t5243 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X562 a_23420_1592# a_23332_1636# VGND.t5775 VGND.t5774 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X563 a_44812_17272# a_44724_17316# VGND.t5714 VGND.t5713 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X564 VGND.t5166 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I VGND.t5165 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X565 VPWR.t5828 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN VPWR.t5827 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X566 _462_.D _365_.ZN VGND.t3409 VGND.t102 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X567 _324_.B.t5 _304_.B a_44948_22020# VPWR.t4701 pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X568 a_31932_26247# a_31844_26344# VGND.t3634 VGND.t3633 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X569 VPWR.t4246 a_2364_15704# a_2276_15748# VPWR.t1085 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X570 a_50084_24328# _398_.C VGND.t3158 VGND.t3157 nfet_06v0 ad=0.176p pd=1.68u as=0.104p ps=0.92u w=0.4u l=0.6u
X571 _330_.A1.t1 a_46198_27060# VPWR.t1622 VPWR.t1621 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X572 _316_.ZN _317_.A2 VGND.t2454 VGND.t2453 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X573 _417_.A2.t0 _419_.A4 VPWR.t4136 VPWR.t4135 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X574 a_47612_12568# a_47524_12612# VGND.t2951 VGND.t2950 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X575 VGND.t1596 a_22992_27555# a_22944_27599# VGND.t1595 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X576 a_31932_23111# a_31844_23208# VGND.t2356 VGND.t2355 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X577 VGND.t231 _325_.A1.t5 _432_.ZN VGND.t230 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X578 a_33164_24679# a_33076_24776# VGND.t3885 VGND.t3884 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X579 _452_.CLK.t0 a_42392_22825.t14 VGND.t6597 VGND.t6596 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X580 a_45644_26399# a_45128_26031# VPWR.t2651 VPWR.t2650 pfet_06v0 ad=43.2f pd=0.6u as=0.1044p ps=0.94u w=0.36u l=0.5u
X581 a_15580_29383# a_15492_29480# VGND.t3706 VGND.t3705 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X582 a_49936_19325.t1 _474_.CLK.t35 VGND.t6449 VGND.t6448 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X583 a_29356_20408# a_29268_20452# VGND.t567 VGND.t566 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X584 VGND.t120 _281_.ZN.t4 _282_.ZN VGND.t119 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X585 VGND.t3942 _247_.B _247_.ZN VGND.t3941 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X586 VPWR.t3728 a_32380_21543# a_32292_21640# VPWR.t3727 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X587 a_66428_15271# a_66340_15368# VGND.t5328 VGND.t5023 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X588 a_42811_19668# _325_.A1.t6 _303_.ZN VGND.t232 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X589 a_29916_1592# a_29828_1636# VGND.t4105 VGND.t2161 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X590 VGND.t5371 _327_.Z a_40684_19368# VGND.t5370 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X591 VPWR.t3964 a_18716_21543# a_18628_21640# VPWR.t3963 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X592 VPWR.t2581 a_27668_31048# a_27668_31048# VPWR.t2580 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X593 VPWR.t6630 _230_.I.t3 a_62564_29032# VPWR.t6629 pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X594 a_28124_1159# a_28036_1256# VGND.t2976 VGND.t2975 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X595 a_36636_1159# a_36548_1256# VGND.t3208 VGND.t3207 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X596 VPWR.t3851 a_67996_18840# a_67908_18884# VPWR.t3850 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X597 _304_.ZN.t3 _304_.B VPWR.t4700 VPWR.t4699 pfet_06v0 ad=0.2808p pd=1.6u as=0.3918p ps=1.815u w=1.08u l=0.5u
X598 VPWR.t4233 a_2812_8999# a_2724_9096# VPWR.t2725 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X599 VPWR.t1604 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I VPWR.t1603 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X600 VPWR.t3920 a_11772_29383# a_11684_29480# VPWR.t3919 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X601 a_48956_30951# a_48868_31048# VGND.t2829 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X602 VPWR.t5206 a_67996_15704# a_67908_15748# VPWR.t5205 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X603 VPWR.t6547 a_48272_25156.t17 _474_.CLK.t3 VPWR.t6546 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X604 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN VPWR.t2526 VPWR.t2525 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X605 clkbuf_1_0__f_clk.I.t31 a_44296_24393.t17 VGND.t243 VGND.t242 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X606 VPWR.t5556 a_52876_10567# a_52788_10664# VPWR.t5555 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X607 VGND.t1652 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN VGND.t1651 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X608 a_26668_23544# a_26580_23588# VGND.t1517 VGND.t1516 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X609 a_44028_15271# a_43940_15368# VGND.t3557 VGND.t3556 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X610 _411_.A2.t1 _397_.A2.t6 VPWR.t7036 VPWR.t7035 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X611 VPWR.t107 _294_.A2.t2 a_35818_29860# VPWR.t106 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X612 a_22452_27599# a_21652_27591.t2 VGND.t98 VGND.t97 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X613 VPWR.t5982 a_18940_1592# a_18852_1636# VPWR.t4612 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X614 VPWR.t3937 a_31932_1159# a_31844_1256# VPWR.t3936 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X615 VGND.t3316 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN VGND.t3315 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X616 a_33152_22091# a_32740_22504.t2 VPWR.t99 VPWR.t98 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X617 a_43344_19001# a_42392_19243# VPWR.t587 VPWR.t586 pfet_06v0 ad=50.4f pd=0.64u as=0.23p ps=1.54u w=0.36u l=0.5u
X618 VPWR.t1462 a_8860_29816# a_8772_29860# VPWR.t1461 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X619 a_49637_28776# _404_.A1 VGND.t3678 VGND.t3677 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X620 VPWR.t1836 a_4940_21543# a_4852_21640# VPWR.t1835 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X621 a_54892_26680# a_54804_26724# VGND.t3114 VGND.t3113 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X622 VPWR.t5562 a_29356_21976# a_29268_22020# VPWR.t5561 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X623 a_26556_30951# a_26468_31048# VGND.t2408 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X624 VPWR.t4046 a_34396_18840# a_34308_18884# VPWR.t4045 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X625 VGND.t5356 a_46848_20893# a_46800_20937# VGND.t5355 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X626 VPWR.t3968 a_64860_9432# a_64772_9476# VPWR.t3967 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X627 a_17036_25112# a_16948_25156# VGND.t5679 VGND.t2124 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X628 a_22300_2727# a_22212_2824# VGND.t5267 VGND.t5266 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X629 a_51644_1592# a_51556_1636# VGND.t3735 VGND.t3734 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X630 VPWR.t4027 a_25660_1159# a_25572_1256# VPWR.t4026 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X631 VPWR.t3404 a_54332_20408# a_54244_20452# VPWR.t3403 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X632 VPWR.t3289 a_1916_21543# a_1828_21640# VPWR.t3288 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X633 a_62396_14136# a_62308_14180# VGND.t5752 VGND.t5751 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X634 a_42252_20936# _303_.ZN _304_.ZN.t1 VGND.t2814 nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X635 a_42161_24776# hold1.Z hold2.I VPWR.t3570 pfet_06v0 ad=0.32805p pd=1.755u as=0.37665p ps=1.835u w=1.215u l=0.5u
X636 VPWR.t3367 a_9532_29383# a_9444_29480# VPWR.t3366 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X637 VPWR.t5964 a_34396_15704# a_34308_15748# VPWR.t5963 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X638 a_17036_21976# a_16948_22020# VGND.t2364 VGND.t2363 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X639 VPWR.t3161 a_41340_2727# a_41252_2824# VPWR.t3160 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X640 a_62396_11000# a_62308_11044# VGND.t1834 VGND.t1833 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X641 VPWR.t3775 a_62956_12135# a_62868_12232# VPWR.t3774 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X642 a_51196_14136# a_51108_14180# VGND.t4078 VGND.t2555 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X643 a_31920_29480# a_31508_29159.t2 VGND.t88 VGND.t87 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X644 VPWR.t4767 a_65084_12568# a_64996_12612# VPWR.t4766 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X645 a_52228_19368# _424_.A2.t7 _424_.ZN VGND.t184 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X646 VPWR.t6646 _452_.CLK.t36 a_35092_19368.t0 VPWR.t6645 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X647 a_25524_26344# _351_.A2 a_25300_26344# VPWR.t3255 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X648 a_51196_11000# a_51108_11044# VGND.t1658 VGND.t1657 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X649 VPWR.t3706 a_35068_15271# a_34980_15368# VPWR.t3705 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X650 a_32088_24831# a_30240_24776# a_31803_24831# VPWR.t6319 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X651 a_3260_25112# a_3172_25156# VGND.t5715 VGND.t2588 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X652 VPWR.t3863 a_1468_13703# a_1380_13800# VPWR.t2216 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X653 VGND.t6310 a_54864_22461.t3 a_54824_22045# VGND.t6309 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X654 VGND.t3992 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I VGND.t3991 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X655 VPWR.t1269 _399_.ZN _424_.B1.t1 VPWR.t1268 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X656 VPWR.t2607 a_15132_1592# a_15044_1636# VPWR.t2606 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X657 VPWR.t3263 a_53324_13703# a_53236_13800# VPWR.t3262 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X658 VPWR.t5134 vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I VPWR.t5133 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X659 a_2364_8999# a_2276_9096# VGND.t3933 VGND.t607 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X660 a_35723_20569# a_33748_20936.t2 a_35088_20893# VPWR.t48 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X661 a_60405_31198# a_60285_30600# VPWR.t360 VPWR.t359 pfet_06v0 ad=61.19999f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X662 VPWR.t4186 a_41160_29083# uo_out[3].t2 VPWR.t4185 pfet_06v0 ad=0.428p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
X663 a_3260_21976# a_3172_22020# VGND.t2193 VGND.t2192 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X664 VPWR.t5557 a_39100_1592# a_39012_1636# VPWR.t627 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X665 a_4156_18407# a_4068_18504# VGND.t5158 VGND.t2194 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X666 VGND.t35 _363_.Z.t2 a_32508_30644# VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X667 VGND.t3516 _296_.ZN uo_out[0].t3 VGND.t1138 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X668 VPWR.t3376 a_23868_2727# a_23780_2824# VPWR.t3375 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X669 a_2364_5863# a_2276_5960# VGND.t4070 VGND.t448 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X670 a_30812_18407# a_30724_18504# VGND.t1401 VGND.t1400 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X671 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN VGND.t5335 VGND.t603 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X672 VPWR.t5581 a_61052_9432# a_60964_9476# VPWR.t5580 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X673 a_62844_12568# a_62756_12612# VGND.t2370 VGND.t2369 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X674 VPWR.t3516 a_65532_14136# a_65444_14180# VPWR.t3515 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X675 a_39324_26247# a_39236_26344# VGND.t3821 VGND.t3820 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X676 a_50076_15704# a_49988_15748# VGND.t1397 VGND.t1396 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X677 VPWR.t6068 a_4940_12135# a_4852_12232# VPWR.t6067 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X678 a_51644_12568# a_51556_12612# VGND.t2989 VGND.t2988 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X679 VGND.t4297 a_45088_29123# a_45040_29167# VGND.t4296 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X680 VPWR.t3948 a_65532_11000# a_65444_11044# VPWR.t3947 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X681 VPWR.t3779 a_17596_2727# a_17508_2824# VPWR.t3778 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X682 _284_.B _282_.ZN VPWR.t777 VPWR.t776 pfet_06v0 ad=0.2808p pd=1.6u as=0.5292p ps=3.14u w=1.08u l=0.5u
X683 a_61164_23111# a_61076_23208# VGND.t5295 VGND.t5294 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X684 a_26556_21543# a_26468_21640# VGND.t2967 VGND.t2966 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X685 VPWR.t4227 _470_.Q _397_.A4 VPWR.t4226 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X686 a_53212_14136# a_53124_14180# VGND.t3783 VGND.t3782 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X687 VPWR.t3106 a_1916_12135# a_1828_12232# VPWR.t2698 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X688 a_43580_27815# a_43492_27912# VGND.t3607 VGND.t3606 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X689 _411_.A2.t7 _402_.A1.t8 VPWR.t6721 VPWR.t6720 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X690 a_50524_2727# a_50436_2824# VGND.t6056 VGND.t6055 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X691 a_53076_24776# _398_.C _478_.D VPWR.t3311 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X692 a_53212_11000# a_53124_11044# VGND.t3570 VGND.t3569 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X693 VPWR.t3583 _371_.A2 a_28596_27916.t7 VPWR.t3582 pfet_06v0 ad=0.312p pd=1.72u as=0.528p ps=3.28u w=1.2u l=0.5u
X694 a_52267_30644# a_51791_30644# VGND.t5272 VGND.t45 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X695 VPWR.t1799 a_22748_21543# a_22660_21640# VPWR.t1798 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X696 a_43916_29816# a_43828_29860# VGND.t3323 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X697 VPWR.t4011 a_67548_9432# a_67460_9476# VPWR.t4010 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X698 VPWR.t6255 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN VPWR.t6254 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X699 VGND.t4517 a_54432_31128# _304_.B VGND.t4514 nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X700 a_32604_18840# a_32516_18884# VGND.t5379 VGND.t2582 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X701 a_38616_24328# _437_.A1.t4 VPWR.t6858 VPWR.t6857 pfet_06v0 ad=0.156p pd=1.12u as=0.40575p ps=2.055u w=0.6u l=0.5u
X702 VGND.t6196 _459_.CLK.t19 a_24452_30344.t1 VGND.t139 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X703 a_51540_24776# _412_.B2 VPWR.t5962 VPWR.t5961 pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X704 a_29835_28776# _352_.A2.t17 _370_.ZN VGND.t6666 nfet_06v0 ad=85.2f pd=0.95u as=0.21175p ps=1.41u w=0.71u l=0.6u
X705 a_3260_15704# a_3172_15748# VGND.t4442 VGND.t2080 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X706 a_52136_20936# _424_.A1 _424_.B2 VGND.t304 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X707 VPWR.t3893 a_17932_27815# a_17844_27912# VPWR.t3892 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X708 a_44252_2727# a_44164_2824# VGND.t2974 VGND.t1176 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X709 a_46837_29076# _383_.A2 VGND.t1016 VGND.t1015 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X710 a_51084_12135# a_50996_12232# VGND.t3206 VGND.t3205 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X711 a_47164_10567# a_47076_10664# VGND.t3704 VGND.t3703 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X712 a_13340_29816# a_13252_29860# VGND.t5374 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X713 VPWR.t5238 a_19164_26247# a_19076_26344# VPWR.t5237 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X714 VPWR.t4198 a_63292_2727# a_63204_2824# VPWR.t4197 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X715 VPWR.t1610 a_55340_24679# a_55252_24776# VPWR.t1609 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X716 VPWR.t2073 a_43356_1592# a_43268_1636# VPWR.t2072 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X717 VGND.t6198 _459_.CLK.t20 a_32180_25640.t1 VGND.t6197 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X718 a_4940_27815# a_4852_27912# VGND.t5333 VGND.t5332 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X719 a_6172_29383# a_6084_29480# VGND.t3555 VGND.t3554 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X720 VPWR.t1754 a_67324_1592# a_67236_1636# VPWR.t1753 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X721 VPWR.t1606 a_19164_23111# a_19076_23208# VPWR.t1605 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X722 VGND.t6358 _452_.CLK.t37 a_45284_19751.t1 VGND.t6357 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X723 a_32268_21976# a_32180_22020# VGND.t3636 VGND.t3635 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X724 a_21068_25112# a_20980_25156# VGND.t5377 VGND.t5376 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X725 a_48956_1159# a_48868_1256# VGND.t3160 VGND.t3159 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X726 VPWR.t4017 a_66092_16839# a_66004_16936# VPWR.t4016 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X727 a_1916_27815# a_1828_27912# VGND.t3123 VGND.t1260 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X728 input9.Z a_52639_30644# VPWR.t4138 VPWR.t4137 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X729 a_3708_2727# a_3620_2824# VGND.t2953 VGND.t2952 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X730 a_21068_21976# a_20980_22020# VGND.t3308 VGND.t3307 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X731 VGND.t3955 a_44340_26183# a_43736_25896# VGND.t3954 nfet_06v0 ad=0.142p pd=1.14u as=0.176p ps=1.68u w=0.4u l=0.6u
X732 VPWR.t2290 a_2812_30951# a_2724_31048# VPWR.t2289 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X733 VGND.t6017 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN VGND.t6016 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X734 VPWR.t1475 a_49740_13703# a_49652_13800# VPWR.t1474 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X735 VGND.t4069 _470_.Q _389_.ZN VGND.t4068 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X736 a_51532_13703# a_51444_13800# VGND.t6019 VGND.t6018 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X737 VPWR.t2664 a_2364_29383# a_2276_29480# VPWR.t2663 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X738 uo_out[6].t3 _287_.A2 VGND.t1932 VGND.t1931 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X739 _284_.ZN.t0 _284_.A2.t2 a_42168_25640.t0 VGND.t26 nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X740 _243_.ZN _241_.Z a_58020_27508# VGND.t3413 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X741 _355_.ZN _355_.B VGND.t2858 VGND.t2857 nfet_06v0 ad=0.21175p pd=1.41u as=0.1209p ps=0.985u w=0.465u l=0.6u
X742 VPWR.t3873 a_34448_25597# a_34440_25273# VPWR.t3872 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X743 a_24204_20408# a_24116_20452# VGND.t3695 VGND.t3694 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X744 a_64300_12135# a_64212_12232# VGND.t5327 VGND.t5326 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X745 VPWR.t349 a_46716_13703# a_46628_13800# VPWR.t348 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X746 _324_.B.t2 _305_.A2 a_42168_22504# VGND.t2875 nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X747 a_53744_22851.t0 _474_.CLK.t36 VPWR.t6747 VPWR.t6746 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X748 VPWR.t5522 a_2364_26247# a_2276_26344# VPWR.t4369 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X749 _355_.B _352_.A2.t18 a_28596_26725# VPWR.t6984 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X750 VPWR.t3966 a_2364_23111# a_2276_23208# VPWR.t3965 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X751 VGND.t20 ui_in[1].t0 a_62532_30736# VGND.t4 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X752 a_65756_26247# a_65668_26344# VGND.t3710 VGND.t3709 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X753 a_46492_15704# a_46404_15748# VGND.t3988 VGND.t3987 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X754 a_49404_18407# a_49316_18504# VGND.t3777 VGND.t3776 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X755 VPWR.t5204 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN VPWR.t1428 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X756 a_50816_19369# a_50280_19369# VGND.t1384 VGND.t1383 nfet_06v0 ad=43.2f pd=0.6u as=0.2637p ps=1.825u w=0.36u l=0.6u
X757 a_43804_30951# a_43716_31048# VGND.t6004 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X758 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I VPWR.t311 VPWR.t310 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X759 VPWR.t4803 _474_.Q _218_.ZN VPWR.t4802 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X760 VPWR.t5241 a_58924_14136# a_58836_14180# VPWR.t1781 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X761 a_47531_21258# _421_.A1 _475_.D VGND.t5749 nfet_06v0 ad=85.2f pd=0.95u as=0.21175p ps=1.41u w=0.71u l=0.6u
X762 a_21516_23544# a_21428_23588# VGND.t3559 VGND.t3558 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X763 _427_.ZN _422_.ZN a_52452_21236# VGND.t1910 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X764 a_65756_23111# a_65668_23208# VGND.t3348 VGND.t3347 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X765 a_35292_15704# a_35204_15748# VGND.t3721 VGND.t3720 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X766 a_52988_9432# a_52900_9476# VGND.t3793 VGND.t3792 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X767 a_10876_1159# a_10788_1256# VGND.t3318 VGND.t3317 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X768 a_64860_4295# a_64772_4392# VGND.t2961 VGND.t2960 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X769 a_43814_21236# a_42982_21730# a_43646_21236# VGND.t5257 nfet_06v0 ad=0.369p pd=2.77u as=43.2f ps=0.6u w=0.36u l=0.6u
X770 a_43932_17800# _325_.A1.t7 _325_.ZN VGND.t6513 nfet_06v0 ad=0.1312p pd=1.14u as=0.2569p ps=1.56u w=0.82u l=0.6u
X771 VPWR.t13 _397_.A1.t2 a_50308_26476# VPWR.t12 pfet_06v0 ad=0.4005p pd=2.12u as=0.1456p ps=1.08u w=0.56u l=0.5u
X772 VPWR.t1612 a_63516_15271# a_63428_15368# VPWR.t1611 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X773 VPWR.t3719 a_40444_15704# a_40356_15748# VPWR.t3718 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X774 VGND.t3358 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I _241_.I0 VGND.t3357 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X775 a_66876_15271# a_66788_15368# VGND.t2985 VGND.t879 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X776 a_59036_12568# a_58948_12612# VGND.t3871 VGND.t3870 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X777 a_46128_20127# a_45696_20072# VPWR.t2599 VPWR.t2598 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X778 a_42728_20452# _452_.Q.t5 a_42460_20452# VPWR.t6949 pfet_06v0 ad=0.33945p pd=1.715u as=0.4599p ps=1.935u w=1.095u l=0.5u
X779 a_30588_21543# a_30500_21640# VGND.t3697 VGND.t3696 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X780 VPWR.t3541 a_1020_19975# a_932_20072# VPWR.t3540 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X781 VGND.t3470 _260_.ZN a_43245_24373# VGND.t3469 nfet_06v0 ad=0.341p pd=2.43u as=92.99999f ps=1.015u w=0.775u l=0.6u
X782 _475_.Q a_47776_20893# VGND.t1808 VGND.t1807 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X783 VPWR.t1416 a_41116_15271# a_41028_15368# VPWR.t1415 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X784 a_44476_15271# a_44388_15368# VGND.t3906 VGND.t3905 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X785 a_45664_26031# a_45128_26031# VGND.t2515 VGND.t2514 nfet_06v0 ad=43.2f pd=0.6u as=0.2637p ps=1.825u w=0.36u l=0.6u
X786 _261_.ZN _447_.Q.t4 a_39796_22504# VGND.t2813 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X787 a_58687_31220# a_58063_30644# a_58519_31220# VPWR.t3241 pfet_06v0 ad=0.3852p pd=2.86u as=61.19999f ps=0.7u w=0.36u l=0.5u
X788 VPWR.t6325 a_50524_17272# a_50436_17316# VPWR.t6324 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X789 VGND.t4869 a_20672_30301# a_20624_30345# VGND.t137 nfet_06v0 ad=0.2333p pd=1.555u as=43.2f ps=0.6u w=0.36u l=0.6u
X790 a_22064_27912# a_21652_27591.t3 VPWR.t103 VPWR.t102 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X791 _359_.ZN _358_.A3 a_34308_26344# VPWR.t479 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X792 VGND.t2181 a_6723_30644# a_6723_30644# VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X793 a_17484_25112# a_17396_25156# VGND.t1409 VGND.t1408 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X794 VPWR.t3777 a_54780_20408# a_54692_20452# VPWR.t3776 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X795 a_42252_20936# _304_.B VGND.t4541 VGND.t4540 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X796 VPWR.t4241 a_21852_2727# a_21764_2824# VPWR.t4240 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X797 VPWR.t6285 a_9980_29383# a_9892_29480# VPWR.t6284 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X798 a_4156_7864# a_4068_7908# VGND.t3106 VGND.t3031 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X799 a_18096_27165# a_17803_26841# VGND.t1271 VGND.t1270 nfet_06v0 ad=0.2119p pd=1.335u as=0.2333p ps=1.555u w=0.815u l=0.6u
X800 a_17484_21976# a_17396_22020# VGND.t1614 VGND.t1613 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X801 a_25884_1592# a_25796_1636# VGND.t6054 VGND.t6053 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X802 a_51868_1159# a_51780_1256# VGND.t2484 VGND.t2483 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X803 _335_.ZN.t16 _459_.Q.t3 VPWR.t6965 VPWR.t6964 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X804 a_2812_1592# a_2724_1636# VGND.t3564 VGND.t1220 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X805 a_43356_1159# a_43268_1256# VGND.t2531 VGND.t2530 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X806 VPWR.t3500 a_23196_23111# a_23108_23208# VPWR.t3499 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X807 a_4156_4728# a_4068_4772# VGND.t1376 VGND.t1375 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X808 a_21404_24679# a_21316_24776# VGND.t3797 VGND.t3796 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X809 a_49852_1592# a_49764_1636# VGND.t3322 VGND.t3321 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X810 VPWR.t3185 a_64972_13703# a_64884_13800# VPWR.t3184 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X811 a_35180_16839# a_35092_16936# VGND.t1942 VGND.t1941 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X812 a_39968_26841# a_39536_26795# VPWR.t3266 VPWR.t3265 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X813 VPWR.t5518 a_15580_2727# a_15492_2824# VPWR.t5517 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X814 VGND.t900 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN VGND.t899 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X815 VPWR.t3125 a_43916_29816# a_43828_29860# VPWR.t3124 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X816 a_34084_28776# _362_.B.t5 a_37324_28776# VGND.t6250 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X817 VGND.t3961 a_43736_25896# _402_.A1.t3 VGND.t3960 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X818 a_21404_21543# a_21316_21640# VGND.t3407 VGND.t3406 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X819 VPWR.t4032 a_53772_13703# a_53684_13800# VPWR.t4031 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X820 a_32156_16839# a_32068_16936# VGND.t4011 VGND.t2877 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X821 a_55228_28248# a_55140_28292# VGND.t5697 VGND.t5696 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X822 a_48272_25156.t7 clkbuf_1_0__f_clk.I.t33 VPWR.t244 VPWR.t243 pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X823 a_67548_4295# a_67460_4392# VGND.t3700 VGND.t3523 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X824 VPWR.t3865 a_33052_19975# a_32964_20072# VPWR.t3864 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X825 VPWR.t5573 a_13340_29816# a_13252_29860# VPWR.t5572 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X826 a_17932_23544# a_17844_23588# VGND.t2368 VGND.t2367 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X827 VPWR.t1616 a_66204_7431# a_66116_7528# VPWR.t1615 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X828 VGND.t916 _384_.A1 _384_.ZN VGND.t915 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X829 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN VPWR.t1732 VPWR.t1731 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X830 a_47924_28292# _381_.Z a_47700_28292# VPWR.t3950 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X831 VPWR.t1774 a_65980_14136# a_65892_14180# VPWR.t1773 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X832 VPWR.t228 _304_.ZN.t11 _324_.B.t19 VPWR.t227 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X833 a_39772_26247# a_39684_26344# VGND.t3996 VGND.t3995 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X834 _427_.B2 _281_.A1 VPWR.t3302 VPWR.t3301 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X835 VPWR.t3380 a_66316_10567# a_66228_10664# VPWR.t3379 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X836 a_47636_25940# _282_.ZN VGND.t760 VGND.t759 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X837 a_17820_30951# a_17732_31048# VGND.t2949 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X838 _454_.Q a_23920_27555# VGND.t612 VGND.t611 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X839 VPWR.t3452 a_65980_11000# a_65892_11044# VPWR.t3451 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X840 a_49628_17272# a_49540_17316# VGND.t5724 VGND.t5723 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X841 VPWR.t5560 a_1916_20408# a_1828_20452# VPWR.t1141 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X842 _313_.ZN _330_.A1.t5 a_36288_23208# VPWR.t207 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X843 a_22076_1592# a_21988_1636# VGND.t1616 VGND.t1615 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X844 _371_.A2 _455_.Q.t3 VPWR.t6847 VPWR.t6846 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X845 VPWR.t5184 a_47164_18407# a_47076_18504# VPWR.t5183 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X846 VPWR.t1275 a_55116_10567# a_55028_10664# VPWR.t1274 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X847 a_47948_23111# a_47860_23208# VGND.t3405 VGND.t3404 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X848 a_59332_29816# _324_.C.t10 VPWR.t6794 VPWR.t6793 pfet_06v0 ad=0.2354p pd=1.95u as=0.1391p ps=1.055u w=0.535u l=0.5u
X849 a_1916_7431# a_1828_7528# VGND.t1 VGND.t0 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X850 a_53660_14136# a_53572_14180# VGND.t5604 VGND.t375 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X851 VPWR.t4853 a_48732_15271# a_48644_15368# VPWR.t4852 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X852 a_46044_1592# a_45956_1636# VGND.t4707 VGND.t638 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X853 a_44864_27165# a_44571_26841# VPWR.t2960 VPWR.t2959 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X854 a_53796_30344# vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN a_53592_30344# VGND.t3612 nfet_06v0 ad=88.2f pd=0.84u as=88.2f ps=0.84u w=0.42u l=0.6u
X855 a_54432_31128# ui_in[7].t0 VPWR.t9 VPWR.t8 pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X856 a_53660_11000# a_53572_11044# VGND.t534 VGND.t533 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X857 VGND.t538 vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN VGND.t537 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X858 a_1020_29383# a_932_29480# VGND.t5322 VGND.t686 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X859 a_45577_27509# _404_.A1 _470_.D VGND.t3676 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X860 a_35756_27216# _460_.Q a_35552_27216# VGND.t3336 nfet_06v0 ad=60.8f pd=0.7u as=79.8f ps=0.8u w=0.38u l=0.6u
X861 VPWR.t1858 a_1468_12568# a_1380_12612# VPWR.t1857 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X862 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I VPWR.t1864 VPWR.t1863 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X863 a_24764_2727# a_24676_2824# VGND.t2444 VGND.t2443 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X864 clkbuf_1_0__f_clk.I.t12 a_44296_24393.t18 VPWR.t242 VPWR.t241 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X865 VGND.t5844 a_17168_27165# a_17120_27209# VGND.t5843 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X866 VPWR.t6648 _452_.CLK.t38 a_36548_27591.t0 VPWR.t6647 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X867 VPWR.t6104 a_46940_17272# a_46852_17316# VPWR.t6103 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X868 VGND.t1405 _399_.A2 a_49405_22805# VGND.t1404 nfet_06v0 ad=0.341p pd=2.43u as=92.99999f ps=1.015u w=0.775u l=0.6u
X869 vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN VPWR.t2603 VPWR.t2602 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X870 VPWR.t4289 a_48508_2727# a_48420_2824# VPWR.t4288 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X871 VPWR.t4290 a_23868_1592# a_23780_1636# VPWR.t2972 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X872 VPWR.t1483 a_35740_17272# a_35652_17316# VPWR.t1482 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X873 a_14684_1159# a_14596_1256# VGND.t1419 VGND.t1418 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X874 VGND.t1069 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN VGND.t1068 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X875 VPWR.t1826 a_62396_27815# a_62308_27912# VPWR.t1825 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X876 a_18492_2727# a_18404_2824# VGND.t5100 VGND.t1120 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X877 a_38288_18191# a_37408_18504# a_37964_18191# VGND.t1754 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X878 VPWR.t2565 a_1468_8999# a_1380_9096# VPWR.t2564 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X879 VPWR.t2566 a_60828_1159# a_60740_1256# VPWR.t1771 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X880 VPWR.t1685 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t1684 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X881 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t1868 VPWR.t1867 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X882 VPWR.t1693 _495_.I a_41160_29083# VPWR.t1692 pfet_06v0 ad=0.3608p pd=2.52u as=0.2542p ps=1.44u w=0.82u l=0.5u
X883 VPWR.t2623 a_16588_26247# a_16500_26344# VPWR.t2622 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X884 VPWR.t2625 a_17596_1592# a_17508_1636# VPWR.t2624 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X885 _303_.ZN _325_.A1.t8 VPWR.t6820 VPWR.t6819 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X886 a_60604_26247# a_60516_26344# VGND.t706 VGND.t705 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X887 VPWR.t4317 a_1916_14136# a_1828_14180# VPWR.t1290 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X888 a_41340_15704# a_41252_15748# VGND.t4156 VGND.t4155 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X889 a_47948_16839# a_47860_16936# VGND.t1560 VGND.t1559 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X890 VPWR.t1644 a_16588_23111# a_16500_23208# VPWR.t1643 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X891 VPWR.t1920 a_4156_7864# a_4068_7908# VPWR.t742 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X892 a_5052_12568# a_4964_12612# VGND.t1695 VGND.t1694 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X893 VPWR.t1786 a_41564_24679# a_41476_24776# VPWR.t1785 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X894 VPWR.t1801 a_1916_11000# a_1828_11044# VPWR.t1800 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X895 a_50972_9432# a_50884_9476# VGND.t1711 VGND.t1710 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X896 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I _274_.A1 VGND.t2525 VGND.t2524 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X897 a_51980_13703# a_51892_13800# VGND.t2527 VGND.t2526 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X898 a_62503_28293# _250_.B a_62279_28293# VPWR.t2507 pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X899 VGND.t2385 _242_.Z a_58020_27508# VGND.t2384 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X900 a_24652_20408# a_24564_20452# VGND.t1792 VGND.t1791 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X901 VGND.t2420 hold2.I a_43192_25640# VGND.t2419 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X902 a_66652_3160# a_66564_3204# VGND.t1794 VGND.t1793 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X903 a_58028_20408# a_57940_20452# VGND.t2387 VGND.t2386 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X904 VPWR.t7 ui_in[2].t0 a_61860_30736# VPWR.t6 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X905 a_61724_15271# a_61636_15368# VGND.t5458 VGND.t5457 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X906 VGND.t237 _304_.ZN.t12 a_43192_22504# VGND.t236 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X907 _452_.D _332_.Z VGND.t4890 VGND.t4889 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X908 a_18352_28777# a_17472_28363# a_18028_28777# VGND.t2504 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X909 a_51084_28248# a_50996_28292# VGND.t5037 VGND.t5036 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X910 a_51540_23588# _417_.A2.t3 VPWR.t130 VPWR.t129 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X911 VPWR.t5203 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN VPWR.t1426 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X912 VGND.t3027 a_35140_26680# _363_.Z.t1 VGND.t3026 nfet_06v0 ad=0.2424p pd=1.635u as=0.341p ps=2.43u w=0.775u l=0.6u
X913 _399_.ZN _399_.A1 a_48321_23208# VPWR.t4237 pfet_06v0 ad=0.3159p pd=1.735u as=0.32805p ps=1.755u w=1.215u l=0.5u
X914 _438_.ZN _438_.A2 VPWR.t5121 VPWR.t5120 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X915 a_21964_23544# a_21876_23588# VGND.t2406 VGND.t2405 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X916 VPWR.t2534 a_55340_23544# a_55252_23588# VPWR.t2533 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X917 a_55676_1159# a_55588_1256# VGND.t2034 VGND.t2033 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X918 a_56684_17272# a_56596_17316# VGND.t2036 VGND.t2035 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X919 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I VGND.t2965 VGND.t2964 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X920 a_47164_1159# a_47076_1256# VGND.t4240 VGND.t4239 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X921 VPWR.t4611 a_53212_27815# a_53124_27912# VPWR.t4610 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X922 _350_.A2.t9 _371_.A1.t10 a_30388_28776# VGND.t6231 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X923 a_45169_27509# _330_.A1.t6 VGND.t209 VGND.t208 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X924 VPWR.t5275 a_63964_15271# a_63876_15368# VPWR.t5274 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X925 a_35628_18407# a_35540_18504# VGND.t5110 VGND.t5109 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X926 _337_.ZN _336_.A1 VPWR.t4212 VPWR.t4211 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X927 a_35710_28776# _460_.Q a_35516_28776# VGND.t3335 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X928 VPWR.t6127 a_48508_10567# a_48420_10664# VPWR.t4725 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X929 VPWR.t2434 a_40892_15704# a_40804_15748# VPWR.t2433 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X930 VPWR.t2440 a_48104_30219# _397_.A2.t1 VPWR.t2439 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X931 a_59484_12568# a_59396_12612# VGND.t4717 VGND.t4716 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X932 VGND.t4222 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I _248_.B1 VGND.t4221 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X933 VPWR.t4863 a_63068_18840# a_62980_18884# VPWR.t4066 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X934 a_23532_21976# a_23444_22020# VGND.t1571 VGND.t1570 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X935 VPWR.t6670 _355_.C.t5 _346_.B VPWR.t6669 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X936 a_32476_29167# _461_.D a_32352_29535# VPWR.t851 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X937 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].I VGND.t5049 VGND.t5048 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X938 VPWR.t2677 a_63068_15704# a_62980_15748# VPWR.t2676 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X939 VPWR.t2643 a_2364_28248# a_2276_28292# VPWR.t2642 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X940 VPWR.t2645 a_41564_15271# a_41476_15368# VPWR.t2644 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X941 VPWR.t6951 _452_.Q.t6 _441_.A3 VPWR.t6950 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X942 _242_.Z a_56516_26344# VPWR.t337 VPWR.t336 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X943 VPWR.t1766 a_60380_12568# a_60292_12612# VPWR.t1765 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X944 a_49604_22020# _384_.A1 _384_.ZN VPWR.t939 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X945 VPWR.t2528 a_46716_12568# a_46628_12612# VPWR.t2527 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X946 a_35232_24029# a_34939_23705# VPWR.t688 VPWR.t687 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X947 VPWR.t5676 a_2364_25112# a_2276_25156# VPWR.t620 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X948 VPWR.t4836 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_57168_26724# VPWR.t4835 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X949 VGND.t6651 _459_.Q.t4 _358_.A2 VGND.t6650 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X950 VGND.t4539 _304_.B _386_.ZN VGND.t4538 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X951 a_28124_26680# a_28036_26724# VGND.t1786 VGND.t1785 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X952 VPWR.t1885 a_51308_16839# a_51220_16936# VPWR.t1884 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X953 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I VGND.t508 VGND.t507 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X954 a_1468_1159# a_1380_1256# VGND.t3488 VGND.t3487 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X955 VPWR.t1502 a_50972_17272# a_50884_17316# VPWR.t1501 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X956 VPWR.t1504 a_40108_16839# a_40020_16936# VPWR.t1503 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X957 VGND.t6239 _284_.ZN.t23 uo_out[0].t11 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X958 VPWR.t2666 a_5052_18840# a_4964_18884# VPWR.t2665 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X959 VPWR.t1722 a_64412_18407# a_64324_18504# VPWR.t1721 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X960 a_50300_1592# a_50212_1636# VGND.t1646 VGND.t1645 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X961 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN VGND.t5911 VGND.t5910 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X962 VPWR.t6217 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN a_53212_29816# VPWR.t6216 pfet_06v0 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X963 a_59796_29480# _238_.ZN _258_.I VPWR.t6178 pfet_06v0 ad=0.3172p pd=1.74u as=0.4016p ps=1.94u w=1.22u l=0.5u
X964 _371_.A2 _349_.A4 VPWR.t2563 VPWR.t2562 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X965 a_53380_20127# _424_.ZN a_52512_19715# VPWR.t5977 pfet_06v0 ad=54f pd=0.66u as=0.1872p ps=1.4u w=0.36u l=0.5u
X966 a_21852_24679# a_21764_24776# VGND.t2486 VGND.t2485 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X967 VPWR.t2617 a_5052_15704# a_4964_15748# VPWR.t2616 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X968 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I VGND.t1429 VGND.t1428 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X969 a_31708_15704# a_31620_15748# VGND.t1431 VGND.t1430 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X970 a_50644_21640# _218_.ZN _474_.D VPWR.t3771 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X971 a_21852_21543# a_21764_21640# VGND.t2539 VGND.t2538 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X972 VGND.t2463 a_16916_31048# uio_oe[0].t0 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X973 a_61836_25515# a_62560_25112# a_62404_25156# VPWR.t2592 pfet_06v0 ad=0.3172p pd=1.74u as=0.4758p ps=2u w=1.22u l=0.5u
X974 a_23420_26247# a_23332_26344# VGND.t5836 VGND.t5835 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X975 a_30596_28292# _337_.ZN VPWR.t5141 VPWR.t5140 pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X976 a_23912_27967# a_22064_27912# a_23627_27967# VPWR.t3413 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X977 a_55676_28248# a_55588_28292# VGND.t2395 VGND.t2394 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X978 a_46940_15271# a_46852_15368# VGND.t2397 VGND.t2396 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X979 a_59372_13703# a_59284_13800# VGND.t4143 VGND.t4142 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X980 a_18492_1159# a_18404_1256# VGND.t4145 VGND.t4144 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X981 _438_.ZN _451_.Q.t2 VPWR.t6419 VPWR.t6418 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X982 a_41776_20072# _328_.A2 a_41572_20072# VPWR.t5665 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X983 a_42853_24373# _260_.ZN VGND.t3468 VGND.t3467 nfet_06v0 ad=92.99999f pd=1.015u as=0.23975p ps=1.475u w=0.775u l=0.6u
X984 VGND.t6145 a_52064_19715.t2 a_53436_19759# VGND.t6144 nfet_06v0 ad=0.1584p pd=1.6u as=43.2f ps=0.6u w=0.36u l=0.6u
X985 VPWR.t4882 _340_.A2 a_25962_29480# VPWR.t4881 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X986 a_1020_8999# a_932_9096# VGND.t4733 VGND.t475 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X987 a_32828_1592# a_32740_1636# VGND.t1625 VGND.t1624 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X988 VPWR.t1705 a_7628_30951# a_7540_31048# VPWR.t1704 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X989 VGND.t103 _294_.A2.t3 _287_.A2 VGND.t102 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X990 a_34348_27208# _334_.A1 _371_.A1.t2 VGND.t2246 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X991 a_64412_29816# a_64324_29860# VGND.t1617 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X992 a_61052_27815# a_60964_27912# VGND.t5460 VGND.t5459 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X993 VPWR.t5663 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t5662 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X994 _337_.ZN _337_.A3.t2 VPWR.t6401 VPWR.t6400 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X995 a_51457_29861# _276_.A2 vgaringosc.workerclkbuff_notouch_.I.t3 VPWR.t2573 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X996 _275_.ZN _416_.A1.t4 VGND.t196 VGND.t195 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X997 a_1020_5863# a_932_5960# VGND.t2482 VGND.t1406 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X998 VPWR.t5669 a_66764_10567# a_66676_10664# VPWR.t5668 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X999 a_21287_29076# _375_.Z a_21103_29076# VGND.t5470 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1000 VPWR.t2536 a_66988_18407# a_66900_18504# VPWR.t2535 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1001 VGND.t5382 a_53212_29816# _274_.A1 VGND.t199 nfet_06v0 ad=0.226p pd=1.515u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1002 VPWR.t1664 a_36860_23111# a_36772_23208# VPWR.t1663 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1003 a_37179_24831# a_35616_24776# a_36544_24419# VGND.t1588 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1004 VPWR.t5261 a_22636_29383# a_22548_29480# VPWR.t5260 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1005 VPWR.t3536 a_33776_29123# _362_.B.t1 VPWR.t3535 pfet_06v0 ad=0.854p pd=3.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1006 _404_.A1 _470_.Q VPWR.t4225 VPWR.t4224 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1007 VGND.t2458 _379_.Z _467_.D VGND.t2457 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1008 VPWR.t2589 a_59036_26247# a_58948_26344# VPWR.t2588 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1009 VPWR.t1679 a_55564_10567# a_55476_10664# VPWR.t1678 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1010 a_50636_10567# a_50548_10664# VGND.t1600 VGND.t1599 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1011 a_62172_19975# a_62084_20072# VGND.t5467 VGND.t5150 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1012 _234_.ZN _436_.B VGND.t5646 VGND.t5645 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1013 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I VGND.t898 VGND.t897 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1014 VPWR.t5651 a_16252_2727# a_16164_2824# VPWR.t5650 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1015 a_45088_29123# a_44795_29535# VGND.t5293 VGND.t5292 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X1016 a_51240_20452# _419_.Z VGND.t4313 VGND.t4312 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1017 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN VPWR.t1740 VPWR.t1739 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1018 VGND.t4564 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I VGND.t4563 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1019 a_42784_25640# hold2.I VGND.t2418 VGND.t2417 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1020 VGND.t6638 _452_.Q.t7 a_42154_21236# VGND.t6637 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1021 VPWR.t209 _330_.A1.t7 a_38506_26724# VPWR.t208 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1022 VPWR.t1630 a_15580_1592# a_15492_1636# VPWR.t1629 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1023 VPWR.t1632 a_48284_15704# a_48196_15748# VPWR.t1631 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1024 a_14796_26247# a_14708_26344# VGND.t5480 VGND.t2217 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1025 VPWR.t5682 a_31820_20408# a_31732_20452# VPWR.t5681 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1026 clkload0.Z a_48384_26724# VGND.t2868 VGND.t2867 nfet_06v0 ad=0.1183p pd=0.975u as=0.2002p ps=1.79u w=0.455u l=0.6u
X1027 a_42784_22504# _304_.ZN.t13 VGND.t239 VGND.t238 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1028 a_63105_28293# vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN _250_.A2 VPWR.t4282 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1029 clkbuf_1_0__f_clk.I.t11 a_44296_24393.t19 VPWR.t276 VPWR.t275 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1030 a_67100_7431# a_67012_7528# VGND.t5477 VGND.t1116 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1031 a_65084_14136# a_64996_14180# VGND.t5479 VGND.t5478 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1032 VPWR.t3885 a_37084_15704# a_36996_15748# VPWR.t3884 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1033 VPWR.t3887 a_61948_12568# a_61860_12612# VPWR.t3886 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1034 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t1012 VGND.t1011 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1035 VPWR.t6298 a_44744_26355# a_46100_26399# VPWR.t6297 pfet_06v0 ad=0.4554p pd=3.25u as=54f ps=0.66u w=0.36u l=0.5u
X1036 a_14796_23111# a_14708_23208# VGND.t6033 VGND.t3977 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1037 a_22059_26399# a_20496_26344# a_21424_25987# VGND.t4670 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1038 VPWR.t5987 a_66204_9432# a_66116_9476# VPWR.t883 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1039 a_39268_18840# _451_.Q.t3 VPWR.t6421 VPWR.t6420 pfet_06v0 ad=0.1456p pd=1.08u as=0.34437p ps=1.895u w=0.56u l=0.5u
X1040 VPWR.t2038 a_27004_1159# a_26916_1256# VPWR.t2037 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1041 VPWR.t3715 a_36524_16839# a_36436_16936# VPWR.t3714 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1042 VGND.t457 a_46624_19715# a_46576_19759# VGND.t456 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X1043 a_34080_22461# a_33708_22505# VPWR.t3717 VPWR.t3716 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X1044 a_65084_11000# a_64996_11044# VGND.t1958 VGND.t1957 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1045 a_59484_1159# a_59396_1256# VGND.t1960 VGND.t1959 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1046 a_67996_1159# a_67908_1256# VGND.t4342 VGND.t4341 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1047 VPWR.t4491 a_50748_12568# a_50660_12612# VPWR.t4490 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1048 VPWR.t6600 _304_.A1.t5 a_39178_23208# VPWR.t6599 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1049 VGND.t3486 _346_.A2 _454_.D VGND.t3485 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X1050 VPWR.t4907 a_67212_13703# a_67124_13800# VPWR.t4906 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1051 _428_.Z a_51240_23340# VPWR.t441 VPWR.t440 pfet_06v0 ad=0.5368p pd=3.32u as=0.389p ps=2.02u w=1.22u l=0.5u
X1052 _371_.A2 _454_.Q VPWR.t4092 VPWR.t4091 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X1053 VPWR.t5207 a_4156_13703# a_4068_13800# VPWR.t3052 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1054 a_58709_29076# _246_.B2 VGND.t5057 VGND.t5056 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1055 VPWR.t2268 a_42012_1592# a_41924_1636# VPWR.t2267 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1056 VPWR.t2270 a_56012_13703# a_55924_13800# VPWR.t2269 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1057 a_21103_29076# _379_.A2 VGND.t2601 VGND.t2600 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1058 a_52408_19759# a_52024_20083# a_51620_19911# VGND.t427 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1059 a_43444_19668# _324_.C.t11 VGND.t6501 VGND.t6500 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1060 a_50972_2727# a_50884_2824# VGND.t2615 VGND.t2614 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1061 a_27004_1159# a_26916_1256# VGND.t1936 VGND.t1935 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1062 a_33500_18407# a_33412_18504# VGND.t2616 VGND.t976 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1063 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN VPWR.t5826 VPWR.t5825 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1064 VGND.t3382 a_33776_29123# a_33728_29167# VGND.t3381 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X1065 a_65532_12568# a_65444_12612# VGND.t2651 VGND.t2650 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1066 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I VGND.t2099 VGND.t2098 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1067 VPWR.t2211 a_5724_1159# a_5636_1256# VPWR.t2210 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1068 vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t2226 VPWR.t2225 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1069 VPWR.t4090 _454_.Q a_24392_28248# VPWR.t4089 pfet_06v0 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X1070 a_49404_2727# a_49316_2824# VGND.t1868 VGND.t1867 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1071 a_58476_20408# a_58388_20452# VGND.t1870 VGND.t1869 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1072 a_47636_23588# _281_.ZN.t5 a_47412_23588# VPWR.t122 pfet_06v0 ad=0.1736p pd=1.18u as=0.1736p ps=1.18u w=0.56u l=0.5u
X1073 VGND.t6360 _452_.CLK.t39 a_35204_24455.t1 VGND.t6359 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1074 VPWR.t1406 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I VPWR.t1405 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1075 a_5276_1159# a_5188_1256# VGND.t1328 VGND.t1327 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1076 VPWR.t2374 a_39100_15704# a_39012_15748# VPWR.t2373 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1077 VPWR.t246 clkbuf_1_0__f_clk.I.t34 a_42392_22825.t7 VPWR.t245 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1078 a_1468_1592# a_1380_1636# VGND.t1293 VGND.t1292 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1079 vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN VGND.t1297 VGND.t1296 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1080 a_29244_21543# a_29156_21640# VGND.t1299 VGND.t1298 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1081 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _275_.A2 VPWR.t2771 VPWR.t2770 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1082 a_5948_29816# a_5860_29860# VGND.t2633 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1083 VPWR.t2195 a_48508_1592# a_48420_1636# VPWR.t2194 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1084 VPWR.t2197 a_36636_21543# a_36548_21640# VPWR.t2196 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1085 VPWR.t2199 a_67772_1592# a_67684_1636# VPWR.t2198 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1086 a_55788_23544# a_55700_23588# VGND.t2075 VGND.t2074 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1087 VPWR.t2178 a_16588_28248# a_16500_28292# VPWR.t633 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1088 VGND.t4318 _416_.A3 _416_.ZN VGND.t4317 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X1089 VPWR.t4469 a_53660_27815# a_53572_27912# VPWR.t4468 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1090 VPWR.t1891 a_25436_21543# a_25348_21640# VPWR.t1890 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1091 a_42376_25640# _284_.B a_42168_25640.t10 VGND.t5393 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1092 a_24080_25227# a_23668_25640.t2 VGND.t6707 VGND.t6706 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1093 VPWR.t2686 a_55228_1159# a_55140_1256# VPWR.t2685 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1094 VPWR.t2687 a_16588_25112# a_16500_25156# VPWR.t1237 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1095 a_20884_26031# a_20084_26023.t2 VGND.t6681 VGND.t6680 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1096 a_42376_22504# _302_.Z a_42168_22504# VGND.t4846 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1097 a_23980_21976# a_23892_22020# VGND.t2585 VGND.t2584 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1098 VGND.t2785 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN VGND.t2784 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1099 a_28364_28776# _337_.A3.t3 _371_.A2 VGND.t6134 nfet_06v0 ad=0.1312p pd=1.14u as=0.4161p ps=1.905u w=0.82u l=0.6u
X1100 a_46156_25112# a_46068_25156# VGND.t2787 VGND.t2786 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1101 a_44484_19668# _325_.A2.t2 VGND.t6121 VGND.t6120 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1102 a_58028_10567# a_57940_10664# VGND.t2148 VGND.t2147 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1103 VPWR.t1828 a_19724_23544# a_19636_23588# VPWR.t1827 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1104 a_45372_9432# a_45284_9476# VGND.t1740 VGND.t339 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1105 uo_out[2].t6 _287_.A1.t12 VGND.t6481 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1106 VGND.t5507 a_27172_24328# a_26548_24372# VGND.t5506 nfet_06v0 ad=0.218p pd=1.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1107 a_59348_29076# _267_.A2 VGND.t3615 VGND.t3614 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1108 VPWR.t2274 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I VPWR.t2273 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1109 VPWR.t2701 a_51756_16839# a_51668_16936# VPWR.t2700 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1110 VGND.t2572 _319_.A3 _319_.ZN VGND.t2571 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X1111 VPWR.t5657 a_64412_29816# a_64324_29860# VPWR.t5656 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1112 VPWR.t2755 a_3260_6296# a_3172_6340# VPWR.t2754 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1113 a_65420_13703# a_65332_13800# VGND.t2623 VGND.t2622 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1114 a_28000_29480# a_27588_29159.t3 VGND.t6557 VGND.t6556 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1115 a_2364_13703# a_2276_13800# VGND.t1840 VGND.t1839 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1116 a_30112_30345# a_29232_29931# a_29788_30345# VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X1117 a_62396_1159# a_62308_1256# VGND.t1962 VGND.t1961 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1118 VPWR.t2065 a_40556_16839# a_40468_16936# VPWR.t2064 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1119 VPWR.t3245 a_28012_20408# a_27924_20452# VPWR.t3244 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1120 a_54220_13703# a_54132_13800# VGND.t3093 VGND.t3092 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1121 VPWR.t5585 a_53212_29816# _274_.A1 VPWR.t5584 pfet_06v0 ad=0.395p pd=2.02u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1122 VPWR.t3440 a_3260_3160# a_3172_3204# VPWR.t1243 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1123 a_30812_1592# a_30724_1636# VGND.t3296 VGND.t2229 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1124 VGND.t3515 _296_.ZN uo_out[0].t2 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1125 VPWR.t2248 a_64860_18407# a_64772_18504# VPWR.t2247 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1126 VGND.t6469 _359_.B.t5 _370_.ZN VGND.t6468 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X1127 VPWR.t1170 _251_.ZN a_60013_26344# VPWR.t1169 pfet_06v0 ad=0.5346p pd=3.31u as=0.37665p ps=1.835u w=1.215u l=0.5u
X1128 a_38336_18147# a_37964_18191# VGND.t4226 VGND.t4225 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X1129 VGND.t4657 _474_.Q _218_.ZN VGND.t4656 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1130 a_45040_29167# a_42820_29159.t4 a_44795_29535# VGND nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1131 VPWR.t2230 a_61612_10567# a_61524_10664# VPWR.t2229 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1132 a_24540_1592# a_24452_1636# VGND.t1713 VGND.t1712 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1133 a_49180_15704# a_49092_15748# VGND.t1715 VGND.t1714 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1134 a_37352_19001# a_35504_18955# a_37067_19001# VPWR.t1330 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X1135 a_5388_26247# a_5300_26344# VGND.t1267 VGND.t1266 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1136 VPWR.t2850 a_4940_16839# a_4852_16936# VPWR.t2849 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1137 _412_.B2 _397_.A1.t3 a_50792_26344# VPWR.t14 pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1138 VPWR.t2852 a_54332_18840# a_54244_18884# VPWR.t2851 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1139 a_5388_23111# a_5300_23208# VGND.t4545 VGND.t4544 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1140 VPWR.t4705 a_54332_15704# a_54244_15748# VPWR.t4704 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1141 VPWR.t2962 a_1916_16839# a_1828_16936# VPWR.t2961 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1142 VPWR.t2964 a_31260_18407# a_31172_18504# VPWR.t2963 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1143 VPWR.t4210 _336_.A1 a_28596_26725# VPWR.t4209 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X1144 VGND.t6411 vgaringosc.workerclkbuff_notouch_.I.t6 a_41048_29816.t5 VGND.t6409 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1145 VGND.t5422 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN VGND.t5421 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1146 a_66204_4295# a_66116_4392# VGND.t2641 VGND.t2640 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1147 VPWR.t2219 a_61052_14136# a_60964_14180# VPWR.t2218 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1148 VPWR.t2220 a_43132_15704# a_43044_15748# VPWR.t450 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1149 VGND.t6192 a_43440_19325.t3 a_44812_19369# VGND.t6191 nfet_06v0 ad=0.1584p pd=1.6u as=43.2f ps=0.6u w=0.36u l=0.6u
X1150 a_33276_21543# a_33188_21640# VGND.t5068 VGND.t5067 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1151 VPWR.t5224 a_55004_15271# a_54916_15368# VPWR.t5223 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1152 VPWR.t6056 a_61052_11000# a_60964_11044# VPWR.t6055 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1153 vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t5805 VGND.t1194 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1154 a_18400_28733# a_18028_28777# VGND.t2506 VGND.t2505 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X1155 _395_.A1 _404_.A1 VPWR.t3828 VPWR.t3827 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1156 _478_.D _428_.Z VPWR.t4909 VPWR.t4908 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1157 VPWR.t5610 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN VPWR.t5609 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1158 VPWR.t1889 a_64412_17272# a_64324_17316# VPWR.t1888 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1159 a_47164_12135# a_47076_12232# VGND.t2928 VGND.t2927 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1160 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I VGND.t3825 VGND.t3824 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1161 VPWR.t798 _223_.ZN _350_.A2.t2 VPWR.t797 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1162 VPWR.t2173 a_53212_17272# a_53124_17316# VPWR.t2172 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1163 VPWR.t1207 _290_.ZN a_34404_31048# VPWR.t1206 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1164 a_48596_28292# _397_.A1.t4 _383_.ZN VPWR.t15 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1165 a_9084_1159# a_8996_1256# VGND.t2547 VGND.t2546 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1166 VPWR.t2684 a_37084_26247# a_36996_26344# VPWR.t397 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1167 VGND.t2630 _275_.A2 _275_.ZN VGND.t2629 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1168 _451_.Q.t1 a_39264_18147# VGND.t6003 VGND.t6002 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1169 _474_.CLK.t4 a_48272_25156.t18 VPWR.t6549 VPWR.t6548 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1170 VPWR.t2693 a_46716_9432# a_46628_9476# VPWR.t2692 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1171 VPWR.t6403 _337_.A3.t4 a_24900_27912# VPWR.t6402 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X1172 a_44320_19369# a_43784_19369# VGND.t2560 VGND.t2559 nfet_06v0 ad=43.2f pd=0.6u as=0.2637p ps=1.825u w=0.36u l=0.6u
X1173 a_60212_25156# _251_.A1.t10 a_60064_25156# VPWR.t7010 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X1174 VPWR.t2732 a_66652_7431# a_66564_7528# VPWR.t2731 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1175 a_5388_16839# a_5300_16936# VGND.t2089 VGND.t2088 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1176 VPWR.t2775 a_5948_29816# a_5860_29860# VPWR.t2774 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1177 VPWR.t2191 a_36972_16839# a_36884_16936# VPWR.t2190 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1178 VGND.t2360 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I VGND.t2359 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1179 a_1468_20408# a_1380_20452# VGND.t2188 VGND.t2187 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1180 a_39178_23208# _301_.A1 _430_.ZN VPWR.t3350 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1181 a_27228_1592# a_27140_1636# VGND.t1780 VGND.t1779 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1182 VPWR.t1880 a_67660_13703# a_67572_13800# VPWR.t1879 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1183 VPWR.t652 a_33948_16839# a_33860_16936# VPWR.t651 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1184 a_30240_24776# a_29828_24455.t2 VGND.t6116 VGND.t6115 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1185 VGND.t1861 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I VGND.t1860 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1186 a_50068_27508# _408_.ZN VGND.t1863 VGND.t1862 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1187 VGND.t867 a_28054_30196# _355_.C.t2 VGND.t71 nfet_06v0 ad=0.2911p pd=1.53u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1188 VPWR.t5458 a_22524_1592# a_22436_1636# VPWR.t5457 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1189 a_47612_13703# a_47524_13800# VGND.t5275 VGND.t2950 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1190 VPWR.t2715 a_56460_13703# a_56372_13800# VPWR.t2714 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1191 a_46492_1592# a_46404_1636# VGND.t2579 VGND.t2578 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1192 VPWR.t2751 a_22636_28248# a_22548_28292# VPWR.t2750 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1193 a_61836_23544# a_61748_23588# VGND.t2620 VGND.t2619 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1194 a_42168_25640.t1 _284_.A2.t3 _284_.ZN.t1 VGND.t27 nfet_06v0 ad=0.3608p pd=2.52u as=0.30965p ps=1.685u w=0.82u l=0.6u
X1195 a_24100_29480# _343_.A2 VPWR.t1259 VPWR.t1258 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1196 _284_.B _397_.A1.t5 a_47636_25940# VGND.t8 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1197 _325_.B _325_.A1.t9 a_43668_19668# VGND.t6514 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1198 a_22304_26031# a_20084_26023.t3 a_22059_26399# VGND.t6682 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1199 VPWR.t6049 a_19328_28733# uio_out[6].t3 VPWR.t6048 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1200 VPWR.t2767 a_58924_18840# a_58836_18884# VPWR.t2766 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1201 VPWR.t2244 a_1916_5863# a_1828_5960# VPWR.t746 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1202 VPWR.t2246 a_22636_25112# a_22548_25156# VPWR.t2245 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1203 a_42168_22504# _305_.A2 _324_.B.t1 VGND.t2874 nfet_06v0 ad=0.3608p pd=2.52u as=0.30965p ps=1.685u w=0.82u l=0.6u
X1204 a_43784_19369# a_43400_18909# a_42996_18840# VGND.t3752 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1205 a_29916_2727# a_29828_2824# VGND.t2162 VGND.t2161 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1206 a_65980_12568# a_65892_12612# VGND.t4608 VGND.t4607 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1207 VPWR.t4761 a_1468_21976# a_1380_22020# VPWR.t4760 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1208 VPWR.t4763 a_53212_1159# a_53124_1256# VPWR.t4762 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1209 a_52512_19715# a_52064_19715.t3 a_52924_20127# VPWR.t6414 pfet_06v0 ad=0.1872p pd=1.4u as=43.2f ps=0.6u w=0.36u l=0.5u
X1210 VPWR.t4740 a_47724_18840# a_47636_18884# VPWR.t4739 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1211 VGND.t247 clkbuf_1_0__f_clk.I.t35 a_42392_22825.t12 VGND.t246 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1212 _358_.A2 _336_.Z a_30036_25940# VGND.t4413 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1213 VPWR.t965 a_1916_2727# a_1828_2824# VPWR.t964 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1214 a_61388_15704# a_61300_15748# VGND.t3025 VGND.t3024 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1215 a_39548_15704# a_39460_15748# VGND.t2575 VGND.t2574 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1216 VPWR.t1572 a_48956_2727# a_48868_2824# VPWR.t1571 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1217 VPWR.t2788 a_4604_20408# a_4516_20452# VPWR.t2787 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1218 VGND.t4311 _419_.Z a_47531_21258# VGND.t4310 nfet_06v0 ad=0.3124p pd=2.3u as=85.2f ps=0.95u w=0.71u l=0.6u
X1219 a_5948_1592# a_5860_1636# VGND.t2649 VGND.t2648 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1220 a_29692_21543# a_29604_21640# VGND.t2742 VGND.t2741 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1221 VPWR.t1014 a_1020_24679# a_932_24776# VPWR.t1013 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1222 a_44132_29535# a_42820_29159.t5 a_43788_29167# VPWR.t7040 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X1223 VPWR.t6467 _459_.CLK.t21 a_15828_27208.t0 VPWR.t6466 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1224 a_1468_14136# a_1380_14180# VGND.t2107 VGND.t2106 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1225 VPWR.t6528 _362_.B.t6 a_32628_26725# VPWR.t6527 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X1226 _290_.ZN _362_.B.t7 VGND.t6252 VGND.t6251 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1227 a_20672_30301# a_20379_29977# VGND.t1854 VGND.t71 nfet_06v0 ad=0.2119p pd=1.335u as=0.2333p ps=1.555u w=0.815u l=0.6u
X1228 VGND.t4894 a_42778_21812# a_43254_21236# VGND.t4893 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X1229 a_39172_22504# _311_.A2.t2 a_38968_22504# VGND.t6103 nfet_06v0 ad=88.2f pd=0.84u as=88.2f ps=0.84u w=0.42u l=0.6u
X1230 uio_out[6].t6 a_19328_28733# VGND.t5795 VGND.t5794 nfet_06v0 ad=0.2119p pd=1.335u as=0.2608p ps=1.455u w=0.815u l=0.6u
X1231 a_1468_11000# a_1380_11044# VGND.t1909 VGND.t1908 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1232 VPWR.t2222 a_25884_21543# a_25796_21640# VPWR.t2221 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1233 VGND.t1703 a_50084_24328# _381_.Z VGND.t1702 nfet_06v0 ad=0.224p pd=1.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1234 VGND.t6523 clk.t1 a_44296_24393.t1 VGND.t6522 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1235 a_17036_26247# a_16948_26344# VGND.t2125 VGND.t2124 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1236 VPWR.t2234 a_4156_12568# a_4068_12612# VPWR.t2233 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1237 a_30388_28776# _335_.ZN.t21 a_32904_28776# VGND.t6678 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1238 VGND.t328 a_42996_18840# a_42392_19243# VGND.t327 nfet_06v0 ad=0.142p pd=1.14u as=0.176p ps=1.68u w=0.4u l=0.6u
X1239 a_34715_22137# a_32740_22504.t3 a_34080_22461# VPWR.t100 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X1240 a_42236_1159# a_42148_1256# VGND.t2139 VGND.t2138 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1241 a_51892_23340# _424_.B1.t8 a_51668_23340# VPWR.t6616 pfet_06v0 ad=0.1736p pd=1.18u as=0.1736p ps=1.18u w=0.56u l=0.5u
X1242 a_17036_23111# a_16948_23208# VGND.t2696 VGND.t2363 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1243 a_26108_2727# a_26020_2824# VGND.t2552 VGND.t2551 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1244 VPWR.t2691 a_29468_1159# a_29380_1256# VPWR.t2690 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1245 a_51196_15271# a_51108_15368# VGND.t2556 VGND.t2555 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1246 a_58476_10567# a_58388_10664# VGND.t4483 VGND.t4482 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1247 VPWR.t4639 a_50748_1592# a_50660_1636# VPWR.t4638 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1248 a_2812_9432# a_2724_9476# VGND.t2587 VGND.t2586 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1249 VPWR.t1016 a_45148_2727# a_45060_2824# VPWR.t1015 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1250 a_3260_26247# a_3172_26344# VGND.t2589 VGND.t2588 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1251 a_39256_28292# _437_.A1.t5 _285_.Z VPWR.t6859 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1252 a_2812_6296# a_2724_6340# VGND.t2087 VGND.t2086 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1253 _258_.I _238_.ZN a_59572_29076# VGND.t5916 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1254 VGND.t394 a_18096_27165# uio_out[7].t7 VGND.t393 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1255 a_1916_12568# a_1828_12612# VGND.t2563 VGND.t1214 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1256 a_3260_23111# a_3172_23208# VGND.t2564 VGND.t2192 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1257 a_52068_29480# _268_.A1.t3 _275_.A2 VPWR.t6735 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1258 VPWR.t2743 a_4604_14136# a_4516_14180# VPWR.t2742 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1259 a_32096_24419# a_31803_24831# VPWR.t3163 VPWR.t3162 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X1260 a_20496_26344# a_20084_26023.t4 VGND.t6684 VGND.t6683 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1261 VGND.t2248 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN VGND.t2247 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1262 _474_.D _218_.ZN a_49988_21236# VGND.t3632 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1263 VPWR.t2786 a_4604_11000# a_4516_11044# VPWR.t2785 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1264 a_32848_29123# a_32476_29167# VPWR.t4997 VPWR.t4996 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X1265 VPWR.t4517 a_28460_20408# a_28372_20452# VPWR.t4516 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1266 VPWR.t3341 a_1020_15271# a_932_15368# VPWR.t3340 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1267 VPWR.t1795 a_50084_24328# _381_.Z VPWR.t1794 pfet_06v0 ad=0.389p pd=2.02u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1268 a_4828_2727# a_4740_2824# VGND.t3196 VGND.t3195 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1269 VPWR.t2213 a_58588_12568# a_58500_12612# VPWR.t2212 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1270 VPWR.t5667 a_62172_19975# a_62084_20072# VPWR.t5666 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1271 VPWR.t2215 a_27900_21543# a_27812_21640# VPWR.t2214 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1272 a_21740_29383# a_21652_29480# VGND.t2064 VGND.t2063 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1273 a_14796_26680# a_14708_26724# VGND.t2066 VGND.t2065 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1274 a_52316_9432# a_52228_9476# VGND.t1844 VGND.t1843 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1275 a_35816_21192# _317_.A2 VPWR.t2579 VPWR.t2578 pfet_06v0 ad=0.156p pd=1.12u as=0.40575p ps=2.055u w=0.6u l=0.5u
X1276 a_64412_15271# a_64324_15368# VGND.t1846 VGND.t1845 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1277 _244_.Z a_60212_25156# VGND.t2593 VGND.t2592 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1278 VPWR.t1876 a_61836_26680# a_61748_26724# VPWR.t1875 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1279 VPWR.t2307 a_25652_31048# a_25652_31048# VPWR.t2306 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1280 a_16140_20408# a_16052_20452# VGND.t2201 VGND.t2200 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1281 a_44736_26031# a_43736_25896# VGND.t3959 VGND.t3958 nfet_06v0 ad=43.2f pd=0.6u as=0.142p ps=1.14u w=0.36u l=0.6u
X1282 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN VPWR.t6279 VPWR.t6278 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1283 _431_.A3 _437_.A1.t6 VGND.t6546 VGND.t6545 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1284 VPWR.t2169 a_4940_4295# a_4852_4392# VPWR.t2168 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1285 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN VPWR.t2605 VPWR.t1708 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1286 VPWR.t2071 a_54780_18840# a_54692_18884# VPWR.t2070 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1287 a_43232_29480# a_42820_29159.t6 VPWR.t7042 VPWR.t7041 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1288 a_9084_30951# a_8996_31048# VGND.t2624 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1289 a_35740_30951# a_35652_31048# VGND.t2625 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1290 VPWR.t2763 a_54780_15704# a_54692_15748# VPWR.t2762 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1291 a_67548_17272# a_67460_17316# VGND.t2637 VGND.t2636 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1292 VPWR.t2779 a_62508_23111# a_62420_23208# VPWR.t2778 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1293 a_18088_26841# a_16240_26795# a_17803_26841# VPWR.t5617 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X1294 a_32604_19975# a_32516_20072# VGND.t2583 VGND.t2582 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1295 VPWR.t2722 a_43580_15704# a_43492_15748# VPWR.t699 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1296 a_3260_16839# a_3172_16936# VGND.t2081 VGND.t2080 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1297 VPWR.t2184 vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I VPWR.t2183 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1298 VPWR.t2024 a_37472_24419# a_37464_24831# VPWR.t2023 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X1299 a_26220_21976# a_26132_22020# VGND.t1924 VGND.t1923 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1300 a_35292_26247# a_35204_26344# VGND.t3212 VGND.t3211 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1301 VPWR.t3359 a_16140_21976# a_16052_22020# VPWR.t2982 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1302 a_19328_28733# a_19035_28409# VGND.t3522 VGND.t3521 nfet_06v0 ad=0.2119p pd=1.335u as=0.2333p ps=1.555u w=0.815u l=0.6u
X1303 VPWR.t2258 a_51956_26183# a_51576_25896# VPWR.t2257 pfet_06v0 ad=0.23p pd=1.54u as=0.352p ps=2.48u w=0.8u l=0.5u
X1304 VPWR.t2264 a_55452_15271# a_55364_15368# VPWR.t2263 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1305 VPWR.t2747 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I VPWR.t2746 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1306 uo_out[4].t0 _287_.A1.t13 a_34708_29860# VPWR.t6778 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1307 a_46716_14136# a_46628_14180# VGND.t2613 VGND.t2612 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1308 VPWR.t1839 a_5052_28248# a_4964_28292# VPWR.t1838 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1309 a_27760_25273# a_27328_25227# VPWR.t6293 VPWR.t6292 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X1310 a_60380_11000# a_60292_11044# VGND.t1338 VGND.t1337 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1311 a_46716_11000# a_46628_11044# VGND.t1340 VGND.t1339 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1312 a_24092_23111# a_24004_23208# VGND.t1342 VGND.t1341 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1313 VPWR.t1854 a_49404_12568# a_49316_12612# VPWR.t1853 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1314 VPWR.t1856 a_64860_17272# a_64772_17316# VPWR.t1855 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1315 VPWR.t4386 a_5052_25112# a_4964_25156# VPWR.t4385 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1316 a_25884_27815# a_25796_27912# VGND.t4230 VGND.t4229 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1317 VPWR.t1969 a_33052_15271# a_32964_15368# VPWR.t1968 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1318 a_39256_28292# a_38584_28292# VPWR.t4050 VPWR.t4049 pfet_06v0 ad=0.3172p pd=1.74u as=0.4005p ps=2.12u w=1.22u l=0.5u
X1319 VGND.t4704 _250_.A2 a_62763_28776# VGND.t4703 nfet_06v0 ad=0.3124p pd=2.3u as=85.2f ps=0.95u w=0.71u l=0.6u
X1320 _416_.A3 _324_.B.t21 VGND.t6414 VGND.t6413 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1321 VPWR.t2719 a_53660_17272# a_53572_17316# VPWR.t2718 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1322 _474_.CLK.t5 a_48272_25156.t19 VPWR.t6551 VPWR.t6550 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1323 a_41996_28777# _265_.ZN a_41828_28777# VGND.t298 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X1324 VPWR.t2895 a_48888_19243# _474_.Q VPWR.t2894 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1325 VGND.t4815 a_38472_30169# _287_.A1.t6 VGND.t1059 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X1326 _352_.A2.t15 _350_.A1.t4 a_29736_27508# VGND.t6338 nfet_06v0 ad=0.2132p pd=1.34u as=98.39999f ps=1.06u w=0.82u l=0.6u
X1327 VPWR.t2897 a_1916_18840# a_1828_18884# VPWR.t2896 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1328 VPWR.t4329 _476_.Q _422_.ZN VPWR.t4328 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1329 VPWR.t3023 _305_.A2 a_44500_22020# VPWR.t3022 pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X1330 a_47376_27912# _304_.B a_47172_27912# VPWR.t4698 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1331 a_35892_19369# a_35092_19368.t2 VGND.t83 VGND.t82 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1332 _452_.D _330_.A1.t8 a_41776_18504# VPWR.t210 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1333 VPWR.t2040 a_1916_15704# a_1828_15748# VPWR.t2039 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1334 VPWR.t6581 _447_.Q.t5 _300_.ZN VPWR.t6580 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1335 VPWR.t2041 a_31260_17272# a_31172_17316# VPWR.t766 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1336 a_24540_24679# a_24452_24776# VGND.t2661 VGND.t2660 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1337 a_28552_25940# _337_.A3.t5 VGND.t6136 VGND.t6135 nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1338 a_46044_1159# a_45956_1256# VGND.t2129 VGND.t2128 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1339 _238_.ZN _238_.I VPWR.t2239 VPWR.t2238 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1340 a_24540_21543# a_24452_21640# VGND.t2135 VGND.t2134 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1341 a_50748_20408# a_50660_20452# VGND.t2150 VGND.t2149 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1342 a_43468_16839# a_43380_16936# VGND.t2152 VGND.t2151 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1343 VPWR.t1123 a_48396_16839# a_48308_16936# VPWR.t1122 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1344 VPWR.t1832 a_40668_20408# a_40580_20452# VPWR.t1831 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1345 a_28908_20408# a_28820_20452# VGND.t1744 VGND.t1743 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1346 VPWR.t6302 a_31932_21543# a_31844_21640# VPWR.t6301 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1347 VPWR.t5124 a_15244_24679# a_15156_24776# VPWR.t666 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1348 _328_.A2 _325_.A2.t3 a_44276_20072# VPWR.t6390 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1349 a_31372_20408# a_31284_20452# VGND.t2224 VGND.t2223 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1350 VPWR.t6047 a_19328_28733# uio_out[6].t2 VPWR.t6046 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1351 VPWR.t1809 a_21292_20408# a_21204_20452# VPWR.t1808 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1352 VPWR.t1810 a_33724_1159# a_33636_1256# VPWR.t673 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1353 a_41432_17801# a_41088_17757.t2 a_40644_17272# VPWR.t161 pfet_06v0 ad=0.1791p pd=1.355u as=0.1665p ps=1.285u w=0.36u l=0.5u
X1354 _337_.A3.t1 a_26160_27165# VGND.t928 VGND.t927 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1355 VPWR.t1850 a_54108_21543# a_54020_21640# VPWR.t1849 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1356 VGND.t249 clkbuf_1_0__f_clk.I.t36 a_42392_22825.t11 VGND.t248 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1357 VPWR.t6553 a_48272_25156.t20 _474_.CLK.t6 VPWR.t6552 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1358 VGND.t6264 a_48272_25156.t21 _474_.CLK.t7 VGND.t6263 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1359 a_51308_19369# _474_.D a_50384_19204# VGND.t2537 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X1360 VPWR.t3238 a_37084_25112# a_36996_25156# VPWR.t3237 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1361 VPWR.t1896 a_66652_9432# a_66564_9476# VPWR.t578 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1362 a_1468_10567# a_1380_10664# VGND.t1800 VGND.t1799 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1363 a_39996_15704# a_39908_15748# VGND.t1952 VGND.t1951 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1364 a_53436_1592# a_53348_1636# VGND.t1954 VGND.t1953 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1365 a_53324_10567# a_53236_10664# VGND.t3384 VGND.t3383 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1366 VPWR.t3539 a_67100_5863# a_67012_5960# VPWR.t995 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1367 a_53548_18407# a_53460_18504# VGND.t3388 VGND.t3387 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1368 a_50796_19001# a_50280_19369# VPWR.t1464 VPWR.t1463 pfet_06v0 ad=43.2f pd=0.6u as=0.1044p ps=0.94u w=0.36u l=0.5u
X1369 a_38616_24328# _438_.A2 a_39004_24463# VGND.t4964 nfet_06v0 ad=0.1606p pd=1.61u as=58.39999f ps=0.685u w=0.365u l=0.6u
X1370 VPWR.t2939 a_28908_21976# a_28820_22020# VPWR.t2938 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1371 a_39860_25156# _416_.A1.t5 _442_.ZN VPWR.t201 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1372 VPWR.t2942 a_33948_18840# a_33860_18884# VPWR.t2941 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1373 VPWR.t2080 a_31372_21976# a_31284_22020# VPWR.t2079 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1374 VPWR.t690 a_67100_2727# a_67012_2824# VPWR.t689 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1375 VGND.t5334 vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN VGND.t605 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1376 a_14908_30951# a_14820_31048# VGND.t1751 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1377 VPWR.t1843 a_42460_1592# a_42372_1636# VPWR.t1842 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1378 a_61948_14136# a_61860_14180# VGND.t1913 VGND.t1912 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1379 VPWR.t2012 a_33948_15704# a_33860_15748# VPWR.t2011 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1380 VPWR.t2014 a_20172_21976# a_20084_22020# VPWR.t2013 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1381 VPWR.t1494 vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I VPWR.t1493 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1382 _437_.ZN _447_.Q.t6 VGND.t6303 VGND.t6302 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1383 a_17484_26247# a_17396_26344# VGND.t2071 VGND.t1408 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1384 VPWR.t686 a_36076_18407# a_35988_18504# VPWR.t685 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1385 VPWR.t5006 _475_.Q _384_.A3.t9 VPWR.t5005 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1386 a_61948_11000# a_61860_11044# VGND.t2091 VGND.t2090 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1387 a_50748_14136# a_50660_14180# VGND.t3030 VGND.t2879 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1388 a_4156_8999# a_4068_9096# VGND.t3032 VGND.t3031 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1389 VPWR.t3191 a_64636_12568# a_64548_12612# VPWR.t3190 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1390 a_17484_23111# a_17396_23208# VGND.t2826 VGND.t1613 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1391 a_28228_25273# a_26916_25640.t5 a_27884_25641# VPWR.t6776 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X1392 a_20844_26680# a_20756_26724# VGND.t3476 VGND.t3475 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1393 a_46156_26031# _402_.ZN a_45232_25987# VGND.t3477 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X1394 VGND.t2816 _352_.ZN _457_.D VGND.t2815 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1395 VPWR.t5958 a_39212_16839# a_39124_16936# VPWR.t5957 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1396 VPWR.t1295 a_52920_22760# _384_.A1 VPWR.t1294 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1397 a_2812_2727# a_2724_2824# VGND.t1221 VGND.t1220 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1398 a_50748_11000# a_50660_11044# VGND.t1223 VGND.t1222 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1399 VPWR.t6872 _229_.I.t4 a_63105_28293# VPWR.t6871 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1400 a_4156_5863# a_4068_5960# VGND.t3299 VGND.t1375 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1401 a_2812_25112# a_2724_25156# VGND.t1290 VGND.t1289 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1402 VPWR.t1361 a_22560_30288# uio_out[4].t0 VPWR.t1360 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1403 VPWR.t1363 a_1916_4728# a_1828_4772# VPWR.t1362 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1404 a_49852_2727# a_49764_2824# VGND.t5766 VGND.t3321 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1405 VGND.t2599 _379_.A2 a_18760_29032# VGND.t2598 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1406 VPWR.t3545 a_57132_12135# a_57044_12232# VPWR.t3544 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1407 a_37464_24831# a_35616_24776# a_37179_24831# VPWR.t1667 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X1408 VGND.t1853 a_20379_29977# a_20672_30301# VGND.t71 nfet_06v0 ad=0.2608p pd=1.455u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1409 a_2812_21976# a_2724_22020# VGND.t3393 VGND.t2943 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1410 VPWR.t1301 a_1916_1592# a_1828_1636# VPWR.t1300 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1411 VPWR.t1303 a_24988_1592# a_24900_1636# VPWR.t1302 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1412 a_46356_24072# _324_.C.t12 VGND.t6503 VGND.t6502 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1413 VPWR.t2393 a_36148_21976# _317_.A2 VPWR.t2392 pfet_06v0 ad=0.4268p pd=2.175u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1414 VPWR.t2397 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t2396 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1415 _350_.A2.t10 _371_.A1.t11 a_30596_28292# VPWR.t6509 pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
X1416 a_3708_18407# a_3620_18504# VGND.t5780 VGND.t5498 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1417 a_46984_23588# _281_.ZN.t6 VGND.t122 VGND.t121 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1418 VPWR.t6030 a_41188_18840# _327_.Z VPWR.t6029 pfet_06v0 ad=0.4268p pd=2.175u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1419 VPWR.t6119 a_19388_2727# a_19300_2824# VPWR.t6118 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1420 VPWR.t3084 a_61948_1159# a_61860_1256# VPWR.t3083 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1421 VPWR.t3086 a_48956_1592# a_48868_1636# VPWR.t3085 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1422 VPWR.t1900 a_1020_23544# a_932_23588# VPWR.t1899 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1423 a_2364_17272# a_2276_17316# VGND.t1803 VGND.t489 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1424 a_37964_18191# _330_.ZN a_37796_18191# VGND.t6042 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X1425 VPWR.t6312 a_58028_17272# a_57940_17316# VPWR.t6311 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1426 a_39004_24463# _437_.A1.t7 VGND.t6548 VGND.t6547 nfet_06v0 ad=58.39999f pd=0.685u as=0.23405p ps=1.555u w=0.365u l=0.6u
X1427 a_17932_24679# a_17844_24776# VGND.t5740 VGND.t2367 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1428 _373_.A2 _350_.A1.t5 a_28672_31048# VPWR.t6622 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1429 a_52316_2727# a_52228_2824# VGND.t2562 VGND.t2561 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1430 VGND.t159 a_41088_17757.t3 a_42460_17801# VGND.t158 nfet_06v0 ad=0.1584p pd=1.6u as=43.2f ps=0.6u w=0.36u l=0.6u
X1431 VPWR.t2139 a_55676_1159# a_55588_1256# VPWR.t2138 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1432 a_51912_20452# a_51240_20452# VPWR.t469 VPWR.t468 pfet_06v0 ad=0.3172p pd=1.74u as=0.4005p ps=2.12u w=1.22u l=0.5u
X1433 a_17932_21543# a_17844_21640# VGND.t370 VGND.t369 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1434 a_18096_27165# a_17803_26841# VPWR.t1340 VPWR.t1339 pfet_06v0 ad=0.2457p pd=1.465u as=0.2619p ps=1.685u w=0.945u l=0.5u
X1435 VPWR.t384 a_2364_4295# a_2276_4392# VPWR.t383 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1436 a_48272_25156.t13 clkbuf_1_0__f_clk.I.t37 VGND.t251 VGND.t250 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1437 VPWR.t637 a_2364_1159# a_2276_1256# VPWR.t356 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1438 VGND.t4562 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN _251_.ZN VGND.t4561 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1439 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN VPWR.t6277 VPWR.t6276 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1440 VPWR.t386 a_50300_15271# a_50212_15368# VPWR.t385 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1441 _452_.CLK.t1 a_42392_22825.t15 VPWR.t6910 VPWR.t6909 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1442 a_53660_15271# a_53572_15368# VGND.t376 VGND.t375 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1443 VGND.t211 _330_.A1.t9 _448_.D VGND.t210 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X1444 a_46044_2727# a_45956_2824# VGND.t639 VGND.t638 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1445 VPWR.t1764 _441_.A3 a_40316_23233# VPWR.t1763 pfet_06v0 ad=0.5913p pd=3.27u as=0.2847p ps=1.615u w=1.095u l=0.5u
X1446 a_30140_23111# a_30052_23208# VGND.t4175 VGND.t4174 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1447 VPWR.t4343 a_6172_30951# a_6084_31048# VPWR.t4342 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1448 VGND.t4419 a_51240_19624# _476_.Q VGND.t4418 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1449 VPWR.t4568 a_54780_26247# a_54692_26344# VPWR.t4567 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1450 a_43936_27165# a_43564_27209# VGND.t4423 VGND.t4422 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X1451 a_46352_22021# _402_.B VPWR.t3274 VPWR.t3273 pfet_06v0 ad=0.44955p pd=1.955u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1452 VGND.t4721 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN VGND.t4720 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1453 _441_.A3 _260_.A2 VPWR.t6289 VPWR.t6288 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1454 VGND.t6039 a_43296_28733# a_43248_28777# VGND.t6038 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X1455 a_48376_27508# _402_.A1.t9 VGND.t6432 VGND.t6431 nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1456 a_49740_10567# a_49652_10664# VGND.t6041 VGND.t6040 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1457 VPWR.t773 a_65084_2727# a_64996_2824# VPWR.t772 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1458 VPWR.t4932 a_45148_1592# a_45060_1636# VPWR.t4931 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1459 a_67996_17272# a_67908_17316# VGND.t4785 VGND.t4784 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1460 a_2812_15704# a_2724_15748# VGND.t1498 VGND.t1497 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1461 a_31260_15271# a_31172_15368# VGND.t1500 VGND.t1499 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1462 VPWR.t3798 a_62956_23111# a_62868_23208# VPWR.t3797 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1463 a_40452_23588# _441_.A3 VPWR.t1762 VPWR.t1761 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1464 a_37312_19369# a_35092_19368.t3 a_37067_19001# VGND.t84 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1465 _358_.A2 _352_.A2.t19 a_29828_26344# VPWR.t6985 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1466 VPWR.t6052 a_1468_27815# a_1380_27912# VPWR.t3823 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1467 a_50636_12135# a_50548_12232# VGND.t5801 VGND.t5800 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1468 VPWR.t4126 a_51048_26680# _284_.A2.t0 VPWR.t4125 pfet_06v0 ad=0.40575p pd=2.055u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1469 VPWR.t4128 a_19276_25112# a_19188_25156# VPWR.t4127 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1470 a_46716_10567# a_46628_10664# VGND.t3976 VGND.t2557 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1471 VPWR.t6259 a_32380_26247# a_32292_26344# VPWR.t6258 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1472 VPWR.t6261 a_18716_26247# a_18628_26344# VPWR.t6260 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1473 a_43788_29167# _480_.Q a_43664_29535# VPWR.t5084 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X1474 VPWR.t1951 a_32380_23111# a_32292_23208# VPWR.t1950 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1475 a_47164_30951# a_47076_31048# VGND.t1857 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1476 a_40038_28720# _234_.ZN VPWR.t3599 VPWR.t3598 pfet_06v0 ad=0.5368p pd=3.32u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1477 a_5724_29383# a_5636_29480# VGND.t5097 VGND.t5096 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1478 VPWR.t5265 a_18716_23111# a_18628_23208# VPWR.t5264 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1479 _441_.A3 _452_.Q.t8 a_39985_24372# VGND.t6639 nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X1480 VPWR.t3674 a_51084_10567# a_50996_10664# VPWR.t3673 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1481 a_30796_24463# _459_.D a_30628_24463# VGND.t2971 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X1482 a_34260_29860# _287_.A1.t14 uo_out[4].t1 VPWR.t6779 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1483 a_34396_17272# a_34308_17316# VGND.t3244 VGND.t3243 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1484 VGND.t3253 _327_.A2 a_42811_19668# VGND.t3252 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1485 a_3260_7864# a_3172_7908# VGND.t3254 VGND.t2269 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1486 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN VGND.t2103 VGND.t2102 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1487 VPWR.t4152 a_49852_12568# a_49764_12612# VPWR.t4151 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1488 a_42908_1159# a_42820_1256# VGND.t4000 VGND.t3999 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1489 a_33483_29535# a_31508_29159.t3 a_32848_29123# VPWR.t94 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X1490 a_3260_4728# a_3172_4772# VGND.t5676 VGND.t2713 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1491 VPWR.t5247 a_54444_16839# a_54356_16936# VPWR.t5246 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1492 a_39536_26795# a_39124_27208.t2 VGND.t226 VGND.t225 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1493 VPWR.t1998 a_4940_26247# a_4852_26344# VPWR.t1997 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1494 VPWR.t2000 a_1916_29383# a_1828_29480# VPWR.t1999 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1495 VPWR.t6882 _448_.Q.t3 a_37384_19624# VPWR.t6881 pfet_06v0 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X1496 VPWR.t1514 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN VPWR.t1513 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1497 a_42320_28777# a_41440_28363# a_41996_28777# VGND.t1455 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X1498 VPWR.t6370 a_52400_25987.t2 a_52360_26355# VPWR.t6369 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1499 VPWR.t3287 a_4940_23111# a_4852_23208# VPWR.t3286 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1500 VPWR.t5340 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I VPWR.t5339 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1501 VGND.t884 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN VGND.t883 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1502 VPWR.t3156 a_1916_26247# a_1828_26344# VPWR.t962 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1503 a_46828_30345# _393_.ZN a_45904_30180# VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X1504 a_4156_1159# a_4068_1256# VGND.t4085 VGND.t4084 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1505 a_22992_27555# a_22620_27599# VGND.t4087 VGND.t4086 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X1506 VPWR.t4254 a_61164_12135# a_61076_12232# VPWR.t4253 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1507 a_66652_4295# a_66564_4392# VGND.t3717 VGND.t1793 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1508 a_62620_18407# a_62532_18504# VGND.t3719 VGND.t3718 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1509 VPWR.t3861 a_1916_23111# a_1828_23208# VPWR.t2669 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1510 VPWR.t499 a_64300_10567# a_64212_10664# VPWR.t498 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1511 a_1468_9432# a_1380_9476# VGND.t4187 VGND.t1799 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1512 VPWR.t4467 _416_.A3 a_47252_18884# VPWR.t4466 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1513 a_34844_15704# a_34756_15748# VGND.t1872 VGND.t1871 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1514 VGND.t129 _417_.A2.t4 _416_.A3 VGND.t128 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1515 VPWR.t1394 a_1468_18407# a_1380_18504# VPWR.t1393 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1516 a_5388_8999# a_5300_9096# VGND.t1874 VGND.t1873 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1517 VGND.t3059 a_29856_29123# a_29808_29167# VGND.t3058 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X1518 _378_.I _346_.B VPWR.t414 VPWR.t413 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1519 a_1468_6296# a_1380_6340# VGND.t3063 VGND.t3062 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1520 a_3260_26680# a_3172_26724# VGND.t4402 VGND.t2751 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1521 VPWR.t2036 a_39268_18840# _330_.A2 VPWR.t2035 pfet_06v0 ad=0.34437p pd=1.895u as=0.31207p ps=1.665u w=1.095u l=0.5u
X1522 a_21180_1592# a_21092_1636# VGND.t4060 VGND.t4059 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1523 a_5388_5863# a_5300_5960# VGND.t4062 VGND.t4061 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1524 VPWR.t2992 a_15692_24679# a_15604_24776# VPWR.t2991 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1525 a_24864_29931# a_24452_30344.t3 VPWR.t159 VPWR.t158 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1526 _441_.A3 _430_.ZN VPWR.t4822 VPWR.t4821 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X1527 _443_.D _437_.A1.t8 VGND.t6550 VGND.t6549 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1528 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I VPWR.t751 VPWR.t750 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1529 a_61052_12568# a_60964_12612# VGND.t3881 VGND.t3880 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1530 VPWR.t4656 a_36656_29123# a_36628_29535# VPWR.t4655 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X1531 VPWR.t2958 a_43936_27165# a_43908_26841# VPWR.t2957 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X1532 VPWR.t1943 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN VPWR.t1942 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1533 VPWR.t1945 a_54556_21543# a_54468_21640# VPWR.t1944 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1534 VGND.t6266 a_48272_25156.t22 _474_.CLK.t8 VGND.t6265 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1535 _408_.ZN _411_.A2.t8 VPWR.t115 VPWR.t114 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1536 VGND.t6505 _324_.C.t13 _416_.A1.t2 VGND.t6504 nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
X1537 a_64972_10567# a_64884_10664# VGND.t2899 VGND.t2898 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1538 uo_out[3].t7 a_41160_29083# VGND.t4033 VGND.t4032 nfet_06v0 ad=0.1183p pd=0.975u as=0.2002p ps=1.79u w=0.455u l=0.6u
X1539 a_64412_18840# a_64324_18884# VGND.t2900 VGND.t2739 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1540 VPWR.t3463 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN VPWR.t3462 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1541 a_20508_23111# a_20420_23208# VGND.t1865 VGND.t1864 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1542 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I VPWR.t2501 VPWR.t2500 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1543 a_1468_29816# a_1380_29860# VGND.t1866 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1544 a_53772_10567# a_53684_10664# VGND.t1916 VGND.t1915 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1545 a_53996_18407# a_53908_18504# VGND.t1918 VGND.t1917 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1546 VPWR.t5691 a_47612_2727# a_47524_2824# VPWR.t5690 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1547 VPWR.t2075 a_67100_17272# a_67012_17316# VPWR.t2074 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1548 a_45920_20523# a_45508_20936.t4 VPWR.t200 VPWR.t199 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1549 a_27676_1592# a_27588_1636# VGND.t1978 VGND.t1977 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1550 a_4604_1592# a_4516_1636# VGND.t5762 VGND.t5761 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1551 a_61276_1159# a_61188_1256# VGND.t5764 VGND.t5763 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1552 VGND.t6001 a_39264_18147# a_39216_18191# VGND.t6000 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X1553 VPWR.t3959 a_22972_1592# a_22884_1636# VPWR.t3958 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1554 a_52852_24372# _427_.B1 _478_.D VGND.t3814 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1555 VPWR.t3871 a_34448_25597# _460_.Q VPWR.t3870 pfet_06v0 ad=0.854p pd=3.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1556 a_58028_12135# a_57940_12232# VGND.t3439 VGND.t3438 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1557 VPWR.t3591 a_37644_23544# a_37556_23588# VPWR.t3590 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1558 VPWR.t3593 a_46940_1592# a_46852_1636# VPWR.t3592 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1559 VPWR.t4779 a_10428_1159# a_10340_1256# VPWR.t4778 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1560 VGND.t4366 a_32848_29123# a_32800_29167# VGND.t4365 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X1561 _474_.CLK.t9 a_48272_25156.t23 VPWR.t6555 VPWR.t6554 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1562 a_34440_25273# a_32592_25227# a_34155_25273# VPWR.t5913 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X1563 VGND.t269 a_44296_24393.t20 clkbuf_1_0__f_clk.I.t30 VGND.t268 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1564 VPWR.t5916 a_16140_27815# a_16052_27912# VPWR.t2872 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1565 VPWR.t4059 a_22748_23111# a_22660_23208# VPWR.t4058 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1566 VPWR.t4652 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN VPWR.t4651 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1567 a_34732_16839# a_34644_16936# VGND.t3914 VGND.t3913 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1568 VPWR.t986 a_39660_16839# a_39572_16936# VPWR.t985 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1569 a_67212_20408# a_67124_20452# VGND.t3653 VGND.t3652 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1570 VPWR.t3804 a_15244_23544# a_15156_23588# VPWR.t3803 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1571 VPWR.t6204 a_53660_1159# a_53572_1256# VPWR.t6203 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1572 VGND.t5704 _293_.A2 uo_out[1].t11 VGND.t3446 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1573 VPWR.t4150 a_3260_7864# a_3172_7908# VPWR.t373 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1574 a_4156_20408# a_4068_20452# VGND.t3055 VGND.t3054 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1575 VPWR.t4145 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I VPWR.t4144 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1576 a_25296_29977# a_24864_29931# VPWR.t4038 VPWR.t4037 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X1577 VPWR.t3214 a_57580_12135# a_57492_12232# VPWR.t3213 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1578 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN VPWR.t2272 VPWR.t2271 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1579 a_20060_2727# a_19972_2824# VGND.t3553 VGND.t3552 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1580 VPWR.t3137 a_28124_1159# a_28036_1256# VPWR.t3136 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1581 a_31708_16839# a_31620_16936# VGND.t1842 VGND.t1430 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1582 a_43664_17317# _325_.B VPWR.t2765 VPWR.t2764 pfet_06v0 ad=0.44955p pd=1.955u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1583 a_46356_24072# _399_.ZN _402_.B VGND.t1187 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1584 a_48141_29480# _388_.B a_47525_29480# VPWR.t4316 pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X1585 VPWR.t2721 a_32604_19975# a_32516_20072# VPWR.t2720 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1586 VPWR.t1596 a_41536_17636# a_41432_17801# VPWR.t1595 pfet_06v0 ad=0.1044p pd=0.94u as=0.1791p ps=1.355u w=0.36u l=0.5u
X1587 a_1468_23544# a_1380_23588# VGND.t3344 VGND.t3343 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1588 VPWR.t4243 a_1020_30951# a_932_31048# VPWR.t4242 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1589 a_28596_27916.t3 _350_.A2.t21 _352_.A2.t3 VPWR.t6574 pfet_06v0 ad=0.528p pd=3.28u as=0.312p ps=1.72u w=1.2u l=0.5u
X1590 a_3708_7431# a_3620_7528# VGND.t4081 VGND.t4080 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1591 VPWR.t4055 a_67100_4728# a_67012_4772# VPWR.t4054 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1592 VPWR.t4057 a_58476_17272# a_58388_17316# VPWR.t4056 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1593 a_32828_2727# a_32740_2824# VGND.t3902 VGND.t1624 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1594 a_47291_25940# _402_.A1.t10 _400_.ZN VGND.t6433 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1595 VPWR.t2008 a_4156_21976# a_4068_22020# VPWR.t2007 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1596 a_46352_20569# a_45920_20523# VPWR.t2078 VPWR.t2077 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X1597 VPWR.t1039 a_51868_2727# a_51780_2824# VPWR.t1038 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1598 a_46716_1159# a_46628_1256# VGND.t1968 VGND.t1967 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1599 VPWR.t978 a_46716_18407# a_46628_18504# VPWR.t977 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1600 VGND.t2645 a_32096_24419# a_32048_24463# VGND.t2644 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X1601 uo_out[3].t1 a_41160_29083# VPWR.t4184 VPWR.t4183 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1602 a_32820_29535# a_31508_29159.t4 a_32476_29167# VPWR.t95 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X1603 a_26556_2727# a_26468_2824# VGND.t5963 VGND.t5962 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1604 VPWR.t6987 _352_.A2.t20 a_30724_26020# VPWR.t6986 pfet_06v0 ad=0.4268p pd=2.175u as=0.1391p ps=1.055u w=0.535u l=0.5u
X1605 _452_.CLK.t2 a_42392_22825.t16 VPWR.t6912 VPWR.t6911 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1606 VPWR.t3597 a_55900_12568# a_55812_12612# VPWR.t3596 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1607 VPWR.t1117 a_45596_2727# a_45508_2824# VPWR.t1116 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1608 a_4156_14136# a_4068_14180# VGND.t3445 VGND.t3444 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1609 a_51196_21543# a_51108_21640# VGND.t2902 VGND.t2901 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1610 a_44816_27209# a_42596_27208.t3 a_44571_26841# VGND.t143 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1611 _452_.CLK.t3 a_42392_22825.t17 VGND.t6599 VGND.t6598 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X1612 _416_.A2 _419_.A4 a_47860_21640# VPWR.t4134 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1613 a_65756_27815# a_65668_27912# VGND.t5777 VGND.t5776 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1614 VGND.t889 _395_.A1 _390_.ZN VGND.t888 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1615 a_60064_25156# vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN VPWR.t4160 VPWR.t4159 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1616 a_4156_11000# a_4068_11044# VGND.t4009 VGND.t4008 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1617 VPWR.t4163 a_54108_14136# a_54020_14180# VPWR.t4162 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1618 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN VGND.t1453 VGND.t1452 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1619 a_65084_15271# a_64996_15368# VGND.t5716 VGND.t5478 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1620 VPWR.t5944 a_54108_11000# a_54020_11044# VPWR.t5943 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1621 VPWR.t2043 a_19388_1592# a_19300_1636# VPWR.t2042 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1622 _334_.A1 a_37584_29123# VPWR.t2049 VPWR.t2048 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1623 VPWR.t2051 a_61948_27815# a_61860_27912# VPWR.t2050 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1624 a_37840_18559# a_37408_18504# VPWR.t1848 VPWR.t1847 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X1625 VPWR.t5981 a_44252_30951# a_44164_31048# VPWR.t5980 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1626 a_35504_18955# a_35092_19368.t4 VGND.t86 VGND.t85 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1627 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN VPWR.t5608 VPWR.t5607 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1628 VGND.t5426 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I VGND.t5425 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1629 a_31120_24463# a_30240_24776# a_30796_24463# VGND.t6050 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X1630 _223_.ZN _223_.I VPWR.t7113 VPWR.t7112 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1631 a_49068_20408# _474_.Q VPWR.t4801 VPWR.t4800 pfet_06v0 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1632 VPWR.t6796 _324_.C.t14 _424_.B1.t3 VPWR.t6795 pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1633 a_4604_12568# a_4516_12612# VGND.t6783 VGND.t6782 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1634 VPWR.t5312 a_54892_16839# a_54804_16936# VPWR.t5311 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1635 a_43888_19204# a_43400_18909# a_44320_19369# VGND.t3751 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X1636 a_43750_23544# a_44162_24120# a_44302_23588# VPWR.t4980 pfet_06v0 ad=0.3852p pd=2.86u as=61.19999f ps=0.7u w=0.36u l=0.5u
X1637 VPWR.t4985 a_30476_23544# a_30388_23588# VPWR.t4984 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1638 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN VGND.t4719 VGND.t4718 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1639 a_51048_26680# _398_.C a_51436_27208# VGND.t3156 nfet_06v0 ad=0.1606p pd=1.61u as=58.39999f ps=0.685u w=0.365u l=0.6u
X1640 uo_out[5].t8 _287_.A1.t15 VGND.t6482 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1641 a_52452_21236# _427_.A2 _427_.ZN VGND.t718 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1642 a_28804_27208# _352_.A2.t21 VGND.t6667 VGND.t3432 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1643 VPWR.t5349 a_61164_20408# a_61076_20452# VPWR.t5348 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1644 a_44028_22020# _305_.A2 VPWR.t3021 VPWR.t3020 pfet_06v0 ad=0.4599p pd=1.935u as=0.3766p ps=1.815u w=1.095u l=0.5u
X1645 a_22188_30951# a_22100_31048# VGND.t5177 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1646 a_28596_27916.t11 _350_.A1.t6 _352_.A2.t11 VPWR.t6623 pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X1647 a_58588_11000# a_58500_11044# VGND.t5187 VGND.t5186 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1648 VPWR.t2016 a_1468_29816# a_1380_29860# VPWR.t2015 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1649 VPWR.t5362 a_65084_1592# a_64996_1636# VPWR.t5361 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1650 a_23872_27599# a_21652_27591.t4 a_23627_27967# VGND.t99 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1651 a_65084_1159# a_64996_1256# VGND.t5859 VGND.t5858 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1652 VPWR.t1949 a_20379_29977# a_20672_30301# VPWR.t1948 pfet_06v0 ad=0.38575p pd=1.92u as=0.2457p ps=1.465u w=0.945u l=0.5u
X1653 _407_.A1 _397_.A2.t7 VGND.t6720 VGND.t6719 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1654 a_40092_27209# _442_.ZN a_39968_26841# VPWR.t2940 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X1655 a_34276_23705# a_32964_24072.t3 a_33932_24073# VPWR.t153 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X1656 _250_.ZN _250_.B VGND.t2383 VGND.t2382 nfet_06v0 ad=0.21175p pd=1.41u as=0.1209p ps=0.985u w=0.465u l=0.6u
X1657 a_62508_13703# a_62420_13800# VGND.t5931 VGND.t5930 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1658 VPWR.t6195 a_1468_26680# a_1380_26724# VPWR.t657 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1659 a_31920_29480# a_31508_29159.t5 VPWR.t97 VPWR.t96 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1660 a_1468_2727# a_1380_2824# VGND.t5933 VGND.t1292 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1661 VGND.t506 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I VGND.t505 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1662 _389_.ZN _397_.A2.t8 VGND.t6722 VGND.t6721 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1663 a_55900_1592# a_55812_1636# VGND.t532 VGND.t531 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1664 VGND.t6384 _355_.C.t6 _355_.ZN VGND.t6383 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X1665 VPWR.t5096 a_43824_18147# a_43796_18559# VPWR.t5095 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X1666 VGND.t3081 a_50384_19204# a_50280_19369# VGND.t3080 nfet_06v0 ad=0.2637p pd=1.825u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1667 a_55788_24679# a_55700_24776# VGND.t4942 VGND.t2074 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1668 _251_.A1.t7 a_63616_31128# VGND.t5884 VGND.t5880 nfet_06v0 ad=0.1183p pd=0.975u as=0.23432p ps=1.94u w=0.455u l=0.6u
X1669 _325_.B _324_.B.t22 VPWR.t6708 VPWR.t2951 pfet_06v0 ad=0.4016p pd=1.94u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1670 a_47173_27208# _402_.A1.t11 VGND.t6435 VGND.t6434 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1671 VPWR.t3508 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I _241_.I0 VPWR.t3507 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1672 VPWR.t3676 a_57020_23111# a_56932_23208# VPWR.t3675 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1673 a_16140_23544# a_16052_23588# VGND.t720 VGND.t719 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1674 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I VPWR.t3339 VPWR.t3338 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1675 VGND.t5909 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I VGND.t5908 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1676 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN VGND.t882 VGND.t881 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1677 a_53696_22895# a_52920_22760# VGND.t1219 VGND.t1218 nfet_06v0 ad=43.2f pd=0.6u as=0.142p ps=1.14u w=0.36u l=0.6u
X1678 VPWR.t4281 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I VPWR.t4280 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1679 VPWR.t2660 _274_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I VPWR.t2659 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1680 VPWR.t5067 a_1916_28248# a_1828_28292# VPWR.t3269 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1681 VGND.t1427 vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I VGND.t1426 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1682 VPWR.t2488 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I VPWR.t2487 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1683 a_44290_21236# a_43814_21236# a_44038_21236# VGND.t3681 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X1684 uo_out[2].t3 _287_.A1.t16 a_37396_29860# VPWR.t6780 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1685 a_49404_14136# a_49316_14180# VGND.t4818 VGND.t4817 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1686 a_64860_18840# a_64772_18884# VGND.t5895 VGND.t3300 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1687 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN VPWR.t6165 VPWR.t6164 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1688 a_20956_23111# a_20868_23208# VGND.t5901 VGND.t5900 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1689 VPWR.t1398 a_1916_25112# a_1828_25156# VPWR.t1397 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1690 a_37360_19325# a_37067_19001# VPWR.t1332 VPWR.t1331 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X1691 a_47728_20937# a_45508_20936.t5 a_47483_20569# VGND.t190 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1692 a_13004_30951# a_12916_31048# VGND.t1318 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1693 a_49404_11000# a_49316_11044# VGND.t1332 VGND.t1331 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1694 a_21376_26031# a_20496_26344# a_21052_26031# VGND.t4669 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X1695 a_49068_20408# _419_.A4 VPWR.t4133 VPWR.t4132 pfet_06v0 ad=0.156p pd=1.12u as=0.395p ps=2.02u w=0.6u l=0.5u
X1696 VGND.t3479 a_45232_25987# a_45128_26031# VGND.t3478 nfet_06v0 ad=0.2637p pd=1.825u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1697 a_49104_30345# a_48104_30219# VGND.t2315 VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=0.142p ps=1.14u w=0.36u l=0.6u
X1698 a_58476_12135# a_58388_12232# VGND.t1344 VGND.t1343 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1699 VGND.t2959 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I VGND.t2958 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1700 a_19744_30301# a_19372_30345# VPWR.t1355 VPWR.t1354 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X1701 a_33396_26344# _358_.A3 VPWR.t478 VPWR.t477 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X1702 _362_.B.t3 a_33776_29123# VGND.t3380 VGND.t3379 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1703 VGND.t6199 _459_.CLK.t22 a_28820_30344.t1 VGND.t139 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1704 VPWR.t5743 a_1468_17272# a_1380_17316# VPWR.t2413 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1705 a_38308_18559# a_36996_18183.t5 a_37964_18191# VPWR.t6942 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X1706 a_31260_18840# a_31172_18884# VGND.t5537 VGND.t3866 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1707 VPWR.t2330 a_4604_18840# a_4516_18884# VPWR.t2329 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1708 VGND.t271 a_44296_24393.t21 clkbuf_1_0__f_clk.I.t29 VGND.t270 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1709 VGND.t3204 _301_.A1 _316_.A3 VGND.t3203 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1710 a_30812_2727# a_30724_2824# VGND.t2230 VGND.t2229 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1711 VPWR.t3831 a_43814_21236# a_44270_21790# VPWR.t3830 pfet_06v0 ad=0.379p pd=2.37u as=61.19999f ps=0.7u w=0.36u l=0.5u
X1712 a_28596_27916.t2 _350_.A2.t22 _352_.A2.t2 VPWR.t6575 pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X1713 VPWR.t1734 a_4604_15704# a_4516_15748# VPWR.t1733 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1714 VPWR.t1736 a_15692_23544# a_15604_23588# VPWR.t1735 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1715 uo_out[4].t11 _294_.ZN.t4 VGND.t147 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1716 VPWR.t2881 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN VPWR.t2880 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1717 _293_.A2 _334_.A1 a_37968_31048# VPWR.t2360 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1718 a_28928_29123# a_28556_29167# VPWR.t1618 VPWR.t1617 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X1719 VPWR.t3439 a_24316_2727# a_24228_2824# VPWR.t3438 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1720 a_53884_1592# a_53796_1636# VGND.t1691 VGND.t1690 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1721 a_58924_13703# a_58836_13800# VGND.t1693 VGND.t1692 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1722 a_4828_1159# a_4740_1256# VGND.t2203 VGND.t2202 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1723 a_46156_16839# a_46068_16936# VGND.t2205 VGND.t2204 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1724 _470_.D _404_.A1 a_44961_27912# VPWR.t3826 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1725 a_20956_1159# a_20868_1256# VGND.t5965 VGND.t5964 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1726 a_12444_1159# a_12356_1256# VGND.t5967 VGND.t5966 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1727 VGND.t1010 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I VGND.t1009 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1728 a_17803_26841# a_16240_26795# a_17168_27165# VGND.t5415 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1729 a_34160_20523# a_33748_20936.t3 VGND.t41 VGND.t40 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1730 a_60604_27815# a_60516_27912# VGND.t2766 VGND.t2765 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1731 VPWR.t5389 a_18044_2727# a_17956_2824# VPWR.t5388 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1732 VPWR.t1874 _244_.Z a_60276_26724# VPWR.t1873 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1733 VPWR.t4993 _302_.Z _324_.B.t15 VPWR.t4992 pfet_06v0 ad=0.3766p pd=1.815u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1734 VGND.t5149 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I VGND.t5148 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1735 a_54864_22461.t1 _474_.CLK.t37 VGND.t6451 VGND.t6450 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1736 a_21396_26399# a_20084_26023.t5 a_21052_26031# VPWR.t7004 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X1737 _407_.ZN _407_.A1 a_51317_27508# VGND.t526 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1738 _402_.A1.t2 a_43736_25896# VGND.t3957 VGND.t3956 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1739 a_41460_22020# _452_.Q.t9 VPWR.t6953 VPWR.t6952 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1740 VPWR.t5135 a_45372_13703# a_45284_13800# VPWR.t3037 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1741 a_60524_25640# _251_.A1.t11 a_60212_25156# VGND.t6686 nfet_06v0 ad=98.39999f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1742 a_43564_27209# _470_.D a_43396_27209# VGND.t5323 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X1743 a_21628_28248# a_21540_28292# VGND.t1619 VGND.t1618 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1744 VPWR.t1701 a_30364_1159# a_30276_1256# VPWR.t1700 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1745 a_55340_25112# a_55252_25156# VGND.t1623 VGND.t1622 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1746 a_59163_30644# a_58687_31220# a_58911_30644# VGND.t45 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X1747 a_67212_10567# a_67124_10664# VGND.t2790 VGND.t2789 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1748 a_29028_24072# _336_.A1 a_28820_24072# VGND.t4057 nfet_06v0 ad=58.39999f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X1749 a_67436_18407# a_67348_18504# VGND.t1638 VGND.t1637 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1750 a_61724_19975# a_61636_20072# VGND.t1640 VGND.t1639 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1751 a_4156_10567# a_4068_10664# VGND.t1642 VGND.t1641 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1752 VPWR.t2946 a_54332_1159# a_54244_1256# VPWR.t2945 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1753 VPWR.t935 a_61052_26247# a_60964_26344# VPWR.t934 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1754 a_31372_23544# a_31284_23588# VGND.t2811 VGND.t2810 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1755 VPWR.t1758 a_1020_4295# a_932_4392# VPWR.t1757 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1756 a_44500_25156# _304_.B _284_.ZN.t12 VPWR.t4697 pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X1757 a_56012_10567# a_55924_10664# VGND.t1677 VGND.t1676 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1758 a_48060_18407# a_47972_18504# VGND.t2718 VGND.t2717 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1759 VPWR.t2856 a_63292_9432# a_63204_9476# VPWR.t2855 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1760 VPWR.t2860 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN VPWR.t2859 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1761 a_20172_23544# a_20084_23588# VGND.t1441 VGND.t1440 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1762 VPWR.t1508 a_1020_1159# a_932_1256# VPWR.t1507 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1763 VPWR.t1510 a_47836_15704# a_47748_15748# VPWR.t1509 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1764 VPWR.t5754 a_48060_1159# a_47972_1256# VPWR.t3127 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1765 a_63068_17272# a_62980_17316# VGND.t5548 VGND.t3919 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1766 a_44296_24393.t2 clk.t2 VPWR.t6833 VPWR.t6832 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1767 a_64636_14136# a_64548_14180# VGND.t5559 VGND.t5558 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1768 VGND.t2097 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN VGND.t2096 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1769 VPWR.t5771 a_54556_14136# a_54468_14180# VPWR.t5770 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1770 VPWR.t5773 a_36636_15704# a_36548_15748# VPWR.t5772 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1771 VGND.t1771 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_62796_25640# VGND.t1770 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X1772 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN VPWR.t2182 VPWR.t2181 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1773 VPWR.t941 a_62172_15271# a_62084_15368# VPWR.t940 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1774 VGND.t253 clkbuf_1_0__f_clk.I.t38 a_48272_25156.t12 VGND.t252 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1775 a_43008_26795# a_42596_27208.t4 VGND.t145 VGND.t144 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1776 VGND.t2322 _393_.A3 _393_.ZN VGND.t2321 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X1777 a_64636_11000# a_64548_11044# VGND.t2324 VGND.t2323 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1778 VPWR.t2452 a_54556_11000# a_54468_11044# VPWR.t2451 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1779 VPWR.t1707 a_67324_12568# a_67236_12612# VPWR.t1706 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1780 VPWR.t1711 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN VPWR.t1710 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1781 _335_.ZN.t5 _334_.A1 a_36828_28776# VGND.t2245 nfet_06v0 ad=0.4161p pd=1.905u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1782 a_28348_23111# a_28260_23208# VGND.t1634 VGND.t1633 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1783 a_57168_26724# a_56404_27208# a_56964_26724# VPWR.t5737 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1784 VPWR.t5742 a_45820_12135# a_45732_12232# VPWR.t3980 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1785 _335_.ZN.t11 _460_.Q VPWR.t3485 VPWR.t3484 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1786 a_52764_2727# a_52676_2824# VGND.t5671 VGND.t5670 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1787 VPWR.t611 a_37308_15271# a_37220_15368# VPWR.t610 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1788 a_56596_29861# _272_.A2 _274_.A2 VPWR.t5895 pfet_06v0 ad=0.3402p pd=1.775u as=0.37665p ps=1.835u w=1.215u l=0.5u
X1789 a_1916_3160# a_1828_3204# VGND.t5675 VGND.t3499 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1790 a_61948_1159# a_61860_1256# VGND.t2932 VGND.t2931 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1791 _384_.A3.t3 _281_.A1 a_51618_22504# VGND.t3148 nfet_06v0 ad=0.2132p pd=1.34u as=0.1517p ps=1.19u w=0.82u l=0.6u
X1792 VPWR.t802 a_3708_13703# a_3620_13800# VPWR.t801 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1793 VPWR.t1658 a_14796_21543# a_14708_21640# VPWR.t1657 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1794 VPWR.t5843 a_7516_1159# a_7428_1256# VPWR.t5842 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1795 a_24864_29931# a_24452_30344.t4 VGND.t156 VGND.t139 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1796 a_58028_18840# a_57940_18884# VGND.t5620 VGND.t5619 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1797 _412_.ZN _424_.B1.t9 a_51540_24776# VPWR.t6617 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1798 VGND.t3001 a_45904_30180# a_45800_30345# VGND.t137 nfet_06v0 ad=0.2637p pd=1.825u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1799 a_22620_27599# _454_.D a_22452_27599# VGND.t5958 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X1800 a_16628_27209# a_15828_27208.t2 VGND.t6102 VGND.t6101 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1801 a_63516_15704# a_63428_15748# VGND.t5094 VGND.t5093 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1802 a_5052_17272# a_4964_17316# VGND.t1668 VGND.t1667 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1803 a_53660_21543# a_53572_21640# VGND.t1670 VGND.t1669 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1804 _447_.Q.t0 a_36016_20893# VPWR.t1752 VPWR.t1751 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1805 a_48308_23588# _397_.Z _399_.A2 VPWR.t896 pfet_06v0 ad=0.2964p pd=1.66u as=0.2964p ps=1.66u w=1.14u l=0.5u
X1806 VPWR.t212 _330_.A1.t10 a_44961_27912# VPWR.t211 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1807 VPWR.t5875 a_45596_1592# a_45508_1636# VPWR.t5874 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1808 a_44300_19001# a_43784_19369# VPWR.t2695 VPWR.t2694 pfet_06v0 ad=43.2f pd=0.6u as=0.1044p ps=0.94u w=0.36u l=0.5u
X1809 VPWR.t5877 a_39772_20408# a_39684_20452# VPWR.t5876 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1810 a_44160_29123# a_43788_29167# VPWR.t5086 VPWR.t5085 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X1811 a_52316_15704# a_52228_15748# VGND.t1415 VGND.t1414 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1812 a_65072_29860# rst_n.t0 VPWR.t6342 VPWR.t6341 pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X1813 VPWR.t248 clkbuf_1_0__f_clk.I.t39 a_42392_22825.t6 VPWR.t247 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1814 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN VGND.t2997 VGND.t2996 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1815 VPWR.t230 _304_.ZN.t14 _324_.B.t18 VPWR.t229 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1816 _393_.A1 _384_.ZN a_47733_29098# VGND.t3023 nfet_06v0 ad=0.21175p pd=1.41u as=85.2f ps=0.95u w=0.71u l=0.6u
X1817 a_45696_20072# a_45284_19751.t2 VGND.t6712 VGND.t6711 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1818 a_63404_23111# a_63316_23208# VGND.t5122 VGND.t5121 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1819 VGND.t1608 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I VGND.t1607 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1820 a_61388_16839# a_61300_16936# VGND.t5123 VGND.t3024 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1821 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I VGND.t1666 VGND.t1665 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1822 VPWR.t2428 a_64972_26680# a_64884_26724# VPWR.t2427 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1823 a_62956_13703# a_62868_13800# VGND.t2308 VGND.t2307 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1824 a_20060_24679# a_19972_24776# VGND.t2310 VGND.t2309 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1825 a_32592_25227# a_32180_25640.t2 VPWR.t38 VPWR.t37 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1826 VPWR.t4041 a_33164_24679# a_33076_24776# VPWR.t4040 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1827 a_53436_9432# a_53348_9476# VGND.t1433 VGND.t1432 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1828 VPWR.t1500 a_25548_20408# a_25460_20452# VPWR.t1499 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1829 a_32508_30644# _334_.A1 _370_.B VGND.t34 nfet_06v0 ad=0.1312p pd=1.14u as=0.2569p ps=1.56u w=0.82u l=0.6u
X1830 a_20060_21543# a_19972_21640# VGND.t5526 VGND.t5525 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1831 a_1468_15271# a_1380_15368# VGND.t5527 VGND.t2106 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1832 VGND.t198 _416_.A1.t6 _416_.ZN VGND.t197 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X1833 _230_.I.t1 a_61860_30736# VGND.t5456 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1834 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN VGND.t1326 VGND.t1325 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1835 a_1468_12135# a_1380_12232# VGND.t5111 VGND.t1908 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1836 a_47164_9432# a_47076_9476# VGND.t5112 VGND.t3703 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1837 VPWR.t4382 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I _248_.B1 VPWR.t4381 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1838 a_44906_24164# a_44786_24120# a_44162_24120# VGND.t1700 nfet_06v0 ad=43.2f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1839 a_37532_25112# a_37444_25156# VGND.t1701 VGND.t493 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1840 VPWR.t1653 a_4156_27815# a_4068_27912# VPWR.t484 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1841 a_53324_12135# a_53236_12232# VGND.t1577 VGND.t1576 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1842 a_46580_28292# _393_.A1 _393_.ZN VPWR.t1490 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1843 VPWR.t5534 a_5052_6296# a_4964_6340# VPWR.t5533 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1844 a_8636_1159# a_8548_1256# VGND.t5341 VGND.t5340 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1845 a_48284_17272# a_48196_17316# VGND.t5343 VGND.t5342 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1846 a_24652_30951# a_24564_31048# VGND.t1582 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1847 a_34084_28776# _362_.B.t8 a_36420_28776# VGND.t6253 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1848 a_24764_1159# a_24676_1256# VGND.t1584 VGND.t1583 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1849 a_49852_14136# a_49764_14180# VGND.t5518 VGND.t2351 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1850 a_16252_1159# a_16164_1256# VGND.t5520 VGND.t5519 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1851 VPWR.t5729 a_51868_15704# a_51780_15748# VPWR.t5728 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1852 VPWR.t5286 a_45820_9432# a_45732_9476# VPWR.t5285 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1853 VPWR.t5288 a_5052_3160# a_4964_3204# VPWR.t5287 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1854 a_4940_13703# a_4852_13800# VGND.t5120 VGND.t5119 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1855 a_37084_17272# a_36996_17316# VGND.t2317 VGND.t2316 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1856 VPWR.t2444 a_24428_21976# a_24340_22020# VPWR.t2443 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1857 a_13452_30951# a_13364_31048# VGND.t2320 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1858 a_49852_11000# a_49764_11044# VGND.t1211 VGND.t1210 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1859 VGND.t6241 _284_.ZN.t24 uo_out[1].t4 VGND.t6240 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1860 _434_.ZN _448_.Q.t4 VPWR.t6884 VPWR.t6883 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X1861 a_1916_13703# a_1828_13800# VGND.t1215 VGND.t1214 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1862 VPWR.t3504 a_22300_2727# a_22212_2824# VPWR.t3503 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1863 a_52204_16839# a_52116_16936# VGND.t5681 VGND.t5680 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1864 VGND.t5685 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I VGND.t5684 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1865 VPWR.t6374 _311_.A2.t3 a_34586_23208# VPWR.t6373 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1866 _375_.Z a_20003_29611# VPWR.t6066 VPWR.t6065 pfet_06v0 ad=0.5368p pd=3.32u as=0.38705p ps=2.08u w=1.22u l=0.5u
X1867 a_26332_1592# a_26244_1636# VGND.t5539 VGND.t5538 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1868 a_41004_16839# a_40916_16936# VGND.t5541 VGND.t5540 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1869 a_52415_31220# a_51791_30644# a_52267_30644# VGND.t45 nfet_06v0 ad=0.369p pd=2.77u as=43.2f ps=0.6u w=0.36u l=0.6u
X1870 a_39264_18147# a_38971_18559# VGND.t1705 VGND.t1704 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X1871 VPWR.t1636 a_31820_25112# a_31732_25156# VPWR.t1635 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1872 vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I VGND.t1558 VGND.t1557 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1873 a_42168_25640.t9 _284_.B a_42784_25640# VGND.t5392 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1874 a_14796_27815# a_14708_27912# VGND.t5561 VGND.t2065 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1875 _371_.A2 _455_.Q.t4 VPWR.t6849 VPWR.t6848 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1876 VPWR.t5776 a_20620_25112# a_20532_25156# VPWR.t5775 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1877 a_48732_15704# a_48644_15748# VGND.t5358 VGND.t5357 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1878 a_42168_22504# _302_.Z a_42784_22504# VGND.t4845 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1879 a_41872_28409# a_41440_28363# VPWR.t1521 VPWR.t1520 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X1880 VGND.t3823 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN VGND.t3822 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1881 a_37532_15704# a_37444_15748# VGND.t5360 VGND.t5359 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1882 VPWR.t3405 a_4156_18407# a_4068_18504# VPWR.t1075 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1883 VGND.t1269 a_17803_26841# a_18096_27165# VGND.t1268 nfet_06v0 ad=0.2608p pd=1.455u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1884 VPWR.t1471 a_30812_18407# a_30724_18504# VPWR.t1081 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1885 a_43296_28733# a_43003_28409# VGND.t1573 VGND.t1572 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X1886 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN VPWR.t5528 VPWR.t5527 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1887 a_53884_20408# a_53796_20452# VGND.t2328 VGND.t2327 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1888 VPWR.t6530 _362_.B.t9 _371_.A1.t7 VPWR.t6529 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1889 clkbuf_1_0__f_clk.I.t28 a_44296_24393.t22 VGND.t273 VGND.t272 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1890 a_42161_24776# _264_.B VPWR.t2458 VPWR.t2457 pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X1891 a_35874_27937# _334_.A1 _365_.ZN VPWR.t2359 pfet_06v0 ad=0.55297p pd=2.105u as=0.31207p ps=1.665u w=1.095u l=0.5u
X1892 a_65756_1159# a_65668_1256# VGND.t5552 VGND.t5551 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1893 a_32828_21543# a_32740_21640# VGND.t5554 VGND.t5553 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1894 a_51048_26680# _384_.A3.t10 VPWR.t182 VPWR.t181 pfet_06v0 ad=0.156p pd=1.12u as=0.40575p ps=2.055u w=0.6u l=0.5u
X1895 VPWR.t1523 a_5388_21543# a_5300_21640# VPWR.t1522 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1896 a_33932_24073# _313_.ZN a_33808_23705# VPWR.t1033 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X1897 VPWR.t1527 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN _249_.A2 VPWR.t1526 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1898 VPWR.t4141 a_10876_1159# a_10788_1256# VPWR.t4140 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1899 a_63313_28776# _229_.I.t5 VGND.t6563 VGND.t6562 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1900 VPWR.t511 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I VPWR.t510 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1901 a_60828_1592# a_60740_1636# VGND.t1686 VGND.t1685 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1902 VGND.t5102 _255_.ZN a_57500_30344# VGND.t325 nfet_06v0 ad=0.3124p pd=2.3u as=85.2f ps=0.95u w=0.71u l=0.6u
X1903 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[1\].I VGND.t1353 VGND.t1352 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1904 a_49740_12135# a_49652_12232# VGND.t5104 VGND.t5103 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1905 a_67660_10567# a_67572_10664# VGND.t5106 VGND.t5105 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1906 VPWR.t250 clkbuf_1_0__f_clk.I.t40 a_48272_25156.t6 VPWR.t249 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1907 a_67884_18407# a_67796_18504# VGND.t1592 VGND.t1591 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1908 a_67100_18840# a_67012_18884# VGND.t1594 VGND.t1593 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1909 VPWR.t5715 a_48508_9432# a_48420_9476# VPWR.t5714 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1910 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t5515 VGND.t71 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1911 VPWR.t6898 uio_out[5].t8 _379_.A2 VPWR.t6897 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1912 VPWR.t6323 a_50524_2727# a_50436_2824# VPWR.t6322 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1913 VPWR.t4724 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I VPWR.t4723 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1914 a_4156_29816# a_4068_29860# VGND.t5555 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1915 a_56460_10567# a_56372_10664# VGND.t5557 VGND.t5556 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1916 a_35516_15271# a_35428_15368# VGND.t1469 VGND.t1468 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1917 a_65196_23544# a_65108_23588# VGND.t1471 VGND.t1470 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1918 a_51956_26183# a_52360_26355# a_52304_26399# VPWR.t3285 pfet_06v0 ad=0.1665p pd=1.285u as=50.4f ps=0.64u w=0.36u l=0.5u
X1919 a_46716_12135# a_46628_12232# VGND.t6059 VGND.t1339 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1920 a_56684_18407# a_56596_18504# VGND.t6060 VGND.t2035 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1921 a_32096_24419# a_31803_24831# VGND.t3003 VGND.t3002 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X1922 _287_.A2 _459_.Q.t5 VGND.t6652 VGND.t102 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1923 a_25212_2727# a_25124_2824# VGND.t6062 VGND.t6061 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1924 VPWR.t5736 a_28572_1159# a_28484_1256# VPWR.t3691 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1925 a_52944_19759# a_52408_19759# VGND.t2605 VGND.t2604 nfet_06v0 ad=43.2f pd=0.6u as=0.2637p ps=1.825u w=0.36u l=0.6u
X1926 a_50084_24328# _281_.ZN.t7 VGND.t124 VGND.t123 nfet_06v0 ad=0.14p pd=1.1u as=0.224p ps=1.52u w=0.4u l=0.6u
X1927 VPWR.t1574 a_36636_26247# a_36548_26344# VPWR.t1573 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1928 a_50384_19204# a_49896_18909# a_50816_19369# VGND.t5242 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X1929 a_19724_25112# a_19636_25156# VGND.t5114 VGND.t5113 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1930 a_39333_20936# _300_.A2 VGND.t939 VGND.t938 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1931 a_65084_30951# a_64996_31048# VGND.t5115 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1932 VPWR.t3133 a_44252_2727# a_44164_2824# VPWR.t3132 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1933 VPWR.t5749 a_14236_29383# a_14148_29480# VPWR.t1547 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1934 a_19724_21976# a_19636_22020# VGND.t5545 VGND.t5544 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1935 VPWR.t3382 a_47164_10567# a_47076_10664# VPWR.t3381 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1936 VPWR.t5753 a_27004_27815# a_26916_27912# VPWR.t5752 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1937 VPWR.t1646 a_67772_12568# a_67684_12612# VPWR.t1645 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1938 VPWR.t6242 a_25436_23111# a_25348_23208# VPWR.t6241 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1939 VGND.t6201 _459_.CLK.t23 a_23892_27208.t1 VGND.t6200 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1940 a_28796_23111# a_28708_23208# VGND.t1568 VGND.t1567 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1941 VPWR.t11 ui_in[7].t1 a_54432_31128# VPWR.t10 pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1942 a_37420_16839# a_37332_16936# VGND.t5550 VGND.t5549 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1943 a_29563_29535# a_27588_29159.t4 a_28928_29123# VPWR.t6865 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X1944 VPWR.t3653 a_37756_15271# a_37668_15368# VPWR.t3652 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1945 _319_.A2 _317_.A2 VGND.t2452 VGND.t2451 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1946 _371_.A2 _349_.A4 VPWR.t2561 VPWR.t2560 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1947 VPWR.t1187 a_18044_1592# a_17956_1636# VPWR.t1186 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1948 VPWR.t1189 a_3708_5863# a_3620_5960# VPWR.t1188 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1949 VPWR.t24 ui_in[1].t1 a_62532_30736# VPWR.t23 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1950 VPWR.t5647 a_45372_12568# a_45284_12612# VPWR.t3902 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1951 VPWR.t278 a_44296_24393.t23 clkbuf_1_0__f_clk.I.t10 VPWR.t277 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1952 a_51420_9432# a_51332_9476# VGND.t5453 VGND.t5452 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1953 VPWR.t3111 a_3708_2727# a_3620_2824# VPWR.t3110 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1954 VPWR.t1624 a_5388_12135# a_5300_12232# VPWR.t1623 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1955 a_25124_28776# _455_.Q.t5 a_28364_28776# VGND.t6535 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1956 VGND.t1545 a_42368_28733# a_42320_28777# VGND.t1544 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X1957 a_58476_18840# a_58388_18884# VGND.t1547 VGND.t1546 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1958 a_21424_25987# a_21052_26031# VGND.t1334 VGND.t1333 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X1959 _328_.A2 _325_.A1.t10 a_44484_19668# VGND.t6515 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1960 a_45232_25987# a_44744_26355# a_45664_26031# VGND.t6032 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X1961 VPWR.t3008 a_48384_26724# clkload0.Z VPWR.t3007 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1962 a_36384_19369# a_35504_18955# a_36060_19369# VGND.t1263 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X1963 a_63964_15704# a_63876_15748# VGND.t5654 VGND.t5653 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1964 a_4156_23544# a_4068_23588# VGND.t5655 VGND.t4832 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1965 VPWR.t5881 _441_.ZN a_40084_25156# VPWR.t5880 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1966 a_67100_3160# a_67012_3204# VGND.t5659 VGND.t5658 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1967 a_28572_1159# a_28484_1256# VGND.t5529 VGND.t5528 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1968 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN VPWR.t5886 VPWR.t5885 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1969 a_43664_17317# _325_.A2.t4 _325_.ZN VPWR.t6391 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1970 a_52764_15704# a_52676_15748# VGND.t5669 VGND.t5668 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1971 _395_.A2 a_49764_26724# VGND.t989 VGND.t988 nfet_06v0 ad=0.3608p pd=2.52u as=0.224p ps=1.52u w=0.82u l=0.6u
X1972 VPWR.t5850 a_60940_15704# a_60852_15748# VPWR.t5849 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1973 a_48708_29816# a_49152_30301.t3 a_49104_30345# VGND.t137 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X1974 VPWR.t6902 uio_out[6].t9 a_20191_29611# VPWR.t6901 pfet_06v0 ad=0.38705p pd=2.08u as=0.1469p ps=1.085u w=0.565u l=0.5u
X1975 a_36004_24463# a_35204_24455.t2 VGND.t6130 VGND.t6129 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1976 a_51457_29861# _274_.ZN VPWR.t1035 VPWR.t1034 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1977 a_30388_28776# _371_.A1.t12 _350_.A2.t11 VGND.t6232 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1978 _337_.ZN _336_.A2.t3 VPWR.t168 VPWR.t167 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1979 a_63852_23111# a_63764_23208# VGND.t1002 VGND.t1001 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1980 VPWR.t6376 _311_.A2.t4 a_34980_22895# VPWR.t6375 pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X1981 VPWR.t3543 a_49404_18407# a_49316_18504# VPWR.t3542 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1982 a_55900_14136# a_55812_14180# VGND.t3067 VGND.t3066 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1983 VPWR.t3227 a_45820_14136# a_45732_14180# VPWR.t3204 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1984 VGND.t6242 _284_.ZN.t25 a_38472_30169# VGND.t71 nfet_06v0 ad=0.2662p pd=2.09u as=0.51425p ps=2.91u w=0.605u l=0.6u
X1985 a_19612_26247# a_19524_26344# VGND.t3034 VGND.t3033 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1986 VGND.t2523 _274_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I VGND.t2522 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1987 a_55900_11000# a_55812_11044# VGND.t3036 VGND.t3035 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1988 VPWR.t3196 a_45820_11000# a_45732_11044# VPWR.t1226 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1989 VPWR.t3678 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN VPWR.t3677 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1990 _250_.ZN _251_.A1.t12 a_62503_28293# VPWR.t7011 pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X1991 a_23196_2727# a_23108_2824# VGND.t3533 VGND.t3532 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1992 _452_.CLK.t4 a_42392_22825.t18 VGND.t6601 VGND.t6600 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1993 a_19612_23111# a_19524_23208# VGND.t3535 VGND.t3534 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1994 VPWR.t3923 a_3708_12568# a_3620_12612# VPWR.t2865 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1995 a_4604_9432# a_4516_9476# VGND.t3780 VGND.t3779 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1996 VPWR.t3927 a_14796_20408# a_14708_20452# VPWR.t3926 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1997 a_64972_12135# a_64884_12232# VGND.t5627 VGND.t5626 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1998 a_47164_2727# a_47076_2824# VGND.t5629 VGND.t5628 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1999 _452_.Q.t1 a_40040_17675# VPWR.t5253 VPWR.t5252 pfet_06v0 ad=0.3172p pd=1.74u as=0.854p ps=3.84u w=1.22u l=0.5u
X2000 a_21052_26031# _455_.D a_20928_26399# VPWR.t866 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X2001 VPWR.t6344 rst_n.t1 a_65072_29860# VPWR.t6343 pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X2002 a_5388_27815# a_5300_27912# VGND.t3655 VGND.t3654 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2003 a_54108_12568# a_54020_12612# VGND.t3657 VGND.t3656 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2004 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I VPWR.t1941 VPWR.t1940 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2005 a_57244_27815# a_57156_27912# VGND.t3659 VGND.t3658 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2006 a_4604_6296# a_4516_6340# VGND.t3582 VGND.t3581 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2007 VGND.t3584 _331_.ZN _452_.D VGND.t3583 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X2008 a_53772_12135# a_53684_12232# VGND.t3586 VGND.t3585 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2009 a_22620_27599# _454_.D a_22496_27967# VPWR.t6215 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X2010 a_50748_15271# a_50660_15368# VGND.t2880 VGND.t2879 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2011 VPWR.t848 a_21740_30951# a_21652_31048# VPWR.t847 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2012 a_2812_26247# a_2724_26344# VGND.t2881 VGND.t1289 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2013 VPWR.t3030 a_17036_21543# a_16948_21640# VPWR.t2489 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2014 VPWR.t6032 a_40668_26247# a_40580_26344# VPWR.t6031 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2015 VGND.t6203 _459_.CLK.t24 a_23668_25640.t1 VGND.t6202 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2016 VPWR.t3941 a_10540_30951# a_10452_31048# VPWR.t3940 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2017 VGND.t1689 a_28928_29123# a_28880_29167# VGND.t1688 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X2018 _371_.A2 _454_.Q VPWR.t4088 VPWR.t4087 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2019 VPWR.t3510 a_24876_21976# a_24788_22020# VPWR.t3509 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2020 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN VGND.t2993 VGND.t2992 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2021 a_2812_23111# a_2724_23208# VGND.t2944 VGND.t2943 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2022 _369_.ZN _371_.A1.t13 a_29680_26724# VPWR.t6510 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X2023 VGND.t5703 _293_.A2 uo_out[1].t10 VGND.t5702 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2024 VPWR.t3103 a_65308_6296# a_65220_6340# VPWR.t3102 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2025 VPWR.t3417 a_42236_27815# a_42148_27912# VPWR.t3416 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2026 a_44795_29535# a_42820_29159.t7 a_44160_29123# VPWR.t7043 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X2027 a_52652_16839# a_52564_16936# VGND.t3274 VGND.t3273 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2028 VGND.t3278 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN VGND.t3277 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2029 VPWR.t5230 a_52988_15271# a_52900_15368# VPWR.t5229 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2030 VPWR.t42 _363_.Z.t3 a_35874_27937# VPWR.t41 pfet_06v0 ad=0.4818p pd=3.07u as=0.55297p ps=2.105u w=1.095u l=0.5u
X2031 VPWR.t3895 a_65308_3160# a_65220_3204# VPWR.t3894 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2032 VPWR.t3672 a_19035_28409# a_19328_28733# VPWR.t3671 pfet_06v0 ad=0.38575p pd=1.92u as=0.2457p ps=1.465u w=0.945u l=0.5u
X2033 VPWR.t1720 a_61724_19975# a_61636_20072# VPWR.t1719 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2034 a_34586_23208# _304_.A1.t6 _312_.ZN VPWR.t6601 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2035 VPWR.t3820 a_3260_21543# a_3172_21640# VPWR.t3819 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2036 a_41452_16839# a_41364_16936# VGND.t3671 VGND.t3670 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2037 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t5719 VPWR.t5718 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2038 a_1468_28248# a_1380_28292# VGND.t3673 VGND.t3672 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2039 a_49828_22020# _473_.Q a_49604_22020# VPWR.t5159 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2040 VPWR.t3946 a_21404_24679# a_21316_24776# VPWR.t3945 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2041 VPWR.t5765 a_4156_29816# a_4068_29860# VPWR.t3430 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2042 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN VPWR.t4143 VPWR.t4142 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2043 VPWR.t5858 a_25936_25597# a_25928_25273# VPWR.t5857 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X2044 VPWR.t4120 a_35180_16839# a_35092_16936# VPWR.t4119 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2045 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I VPWR.t5132 VPWR.t5131 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2046 VPWR.t3256 a_54444_25112# a_54356_25156# VPWR.t1441 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2047 VPWR.t3257 a_4156_26680# a_4068_26724# VPWR.t1443 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2048 _474_.CLK.t10 a_48272_25156.t24 VGND.t6268 VGND.t6267 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X2049 a_31484_1159# a_31396_1256# VGND.t3111 VGND.t3110 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2050 VPWR.t4164 a_32156_16839# a_32068_16936# VPWR.t2905 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2051 VGND.t1746 a_38336_18147# a_38288_18191# VGND.t1745 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X2052 a_37980_15704# a_37892_15748# VGND.t3627 VGND.t3626 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2053 VPWR.t4063 vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN VPWR.t4062 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2054 a_58924_17272# a_58836_17316# VGND.t3629 VGND.t3628 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2055 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I VGND.t1604 VGND.t1603 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2056 uo_out[0].t10 _284_.ZN.t26 VGND.t6243 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2057 a_52540_1592# a_52452_1636# VGND.t3007 VGND.t3006 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2058 a_27172_24328# _336_.A2.t4 VPWR.t170 VPWR.t169 pfet_06v0 ad=0.1456p pd=1.08u as=0.34437p ps=1.895u w=0.56u l=0.5u
X2059 a_2812_16839# a_2724_16936# VGND.t3008 VGND.t1497 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2060 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN VGND.t5683 VGND.t5682 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2061 a_28900_29535# a_27588_29159.t5 a_28556_29167# VPWR.t6866 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X2062 VGND.t2447 _276_.A2 a_52073_30344# VGND.t199 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2063 VPWR.t3057 a_65308_18840# a_65220_18884# VPWR.t3056 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2064 a_33720_28776# _223_.ZN VGND.t777 VGND.t776 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2065 a_30132_29977# a_28820_30344.t2 a_29788_30345# VPWR.t6365 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X2066 VPWR.t4605 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].I VPWR.t4604 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2067 a_26750_28776# _454_.Q a_26556_28776# VGND.t3940 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2068 VPWR.t1614 a_65308_15704# a_65220_15748# VPWR.t1613 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2069 VGND.t2866 a_48384_26724# clkload0.Z VGND.t2865 nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X2070 VPWR.t1211 a_4604_28248# a_4516_28292# VPWR.t1210 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2071 VPWR.t3 a_1916_7431# a_1828_7528# VPWR.t2 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2072 VGND.t1242 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t1241 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2073 a_58116_30344# _255_.ZN VGND.t5101 VGND.t71 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2074 VPWR.t5021 a_20672_30301# a_20664_29977# VPWR.t5020 pfet_06v0 ad=0.2619p pd=1.685u as=50.4f ps=0.64u w=0.36u l=0.5u
X2075 a_23644_23111# a_23556_23208# VGND.t1248 VGND.t1247 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2076 VPWR.t2388 a_4604_25112# a_4516_25156# VPWR.t2387 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2077 VGND.t1632 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN VGND.t1631 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2078 VPWR.t3952 a_32604_15271# a_32516_15368# VPWR.t3951 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2079 a_3260_8999# a_3172_9096# VGND.t2270 VGND.t2269 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2080 VPWR.t2391 a_3260_12135# a_3172_12232# VPWR.t2390 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2081 a_35964_15271# a_35876_15368# VGND.t2710 VGND.t2709 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2082 VPWR.t5050 a_48708_29816# a_48104_30219# VPWR.t5049 pfet_06v0 ad=0.23p pd=1.54u as=0.352p ps=2.48u w=0.8u l=0.5u
X2083 VGND.t1788 a_18400_28733# a_18352_28777# VGND.t1787 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X2084 a_1468_18840# a_1380_18884# VGND.t2712 VGND.t2711 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2085 a_3260_5863# a_3172_5960# VGND.t2714 VGND.t2713 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2086 VPWR.t2568 a_24764_2727# a_24676_2824# VPWR.t2567 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2087 a_33508_31048# _287_.A1.t17 uo_out[5].t5 VPWR.t6781 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2088 VPWR.t4425 a_24092_21543# a_24004_21640# VPWR.t4424 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2089 VPWR.t2738 a_51620_19911# a_51240_19624# VPWR.t2737 pfet_06v0 ad=0.23p pd=1.54u as=0.352p ps=2.48u w=0.8u l=0.5u
X2090 VPWR.t5530 a_48508_30951# a_48420_31048# VPWR.t5529 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2091 VPWR.t4426 a_14684_29383# a_14596_29480# VPWR.t655 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2092 VPWR.t2303 a_4156_17272# a_4068_17316# VPWR.t926 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2093 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN _245_.I1 VGND.t5232 VGND.t5231 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2094 VPWR.t2304 a_36188_26680# a_36100_26724# VPWR.t928 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2095 VPWR.t2305 a_30812_17272# a_30724_17316# VPWR.t930 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2096 _370_.B _223_.I VGND.t6794 VGND.t6793 nfet_06v0 ad=0.2569p pd=1.56u as=0.2244p ps=1.9u w=0.51u l=0.6u
X2097 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN VPWR.t609 VPWR.t608 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2098 VGND.t2220 a_31168_24419# a_31120_24463# VGND.t2219 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X2099 VPWR.t5267 a_18492_2727# a_18404_2824# VPWR.t5266 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2100 VPWR.t5575 a_25884_23111# a_25796_23208# VPWR.t5574 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2101 a_17036_27815# a_16948_27912# VGND.t2222 VGND.t2221 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2102 a_35044_21640# _330_.A1.t11 _316_.ZN VPWR.t213 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2103 VPWR.t6770 _359_.B.t6 a_34308_26344# VPWR.t6769 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X2104 VPWR.t5834 a_18380_23544# a_18292_23588# VPWR.t5833 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2105 VPWR.t1957 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I VPWR.t1956 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2106 VPWR.t465 a_46624_19715# a_46596_20127# VPWR.t464 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X2107 VPWR.t4154 a_26108_30951# a_26020_31048# VPWR.t4153 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2108 a_52073_30344# _416_.A1.t7 vgaringosc.workerclkbuff_notouch_.I.t0 VGND.t199 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X2109 uo_out[2].t8 _288_.ZN.t3 VGND.t6063 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X2110 VGND.t2254 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN VGND.t2253 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2111 VGND.t2798 a_54192_22851# a_54088_22895# VGND.t2797 nfet_06v0 ad=0.2637p pd=1.825u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2112 a_51420_2727# a_51332_2824# VGND.t2802 VGND.t2801 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2113 a_43888_27209# a_43008_26795# a_43564_27209# VGND.t5759 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X2114 VPWR.t2937 a_54780_1159# a_54692_1256# VPWR.t2936 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2115 VPWR.t280 a_44296_24393.t24 clkbuf_1_0__f_clk.I.t9 VPWR.t279 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2116 VPWR.t1642 a_47948_16839# a_47860_16936# VPWR.t1641 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2117 a_18268_30951# a_18180_31048# VGND.t2182 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2118 _437_.ZN _437_.A1.t9 a_37408_23208# VPWR.t6860 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X2119 a_30924_20408# a_30836_20452# VGND.t2184 VGND.t2183 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2120 VPWR.t2884 a_20844_20408# a_20756_20452# VPWR.t2883 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2121 a_3260_27815# a_3172_27912# VGND.t2752 VGND.t2751 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2122 a_55228_1592# a_55140_1636# VGND.t2754 VGND.t2753 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2123 VPWR.t2889 a_65868_12135# a_65780_12232# VPWR.t2888 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2124 VGND.t6205 _459_.CLK.t25 a_42820_29159.t0 VGND.t6204 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2125 a_28000_29480# a_27588_29159.t6 VPWR.t6868 VPWR.t6867 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2126 a_27460_28776# _337_.A3.t6 _371_.A2 VGND.t6137 nfet_06v0 ad=0.1312p pd=1.14u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2127 VPWR.t6219 a_54668_12135# a_54580_12232# VPWR.t6218 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2128 VPWR.t467 a_20284_1592# a_20196_1636# VPWR.t466 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2129 VPWR.t6221 a_36636_25112# a_36548_25156# VPWR.t6220 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2130 VPWR.t2871 a_16700_29383# a_16612_29480# VPWR.t2403 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2131 a_16140_28248# a_16052_28292# VGND.t2738 VGND.t2737 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2132 VPWR.t3567 a_48060_13703# a_47972_13800# VPWR.t3566 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2133 VPWR.t1252 a_44252_1592# a_44164_1636# VPWR.t1251 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2134 a_64412_19975# a_64324_20072# VGND.t2740 VGND.t2739 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2135 vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN VPWR.t2827 VPWR.t2826 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2136 VPWR.t2833 a_47388_17272# a_47300_17316# VPWR.t2832 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2137 a_43668_19668# _324_.B.t23 a_43444_19668# VGND.t6415 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2138 VPWR.t6269 a_27900_23111# a_27812_23208# VPWR.t6268 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2139 a_1468_30951# a_1380_31048# VGND.t2695 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2140 VPWR.t2909 a_30924_21976# a_30836_22020# VPWR.t2908 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2141 a_49404_1159# a_49316_1256# VGND.t2777 VGND.t2776 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2142 a_31140_24831# a_29828_24455.t3 a_30796_24463# VPWR.t6386 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X2143 a_38576_22504# _311_.A2.t5 VPWR.t6378 VPWR.t6377 pfet_06v0 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X2144 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t2781 VGND.t2780 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2145 VPWR.t4116 a_4940_8999# a_4852_9096# VPWR.t4115 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2146 VPWR.t2147 a_36188_17272# a_36100_17316# VPWR.t2146 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2147 VGND.t2044 a_24196_31048# uio_out[3].t0 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2148 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I _258_.ZN VGND.t2048 VGND.t2047 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2149 a_27676_2727# a_27588_2824# VGND.t2049 VGND.t1977 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2150 VPWR.t6206 a_7964_1159# a_7876_1256# VPWR.t6205 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2151 VPWR.t6997 _335_.ZN.t22 _350_.A2.t16 VPWR.t6996 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2152 VPWR.t6207 a_3708_4728# a_3620_4772# VPWR.t5464 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2153 VPWR.t5277 a_35628_18407# a_35540_18504# VPWR.t5276 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2154 a_41708_30644# _388_.B _495_.I VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2155 a_54556_12568# a_54468_12612# VGND.t5948 VGND.t5947 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2156 a_67324_14136# a_67236_14180# VGND.t2037 VGND.t968 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2157 VPWR.t2145 a_57244_14136# a_57156_14180# VPWR.t2144 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2158 a_42392_22825.t5 clkbuf_1_0__f_clk.I.t41 VPWR.t252 VPWR.t251 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X2159 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN VPWR.t4279 VPWR.t4278 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2160 VPWR.t650 a_3708_1592# a_3620_1636# VPWR.t649 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2161 a_35292_1159# a_35204_1256# VGND.t2041 VGND.t2040 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2162 VGND.t5985 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t5984 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2163 hold2.I hold1.Z a_42853_24373# VGND.t3419 nfet_06v0 ad=0.2015p pd=1.295u as=92.99999f ps=1.015u w=0.775u l=0.6u
X2164 a_22944_27599# a_22064_27912# a_22620_27599# VGND.t3268 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X2165 VGND.t6564 _229_.I.t6 a_61297_30300# VGND.t1077 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2166 a_67324_11000# a_67236_11044# VGND.t5826 VGND.t5825 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2167 VPWR.t6086 a_57244_11000# a_57156_11044# VPWR.t6085 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2168 a_41536_17636# a_41088_17757.t4 a_41948_17433# VPWR.t162 pfet_06v0 ad=0.1872p pd=1.4u as=43.2f ps=0.6u w=0.36u l=0.5u
X2169 a_60276_29032# _238_.I a_60916_29612# VPWR.t2237 pfet_06v0 ad=0.2464p pd=2u as=0.1736p ps=1.18u w=0.56u l=0.5u
X2170 VPWR.t476 _358_.A3 a_31348_25156# VPWR.t475 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2171 VPWR.t6100 a_17484_21543# a_17396_21640# VPWR.t1696 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2172 a_66988_19975# a_66900_20072# VGND.t5842 VGND.t5841 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2173 a_51665_30344# _275_.ZN VGND.t2481 VGND.t199 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2174 a_3708_1159# a_3620_1256# VGND.t1301 VGND.t1300 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2175 VPWR.t1376 a_57468_1159# a_57380_1256# VPWR.t1375 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2176 VGND.t2591 a_60212_25156# _244_.Z VGND.t2590 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2177 VPWR.t1378 a_4156_4295# a_4068_4392# VPWR.t1377 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2178 a_53884_9432# a_53796_9476# VGND.t5862 VGND.t5861 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2179 a_11324_1159# a_11236_1256# VGND.t5864 VGND.t5863 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2180 VPWR.t6126 a_42684_27815# a_42596_27912# VPWR.t6125 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2181 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN VPWR.t2366 VPWR.t2365 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2182 a_33376_23659# a_32964_24072.t4 VPWR.t155 VPWR.t154 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2183 VPWR.t406 a_18096_27165# uio_out[7].t3 VPWR.t405 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2184 a_1916_17272# a_1828_17316# VGND.t5837 VGND.t2849 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2185 a_51668_23340# _384_.A3.t11 a_51428_23340# VPWR.t183 pfet_06v0 ad=0.1736p pd=1.18u as=0.196p ps=1.26u w=0.56u l=0.5u
X2186 VGND.t6105 _311_.A2.t6 _312_.ZN VGND.t6104 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2187 a_20664_29977# a_18816_29931# a_20379_29977# VPWR.t6099 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X2188 uo_out[5].t11 _287_.A1.t18 a_33060_31048# VPWR.t6782 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2189 a_41708_30644# a_41056_30669# VGND.t5968 VGND.t34 nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X2190 VPWR.t4250 a_4156_1159# a_4068_1256# VPWR.t4249 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2191 a_1468_24679# a_1380_24776# VGND.t5969 VGND.t3343 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2192 a_66204_15704# a_66116_15748# VGND.t5971 VGND.t5970 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2193 _272_.A2 _255_.ZN VPWR.t5271 VPWR.t5270 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2194 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN VPWR.t6175 VPWR.t6174 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2195 VPWR.t2864 vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I VPWR.t2863 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2196 a_1468_21543# a_1380_21640# VGND.t5814 VGND.t2187 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2197 VGND.t6064 _288_.ZN.t4 uo_out[2].t9 VGND.t146 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2198 a_9084_29383# a_8996_29480# VGND.t5816 VGND.t5815 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2199 VPWR.t2615 a_21852_24679# a_21764_24776# VPWR.t2614 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2200 VPWR.t176 a_44784_25987.t2 a_44744_26355# VPWR.t175 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2201 a_64076_16839# a_63988_16936# VGND.t2051 VGND.t2050 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2202 VGND.t2101 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I VGND.t2100 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2203 a_45012_29816# a_45416_29885# a_45360_29977# VPWR.t2160 pfet_06v0 ad=0.1665p pd=1.285u as=50.4f ps=0.64u w=0.36u l=0.5u
X2204 VPWR.t2163 a_54892_25112# a_54804_25156# VPWR.t1143 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2205 vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN VPWR.t2879 VPWR.t2878 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2206 a_41056_30669# _388_.B VPWR.t4315 VPWR.t4314 pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X2207 VPWR.t542 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN _231_.I VPWR.t541 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2208 VPWR.t341 a_59955_30600# _237_.A1 VPWR.t340 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2209 VPWR.t3766 a_5724_30951# a_5636_31048# VPWR.t3765 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2210 a_38316_20408# a_38228_20452# VGND.t5905 VGND.t5904 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2211 VPWR.t6171 a_5276_29383# a_5188_29480# VPWR.t6170 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2212 a_4156_15271# a_4068_15368# VGND.t5972 VGND.t3444 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2213 a_13340_29383# a_13252_29480# VGND.t5974 VGND.t5973 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2214 a_27116_20408# a_27028_20452# VGND.t5976 VGND.t5975 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2215 a_50076_9432# a_49988_9476# VGND.t5978 VGND.t5977 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2216 VPWR.t2130 a_17036_20408# a_16948_20452# VPWR.t2129 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2217 a_30812_15271# a_30724_15368# VGND.t2028 VGND.t2027 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2218 a_67212_12135# a_67124_12232# VGND.t2030 VGND.t2029 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2219 a_36432_19325# a_36060_19369# VGND.t1612 VGND.t1611 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X2220 VPWR.t2137 a_30140_21543# a_30052_21640# VPWR.t2136 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2221 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I VGND.t3276 VGND.t3275 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2222 VPWR.t6211 a_18828_25112# a_18740_25156# VPWR.t6210 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2223 _370_.ZN _370_.B VGND.t5524 VGND.t5523 nfet_06v0 ad=0.21175p pd=1.41u as=0.1209p ps=0.985u w=0.465u l=0.6u
X2224 a_4156_12135# a_4068_12232# VGND.t5953 VGND.t4008 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2225 _460_.D _360_.ZN VGND.t5955 VGND.t5954 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2226 VPWR.t3493 a_31932_26247# a_31844_26344# VPWR.t3492 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2227 VPWR.t6074 a_57580_18840# a_57492_18884# VPWR.t4926 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2228 a_5052_7864# a_4964_7908# VGND.t5821 VGND.t5820 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2229 VPWR.t6078 a_65756_18840# a_65668_18884# VPWR.t6077 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2230 VGND.t2468 a_61836_25515# _245_.Z VGND.t2467 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2231 VPWR.t591 a_60268_13703# a_60180_13800# VPWR.t590 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2232 a_56012_12135# a_55924_12232# VGND.t5830 VGND.t5829 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2233 a_26780_1592# a_26692_1636# VGND.t5832 VGND.t5831 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2234 VPWR.t2067 a_38616_24328# _311_.A2.t0 VPWR.t2066 pfet_06v0 ad=0.40575p pd=2.055u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2235 a_52316_1159# a_52228_1256# VGND.t5834 VGND.t5833 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2236 a_60828_1159# a_60740_1256# VGND.t2442 VGND.t2441 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2237 VPWR.t2480 a_31932_23111# a_31844_23208# VPWR.t2479 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2238 VGND.t6139 _337_.A3.t7 a_29348_25940# VGND.t6138 nfet_06v0 ad=0.3608p pd=2.52u as=0.1148p ps=1.1u w=0.82u l=0.6u
X2239 a_65072_29860# rst_n.t2 VGND.t6072 VGND.t71 nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X2240 a_46716_30951# a_46628_31048# VGND.t5352 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2241 a_5052_4728# a_4964_4772# VGND.t5354 VGND.t5353 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2242 VPWR.t410 a_65756_15704# a_65668_15748# VPWR.t409 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2243 VPWR.t6557 a_48272_25156.t25 _474_.CLK.t11 VPWR.t6556 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2244 VPWR.t1681 a_50636_10567# a_50548_10664# VPWR.t1680 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2245 a_24428_23544# a_24340_23588# VGND.t5440 VGND.t5439 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2246 a_32980_25641# a_32180_25640.t3 VGND.t31 VGND.t30 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2247 a_33812_29860# _294_.ZN.t5 VPWR.t148 VPWR.t147 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X2248 a_33948_17272# a_33860_17316# VGND.t5442 VGND.t5441 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2249 VPWR.t5640 a_3260_20408# a_3172_20452# VPWR.t5639 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2250 VGND.t1075 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN VGND.t1074 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2251 a_36172_24463# _444_.D a_36004_24463# VGND.t5444 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X2252 _352_.A2.t10 _350_.A1.t7 a_28596_27916.t10 VPWR.t6624 pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X2253 VPWR.t5645 a_27116_21976# a_27028_22020# VPWR.t5644 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2254 a_60828_26680# a_60740_26724# VGND.t5179 VGND.t5178 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2255 VPWR.t5940 a_66428_15271# a_66340_15368# VPWR.t5939 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2256 VPWR.t5354 a_32156_18840# a_32068_18884# VPWR.t4443 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2257 VPWR.t3993 _359_.ZN _360_.ZN VPWR.t3992 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X2258 VPWR.t1744 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I VPWR.t1743 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2259 a_48921_22020# _473_.Q VPWR.t5158 VPWR.t5157 pfet_06v0 ad=0.1469p pd=1.085u as=0.38705p ps=2.08u w=0.565u l=0.5u
X2260 a_39884_27815# a_39796_27912# VGND.t5183 VGND.t5182 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2261 a_33956_31048# _290_.ZN VPWR.t1205 VPWR.t1204 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2262 VPWR.t5677 a_67100_7431# a_67012_7528# VPWR.t5034 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2263 VPWR.t5890 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN VPWR.t5889 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2264 VGND.t5369 _327_.Z a_40636_18180# VGND.t5368 nfet_06v0 ad=0.2424p pd=1.635u as=79.8f ps=0.8u w=0.38u l=0.6u
X2265 VPWR.t2981 a_32156_15704# a_32068_15748# VPWR.t1974 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2266 a_25204_26841# a_23892_27208.t2 a_24860_27209# VPWR.t6337 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X2267 VPWR.t2969 a_48956_30951# a_48868_31048# VPWR.t2968 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2268 _359_.B.t1 a_45088_29123# VGND.t4295 VGND.t4294 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2269 a_19035_28409# a_17472_28363# a_18400_28733# VGND.t2503 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2270 VPWR.t5542 a_60716_12135# a_60628_12232# VPWR.t5541 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2271 VPWR.t3704 a_44028_15271# a_43940_15368# VPWR.t3703 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2272 a_47388_15271# a_47300_15368# VGND.t5349 VGND.t5348 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2273 a_17484_27815# a_17396_27912# VGND.t5351 VGND.t5350 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2274 a_21052_26031# _455_.D a_20884_26031# VGND.t847 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X2275 a_52848_25987# a_52400_25987.t3 a_53260_26399# VPWR.t6371 pfet_06v0 ad=0.1872p pd=1.4u as=43.2f ps=0.6u w=0.36u l=0.5u
X2276 a_1020_25112# a_932_25156# VGND.t5171 VGND.t2175 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2277 a_2812_7431# a_2724_7528# VGND.t5172 VGND.t2086 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2278 VPWR.t5347 a_45260_17272# a_45172_17316# VPWR.t1978 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2279 vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t1240 VGND.t1239 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2280 VPWR.t2585 a_26556_30951# a_26468_31048# VPWR.t2584 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2281 a_31932_2727# a_31844_2824# VGND.t3338 VGND.t3337 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2282 VPWR.t3488 a_1916_9432# a_1828_9476# VPWR.t1981 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2283 VPWR.t1518 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I VPWR.t1517 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2284 VGND.t322 a_9635_30644# a_9635_30644# VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2285 VPWR.t3753 _267_.A2 _267_.ZN VPWR.t3752 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X2286 a_1020_21976# a_932_22020# VGND.t3831 VGND.t2681 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2287 VPWR.t333 a_42996_18840# a_42392_19243# VPWR.t332 pfet_06v0 ad=0.23p pd=1.54u as=0.352p ps=2.48u w=0.8u l=0.5u
X2288 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN VGND.t1630 VGND.t1629 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2289 a_2812_26680# a_2724_26724# VGND.t3832 VGND.t2683 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2290 VPWR.t2749 a_50972_2727# a_50884_2824# VPWR.t2748 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2291 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t724 VGND.t723 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2292 VPWR.t3757 a_3260_14136# a_3172_14180# VPWR.t3756 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2293 VPWR.t2792 a_33500_18407# a_33412_18504# VPWR.t2791 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2294 a_25660_2727# a_25572_2824# VGND.t3620 VGND.t3619 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2295 a_49292_16839# a_49204_16936# VGND.t3622 VGND.t3621 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2296 a_57468_16839# a_57380_16936# VGND.t3624 VGND.t3623 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2297 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I VPWR.t2205 VPWR.t2204 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2298 a_17472_28363# a_17060_28776.t4 VPWR.t6906 VPWR.t6905 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2299 VPWR.t3368 a_3260_11000# a_3172_11044# VPWR.t1987 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2300 a_16140_24679# a_16052_24776# VGND.t3222 VGND.t719 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2301 a_35268_21640# _317_.A2 a_35044_21640# VPWR.t2577 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2302 VPWR.t1963 a_49404_2727# a_49316_2824# VPWR.t1962 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2303 a_29468_1592# a_29380_1636# VGND.t3223 VGND.t3126 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2304 a_7516_1159# a_7428_1256# VGND.t5618 VGND.t5617 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2305 VPWR.t5123 a_60401_30300# _255_.I VPWR.t5122 pfet_06v0 ad=0.38705p pd=2.08u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2306 VPWR.t3838 a_5388_4295# a_5300_4392# VPWR.t3837 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2307 a_49952_26724# _412_.A1 a_49764_26724# VPWR.t3841 pfet_06v0 ad=0.1736p pd=1.18u as=0.2464p ps=2u w=0.56u l=0.5u
X2308 a_15132_1159# a_15044_1256# VGND.t3693 VGND.t3692 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2309 a_53108_21640# _422_.ZN _427_.ZN VPWR.t2004 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2310 a_16140_21543# a_16052_21640# VGND.t2846 VGND.t2200 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2311 VPWR.t6469 _459_.CLK.t26 a_35316_29159.t0 VPWR.t6468 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2312 VPWR.t4081 a_2364_8999# a_2276_9096# VPWR.t4000 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2313 VPWR.t2985 a_32268_20408# a_32180_20452# VPWR.t2984 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2314 a_62564_29032# _230_.I.t4 a_62944_29101# VGND.t6345 nfet_06v0 ad=0.1584p pd=1.6u as=57.59999f ps=0.68u w=0.36u l=0.6u
X2315 a_64860_19975# a_64772_20072# VGND.t3301 VGND.t3300 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2316 a_47636_25940# _397_.A1.t6 _284_.B VGND.t9 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2317 VPWR.t3667 _296_.ZN a_40644_31048# VPWR.t3666 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2318 VPWR.t3222 _378_.I _378_.ZN VPWR.t3221 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2319 a_43668_19668# _325_.A2.t5 _325_.B VGND.t6122 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2320 a_19500_27815# a_19412_27912# VGND.t3304 VGND.t3303 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2321 VPWR.t1191 a_18492_1592# a_18404_1636# VPWR.t1190 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2322 VPWR.t3259 a_31484_1159# a_31396_1256# VPWR.t3258 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2323 a_52852_24372# _428_.Z VGND.t4759 VGND.t4758 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2324 VGND.t5770 a_43888_19204# a_43784_19369# VGND.t5769 nfet_06v0 ad=0.2637p pd=1.825u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2325 a_41488_24072# _260_.A1 VPWR.t3916 VPWR.t3915 pfet_06v0 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X2326 VPWR.t3918 a_20508_21543# a_20420_21640# VPWR.t3917 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2327 _352_.A2.t1 _350_.A2.t23 a_28596_27916.t1 VPWR.t6576 pfet_06v0 ad=0.312p pd=1.72u as=0.48p ps=2u w=1.2u l=0.5u
X2328 VPWR.t5019 a_20672_30301# uio_out[5].t2 VPWR.t5018 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2329 VPWR.t6076 a_5052_7864# a_4964_7908# VPWR.t6075 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2330 VPWR.t3971 a_39324_26247# a_39236_26344# VPWR.t3970 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2331 a_1020_15704# a_932_15748# VGND.t4043 VGND.t3970 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2332 a_67772_14136# a_67684_14180# VGND.t4044 VGND.t3921 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2333 VPWR.t765 a_61164_23111# a_61076_23208# VPWR.t764 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2334 a_26756_24801# _352_.A2.t22 VPWR.t6989 VPWR.t6988 pfet_06v0 ad=0.55297p pd=2.105u as=0.4818p ps=3.07u w=1.095u l=0.5u
X2335 VPWR.t4019 a_57692_14136# a_57604_14180# VPWR.t4018 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2336 a_44864_27165# a_44571_26841# VGND.t2821 VGND.t2820 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X2337 a_51196_1592# a_51108_1636# VGND.t3865 VGND.t3864 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2338 a_31260_19975# a_31172_20072# VGND.t3867 VGND.t3866 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2339 a_35716_20072# _319_.A2 a_35492_20072# VPWR.t1185 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2340 VPWR.t6060 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t6059 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2341 a_29620_30345# a_28820_30344.t3 VGND.t6094 VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2342 a_11100_29816# a_11012_29860# VGND.t3167 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2343 VPWR.t2250 a_58028_10567# a_57940_10664# VPWR.t2249 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2344 _424_.A2.t3 _324_.C.t15 VPWR.t6798 VPWR.t6797 pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X2345 VPWR.t3316 a_60940_28248# a_60852_28292# VPWR.t3315 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2346 a_67772_11000# a_67684_11044# VGND.t3171 VGND.t3170 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2347 a_3708_20408# a_3620_20452# VGND.t2884 VGND.t2883 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2348 VPWR.t3036 a_57692_11000# a_57604_11044# VPWR.t3035 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2349 a_33152_22091# a_32740_22504.t4 VGND.t93 VGND.t92 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2350 a_45372_14136# a_45284_14180# VGND.t2888 VGND.t2887 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2351 a_43646_21236# a_42982_21730# VGND.t5256 VGND.t5255 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2352 a_40436_26841# a_39124_27208.t3 a_40092_27209# VPWR.t220 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X2353 VGND.t6437 _402_.A1.t12 a_49172_27508# VGND.t6436 nfet_06v0 ad=0.3608p pd=2.52u as=0.1148p ps=1.1u w=0.82u l=0.6u
X2354 a_43890_24164# a_43750_23544# a_43126_24119# VGND.t4841 nfet_06v0 ad=43.2f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X2355 a_44296_24393.t3 clk.t3 VGND.t6525 VGND.t6524 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2356 VPWR.t3975 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN VPWR.t3974 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2357 a_45372_11000# a_45284_11044# VGND.t3218 VGND.t3217 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2358 a_51240_23340# _424_.B1.t10 VGND.t6334 VGND.t6333 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2359 a_53616_29480# _274_.A2 a_53412_29480# VPWR.t5896 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2360 VPWR.t4101 a_48060_12568# a_47972_12612# VPWR.t4100 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2361 a_64636_1159# a_64548_1256# VGND.t3951 VGND.t3950 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2362 a_43440_19325.t0 _452_.CLK.t40 VPWR.t6650 VPWR.t6649 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2363 a_56124_1159# a_56036_1256# VGND.t3953 VGND.t3952 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2364 a_62944_29101# _229_.I.t7 VGND.t6566 VGND.t6565 nfet_06v0 ad=57.59999f pd=0.68u as=0.218p ps=1.52u w=0.36u l=0.6u
X2365 VGND.t1451 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I VGND.t1450 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2366 a_43245_24373# hold1.Z hold2.I VGND.t3418 nfet_06v0 ad=92.99999f pd=1.015u as=0.2015p ps=1.295u w=0.775u l=0.6u
X2367 _457_.D _355_.C.t7 VGND.t6386 VGND.t6385 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X2368 VPWR.t5536 a_8636_1159# a_8548_1256# VPWR.t5535 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2369 VPWR.t3318 a_68108_12135# a_68020_12232# VPWR.t3317 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2370 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I VGND.t2172 VGND.t2171 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2371 VPWR.t6251 a_52988_1592# a_52900_1636# VPWR.t6250 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2372 a_66652_15704# a_66564_15748# VGND.t2934 VGND.t2933 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2373 VGND.t1511 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_56828_25940# VGND.t1009 nfet_06v0 ad=0.2132p pd=1.34u as=98.39999f ps=1.06u w=0.82u l=0.6u
X2374 VPWR.t3090 a_3708_21976# a_3620_22020# VPWR.t3089 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2375 VPWR.t6471 _459_.CLK.t27 a_29828_24455.t0 VPWR.t6470 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2376 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t5983 VGND.t5982 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2377 a_34400_25641# a_32180_25640.t4 a_34155_25273# VGND nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2378 a_58519_31220# a_58063_30644# VPWR.t3240 VPWR.t3239 pfet_06v0 ad=61.19999f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2379 a_20624_30345# a_18404_30344.t2 a_20379_29977# VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2380 a_45820_12568# a_45732_12612# VGND.t3826 VGND.t3044 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2381 a_3708_14136# a_3620_14180# VGND.t3827 VGND.t3542 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2382 a_49988_21236# _424_.A2.t8 _474_.D VGND.t185 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2383 a_54192_22851# a_53704_23219# a_54624_22895# VGND.t3829 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X2384 a_33052_15704# a_32964_15748# VGND.t3830 VGND.t3546 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2385 a_38764_20408# a_38676_20452# VGND.t3040 VGND.t3039 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2386 a_47271_21640# _421_.B a_47047_21640# VPWR.t3200 pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X2387 VGND.t3973 a_51048_26680# _284_.A2.t1 VGND.t3972 nfet_06v0 ad=0.23405p pd=1.555u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2388 VGND.t6234 _371_.A1.t14 _369_.ZN VGND.t6233 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2389 a_3708_11000# a_3620_11044# VGND.t3043 VGND.t2729 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2390 a_41116_26247# a_41028_26344# VGND.t3537 VGND.t3536 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2391 a_27564_20408# a_27476_20452# VGND.t3539 VGND.t3538 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2392 VPWR.t3688 a_17484_20408# a_17396_20452# VPWR.t3687 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2393 a_40092_27209# _442_.ZN a_39924_27209# VGND.t2807 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X2394 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t5661 VPWR.t5660 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2395 VPWR.t3690 a_65756_6296# a_65668_6340# VPWR.t3689 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2396 a_41488_24072# _304_.A1.t7 VPWR.t6603 VPWR.t6602 pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X2397 a_67660_12135# a_67572_12232# VGND.t4037 VGND.t4036 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2398 VPWR.t3300 _281_.A1 _384_.A3.t1 VPWR.t3299 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2399 _251_.ZN _251_.A1.t13 VGND.t6688 VGND.t6687 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X2400 VGND.t4963 _438_.A2 _431_.A3 VGND.t4962 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2401 VPWR.t4191 a_65756_3160# a_65668_3204# VPWR.t862 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2402 VPWR.t4235 a_65756_26247# a_65668_26344# VPWR.t4234 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2403 VGND.t3853 a_22352_25987# a_22304_26031# VGND.t3852 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X2404 a_56460_12135# a_56372_12232# VGND.t3855 VGND.t3854 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2405 VPWR.t5918 a_43804_30951# a_43716_31048# VPWR.t5917 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2406 _424_.A2.t1 _324_.B.t24 VPWR.t6710 VPWR.t6709 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2407 _301_.A1 a_35008_22461# VPWR.t6036 VPWR.t6035 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2408 VPWR.t6416 a_52064_19715.t4 a_52024_20083# VPWR.t6415 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2409 VPWR.t3496 a_65756_23111# a_65668_23208# VPWR.t3495 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2410 a_24876_23544# a_24788_23588# VGND.t3494 VGND.t3493 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2411 a_30796_24463# _459_.D a_30672_24831# VPWR.t3129 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X2412 VPWR.t3647 a_31484_26680# a_31396_26724# VPWR.t3646 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2413 a_42236_15271# a_42148_15368# VGND.t3498 VGND.t3497 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2414 a_48321_23208# _324_.B.t25 VPWR.t6712 VPWR.t6711 pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X2415 a_1916_4295# a_1828_4392# VGND.t3500 VGND.t3499 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2416 VGND.t6470 _359_.B.t7 _462_.D VGND.t102 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2417 a_65308_7864# a_65220_7908# VGND.t3310 VGND.t3309 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2418 VPWR.t3457 a_56124_27815# a_56036_27912# VPWR.t3456 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2419 a_36148_21976# _311_.A2.t7 VPWR.t6380 VPWR.t6379 pfet_06v0 ad=0.1391p pd=1.055u as=0.4268p ps=2.175u w=0.535u l=0.5u
X2420 _284_.ZN.t7 hold2.I VPWR.t2546 VPWR.t2545 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2421 VPWR.t3459 a_27564_21976# a_27476_22020# VPWR.t3458 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2422 a_41188_18840# _325_.A2.t6 VPWR.t6393 VPWR.t6392 pfet_06v0 ad=0.1391p pd=1.055u as=0.4268p ps=2.175u w=0.535u l=0.5u
X2423 a_65308_4728# a_65220_4772# VGND.t3097 VGND.t3096 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2424 a_66540_16839# a_66452_16936# VGND.t3099 VGND.t3098 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2425 VPWR.t3145 a_66876_15271# a_66788_15368# VPWR.t3144 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2426 VGND.t3251 _327_.A2 _328_.A2 VGND.t3250 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X2427 a_54816_22505# a_54040_22366# VGND.t3103 VGND.t3102 nfet_06v0 ad=43.2f pd=0.6u as=0.142p ps=1.14u w=0.36u l=0.6u
X2428 a_15244_25112# a_15156_25156# VGND.t661 VGND.t660 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2429 a_37291_29535# a_35728_29480# a_36656_29123# VGND.t663 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2430 a_23060_26724# _355_.C.t8 _454_.D VPWR.t6671 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2431 a_33724_1592# a_33636_1636# VGND.t667 VGND.t666 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2432 VGND.t2438 _349_.A4 a_25332_28776# VGND.t2437 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2433 VPWR.t2189 a_5388_16839# a_5300_16936# VPWR.t2188 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2434 a_15244_21976# a_15156_22020# VGND.t2344 VGND.t2343 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2435 VPWR.t2875 a_64412_19975# a_64324_20072# VPWR.t2874 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2436 VPWR.t2470 a_19500_20408# a_19412_20452# VPWR.t2469 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2437 VPWR.t1895 a_44476_15271# a_44388_15368# VPWR.t1894 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2438 VPWR.t2472 a_63292_12568# a_63204_12612# VPWR.t2471 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2439 a_4156_28248# a_4068_28292# VGND.t484 VGND.t483 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2440 a_40220_20408# a_40132_20452# VGND.t486 VGND.t485 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2441 VPWR.t489 a_52092_12568# a_52004_12612# VPWR.t488 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2442 VGND.t1217 a_52920_22760# _384_.A1 VGND.t1216 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2443 VPWR.t6177 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN VPWR.t2523 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2444 VPWR.t6283 a_51532_13703# a_51444_13800# VPWR.t6282 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2445 a_2364_18407# a_2276_18504# VGND.t490 VGND.t489 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2446 VPWR.t2516 a_45820_18840# a_45732_18884# VPWR.t2515 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2447 a_59226_25156# _251_.A1.t14 _251_.ZN VPWR.t7012 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2448 VPWR.t3314 a_11100_29816# a_11012_29860# VPWR.t3313 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2449 VPWR.t2266 a_29916_2727# a_29828_2824# VPWR.t2265 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2450 VPWR.t3657 a_45820_15704# a_45732_15748# VPWR.t3656 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2451 VPWR.t2518 a_63740_14136# a_63652_14180# VPWR.t2517 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2452 _335_.ZN.t15 _362_.B.t10 VPWR.t6532 VPWR.t6531 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2453 VPWR.t1580 a_67100_9432# a_67012_9476# VPWR.t1579 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2454 a_37532_26247# a_37444_26344# VGND.t494 VGND.t493 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2455 VPWR.t1373 a_66988_19975# a_66900_20072# VPWR.t1372 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2456 a_52408_19759# a_52064_19715.t5 a_51620_19911# VPWR.t6417 pfet_06v0 ad=0.1791p pd=1.355u as=0.1665p ps=1.285u w=0.36u l=0.5u
X2457 VPWR.t4327 _476_.Q _384_.A3.t5 VPWR.t4326 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2458 VPWR.t493 a_63740_11000# a_63652_11044# VPWR.t492 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2459 VPWR.t495 a_52540_14136# a_52452_14180# VPWR.t494 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2460 VPWR.t6652 _452_.CLK.t41 a_39124_27208.t0 VPWR.t6651 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2461 VPWR.t2474 a_52540_11000# a_52452_11044# VPWR.t2473 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2462 a_49852_15271# a_49764_15368# VGND.t2352 VGND.t2351 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2463 a_50120_26476# _411_.A2.t9 VGND.t111 VGND.t110 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2464 a_21600_26725# _346_.A2 _455_.D VPWR.t3636 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2465 VGND.t5748 _421_.A1 a_47291_25940# VGND.t5747 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2466 a_7292_29816# a_7204_29860# VGND.t2421 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2467 a_40196_31048# _296_.ZN VPWR.t3665 VPWR.t3664 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2468 _324_.C.t3 a_65072_29860# VPWR.t1112 VPWR.t1111 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2469 VPWR.t2550 a_20956_21543# a_20868_21640# VPWR.t2549 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2470 VPWR.t6273 a_49628_9432# a_49540_9476# VPWR.t6272 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2471 VPWR.t2552 a_59932_1159# a_59844_1256# VPWR.t2551 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2472 a_20396_20408# a_20308_20452# VGND.t2427 VGND.t2426 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2473 _284_.ZN.t18 _284_.B VPWR.t5595 VPWR.t5594 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2474 a_4156_18840# a_4068_18884# VGND.t1031 VGND.t1030 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2475 VPWR.t4149 a_39772_26247# a_39684_26344# VPWR.t4148 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2476 VPWR.t3587 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t3586 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2477 VPWR.t1174 a_31708_1592# a_31620_1636# VPWR.t1173 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2478 a_30812_18840# a_30724_18884# VGND.t1037 VGND.t1036 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2479 VPWR.t3108 a_17820_30951# a_17732_31048# VPWR.t3107 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2480 VPWR.t2689 a_26108_2727# a_26020_2824# VPWR.t2688 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2481 VPWR.t345 a_6620_1159# a_6532_1256# VPWR.t344 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2482 VPWR.t1 a_47948_23111# a_47860_23208# VPWR.t0 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2483 a_45372_10567# a_45284_10664# VGND.t340 VGND.t339 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2484 VPWR.t4637 a_58476_10567# a_58388_10664# VPWR.t4636 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2485 VPWR.t1400 a_62284_23544# a_62196_23588# VPWR.t1399 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2486 VPWR.t3668 a_33500_17272# a_33412_17316# VPWR.t417 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2487 VPWR.t3455 a_65308_7864# a_65220_7908# VPWR.t3454 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2488 a_40084_25156# _436_.ZN a_39860_25156# VPWR.t569 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2489 VPWR.t353 a_60156_27815# a_60068_27912# VPWR.t352 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2490 a_30476_25112# a_30388_25156# VGND.t346 VGND.t345 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2491 a_2364_1592# a_2276_1636# VGND.t348 VGND.t347 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2492 VPWR.t6257 a_25436_1592# a_25348_1636# VPWR.t6256 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2493 a_30364_1159# a_30276_1256# VGND.t1621 VGND.t1620 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2494 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I _241_.I0 VGND.t3741 VGND.t3740 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2495 a_19372_30345# _465_.D a_19248_29977# VPWR.t1177 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X2496 VPWR.t3494 a_49404_1592# a_49316_1636# VPWR.t2910 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2497 a_30476_21976# a_30388_22020# VGND.t1123 VGND.t1122 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2498 _250_.B _249_.A2 a_63952_29480# VPWR.t1532 pfet_06v0 ad=0.37665p pd=1.835u as=0.3402p ps=1.775u w=1.215u l=0.5u
X2499 a_45708_16839# a_45620_16936# VGND.t1125 VGND.t1124 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2500 VPWR.t1182 a_68108_20408# a_68020_20452# VPWR.t1181 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2501 _378_.I _379_.A2 VPWR.t2736 VPWR.t2735 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2502 VPWR.t4104 a_56124_1159# a_56036_1256# VPWR.t4103 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2503 VPWR.t3343 a_4828_2727# a_4740_2824# VPWR.t3342 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2504 a_22412_20408# a_22324_20452# VGND.t996 VGND.t995 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2505 a_3708_10567# a_3620_10664# VGND.t998 VGND.t997 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2506 a_7180_30951# a_7092_31048# VGND.t999 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2507 VPWR.t716 a_60604_26247# a_60516_26344# VPWR.t715 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2508 a_60828_2727# a_60740_2824# VGND.t4808 VGND.t1685 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2509 a_30924_23544# a_30836_23588# VGND.t4810 VGND.t4809 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2510 _424_.A2.t5 _324_.C.t16 a_45156_21236# VGND.t6506 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2511 a_47612_18407# a_47524_18504# VGND.t4812 VGND.t4811 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2512 a_36060_19369# _448_.D a_35892_19369# VGND.t637 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X2513 VPWR.t4410 a_64300_23544# a_64212_23588# VPWR.t4409 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2514 VPWR.t1273 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t1272 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2515 _355_.B _336_.A2.t5 a_28804_27208# VGND.t163 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2516 VGND.t4232 a_18760_29032# _379_.Z VGND.t4231 nfet_06v0 ad=0.218p pd=1.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2517 uo_out[6].t5 _287_.A1.t19 a_33028_27912# VPWR.t6783 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2518 a_1468_7431# a_1380_7528# VGND.t5856 VGND.t3062 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2519 a_42168_25640.t7 _304_.B _284_.ZN.t11 VGND.t4537 nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X2520 VPWR.t6980 _381_.A2.t3 a_49212_26369# VPWR.t6979 pfet_06v0 ad=0.4818p pd=3.07u as=0.4599p ps=1.935u w=1.095u l=0.5u
X2521 a_4156_30951# a_4068_31048# VGND.t5857 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2522 _244_.Z a_60212_25156# VPWR.t2730 VPWR.t2729 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2523 a_44296_24393.t4 clk.t4 VPWR.t6835 VPWR.t6834 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X2524 a_34448_25597# a_34155_25273# VPWR.t5915 VPWR.t5914 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X2525 a_41564_26247# a_41476_26344# VGND.t4937 VGND.t4936 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2526 a_3708_3160# a_3620_3204# VGND.t4939 VGND.t4938 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2527 VPWR.t5655 a_61724_15271# a_61636_15368# VPWR.t5654 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2528 VPWR.t2180 a_3260_16839# a_3172_16936# VPWR.t2179 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2529 VGND.t255 clkbuf_1_0__f_clk.I.t42 a_48272_25156.t11 VGND.t254 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2530 a_56516_26344# _251_.A1.t15 a_56368_26344# VPWR.t7013 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X2531 a_61940_29076# _229_.I.t8 _250_.C VGND.t6567 nfet_06v0 ad=0.2132p pd=1.34u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2532 a_57244_12568# a_57156_12612# VGND.t4908 VGND.t4907 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2533 VPWR.t6914 a_42392_22825.t19 _452_.CLK.t5 VPWR.t6913 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2534 VGND.t1664 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I VGND.t1663 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2535 a_24952_29032# _340_.A2 VPWR.t4880 VPWR.t4879 pfet_06v0 ad=0.156p pd=1.12u as=0.40575p ps=2.055u w=0.6u l=0.5u
X2536 _397_.A4 _470_.Q a_47173_27208# VGND.t4067 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2537 a_42684_15271# a_42596_15368# VGND.t4912 VGND.t4911 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2538 a_53436_19759# _424_.ZN a_52512_19715# VGND.t5734 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X2539 VPWR.t3243 a_47388_1592# a_47300_1636# VPWR.t3242 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2540 VGND.t118 a_49936_19325.t2 a_51308_19369# VGND.t117 nfet_06v0 ad=0.1584p pd=1.6u as=43.2f ps=0.6u w=0.36u l=0.6u
X2541 a_27908_27912# _371_.A3 VPWR.t980 VPWR.t979 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2542 VPWR.t6188 a_28348_21543# a_28260_21640# VPWR.t6187 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2543 a_22188_29383# a_22100_29480# VGND.t5929 VGND.t5928 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2544 VGND.t1324 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I VGND.t1323 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2545 a_4604_17272# a_4516_17316# VGND.t4827 VGND.t4826 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2546 VGND.t4973 vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I VGND.t4972 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2547 _323_.A3 _448_.Q.t5 a_38304_20072# VPWR.t6885 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X2548 a_15692_25112# a_15604_25156# VGND.t4829 VGND.t4828 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2549 a_55228_9432# a_55140_9476# VGND.t4831 VGND.t4830 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2550 a_4156_24679# a_4068_24776# VGND.t4833 VGND.t4832 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2551 a_67100_4295# a_67012_4392# VGND.t5877 VGND.t5658 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2552 a_15692_21976# a_15604_22020# VGND.t5878 VGND.t5062 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2553 VPWR.t3447 a_64860_19975# a_64772_20072# VPWR.t3446 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2554 a_61689_29860# _230_.I.t5 VPWR.t6632 VPWR.t6631 pfet_06v0 ad=0.1469p pd=1.085u as=0.38705p ps=2.08u w=0.565u l=0.5u
X2555 VPWR.t6394 _325_.A2.t7 a_43892_20072# VPWR.t4684 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2556 VPWR.t2153 _258_.ZN vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I VPWR.t2152 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2557 a_4156_21543# a_4068_21640# VGND.t5879 VGND.t3054 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2558 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I VPWR.t1955 VPWR.t1954 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2559 VPWR.t2802 a_24540_24679# a_24452_24776# VPWR.t2801 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2560 VPWR.t6967 _459_.Q.t6 a_29828_26344# VPWR.t6966 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X2561 VPWR.t2548 a_7292_29816# a_7204_29860# VPWR.t2547 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2562 VGND.t22 a_53744_22851.t2 a_53704_23219# VGND.t21 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2563 a_33148_25641# _460_.D a_33024_25273# VPWR.t6073 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X2564 a_55900_15271# a_55812_15368# VGND.t5892 VGND.t3066 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2565 VGND.t172 a_44784_25987.t3 a_46156_26031# VGND.t171 nfet_06v0 ad=0.1584p pd=1.6u as=43.2f ps=0.6u w=0.36u l=0.6u
X2566 VPWR.t6969 _459_.Q.t7 a_30724_26020# VPWR.t6968 pfet_06v0 ad=0.1391p pd=1.055u as=0.2354p ps=1.95u w=0.535u l=0.5u
X2567 VPWR.t2662 a_51980_13703# a_51892_13800# VPWR.t2661 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2568 vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN VPWR.t1121 VPWR.t1120 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2569 a_23284_26724# _345_.A2 a_23060_26724# VPWR.t3228 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2570 VPWR.t2256 a_43468_16839# a_43380_16936# VPWR.t2255 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2571 a_18472_29076# _379_.A2 VGND.t2597 VGND.t2596 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2572 a_40264_30320# _285_.Z VGND.t5707 VGND.t5706 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2573 a_57132_13703# a_57044_13800# VGND.t3075 VGND.t3074 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2574 VPWR.t4023 a_31260_19975# a_31172_20072# VPWR.t4022 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2575 uo_out[0].t6 _284_.ZN.t27 a_39300_31048# VPWR.t6516 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2576 a_23627_27967# a_22064_27912# a_22992_27555# VGND.t3267 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2577 a_34172_1159# a_34084_1256# VGND.t3284 VGND.t3283 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2578 a_33500_15271# a_33412_15368# VGND.t3286 VGND.t3285 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2579 VPWR.t5839 a_47612_9432# a_47524_9476# VPWR.t5838 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2580 a_36496_24463# a_35616_24776# a_36172_24463# VGND.t1587 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X2581 VPWR.t3429 a_3708_27815# a_3620_27912# VPWR.t3428 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2582 VGND.t1556 vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I VGND.t1555 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2583 VGND.t4906 _250_.C _250_.ZN VGND.t4905 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X2584 a_41572_18504# _332_.Z VPWR.t5044 VPWR.t5043 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2585 VPWR.t3169 a_50188_12135# a_50100_12232# VPWR.t3168 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2586 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I VGND.t1523 VGND.t1522 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2587 a_37980_26247# a_37892_26344# VGND.t3014 VGND.t3013 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2588 VPWR.t3175 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN VPWR.t3174 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2589 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t1246 VGND.t1245 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2590 VPWR.t1898 a_1468_10567# a_1380_10664# VPWR.t1897 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2591 a_47836_17272# a_47748_17316# VGND.t2910 VGND.t2909 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2592 VPWR.t6095 a_23420_26247# a_23332_26344# VPWR.t6094 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2593 VPWR.t2591 a_16916_31048# a_16916_31048# VPWR.t2590 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2594 a_49404_30951# a_49316_31048# VGND.t2911 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2595 VPWR.t3069 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I VPWR.t3068 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2596 VPWR.t7051 ui_in[0].t0 a_63616_31128# VPWR.t7050 pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X2597 VPWR.t3538 a_53324_10567# a_53236_10664# VPWR.t3537 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2598 VPWR.t3625 a_53548_18407# a_53460_18504# VPWR.t3624 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2599 a_58588_21543# a_58500_21640# VGND.t3944 VGND.t3943 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2600 a_27116_23544# a_27028_23588# VGND.t3946 VGND.t3945 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2601 a_28124_1592# a_28036_1636# VGND.t3948 VGND.t3947 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2602 VPWR.t4306 a_46940_15271# a_46852_15368# VPWR.t4305 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2603 a_36500_29860# _288_.ZN.t5 VPWR.t6330 VPWR.t6329 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X2604 a_36636_17272# a_36548_17316# VGND.t592 VGND.t591 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2605 VPWR.t6023 a_23420_1592# a_23332_1636# VPWR.t6022 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2606 VPWR.t2448 _393_.A3 a_46804_28292# VPWR.t2447 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2607 VPWR.t4884 a_1020_8999# a_932_9096# VPWR.t4883 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2608 VPWR.t2370 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN VPWR.t2369 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2609 a_55340_26680# a_55252_26724# VGND.t594 VGND.t593 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2610 a_33728_29167# a_31508_29159.t6 a_33483_29535# VGND.t89 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2611 a_40565_24394# _435_.ZN VGND.t4681 VGND.t4680 nfet_06v0 ad=85.2f pd=0.95u as=0.3124p ps=2.3u w=0.71u l=0.6u
X2612 VPWR.t3115 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I VPWR.t3114 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2613 a_27004_30951# a_26916_31048# VGND.t761 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2614 VPWR.t1584 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I a_60416_25156# VPWR.t1583 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X2615 VPWR.t1369 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I VPWR.t1368 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2616 vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I VPWR.t2831 VPWR.t2830 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2617 _474_.CLK.t12 a_48272_25156.t26 VGND.t6270 VGND.t6269 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2618 VPWR.t781 a_2812_5863# a_2724_5960# VPWR.t780 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2619 a_32352_29535# a_31920_29480# VPWR.t3292 VPWR.t3291 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X2620 VGND.t4031 a_41160_29083# uo_out[3].t6 VGND.t4030 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X2621 VPWR.t1297 a_2812_2727# a_2724_2824# VPWR.t1296 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2622 VPWR.t783 a_63404_12135# a_63316_12232# VPWR.t782 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2623 a_53436_18840# a_53348_18884# VGND.t4274 VGND.t4273 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2624 a_51877_21236# _281_.A1 _281_.ZN.t1 VGND.t3147 nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2625 VGND.t5503 a_37360_19325# a_37312_19369# VGND.t5502 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X2626 VPWR.t6014 a_49852_2727# a_49764_2824# VPWR.t6013 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2627 VPWR.t4432 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I VPWR.t4431 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2628 VGND.t5514 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2629 VPWR.t5897 a_42908_1159# a_42820_1256# VPWR.t5308 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2630 VPWR.t3563 a_29916_1592# a_29828_1636# VPWR.t1823 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2631 a_6844_1592# a_6756_1636# VGND.t423 VGND.t422 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2632 VPWR.t1110 a_65072_29860# _324_.C.t2 VPWR.t1109 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2633 a_45128_26031# a_44744_26355# a_44340_26183# VGND.t6031 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2634 VPWR.t2728 a_60212_25156# _244_.Z VPWR.t2727 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X2635 VPWR.t6028 a_3708_18407# a_3620_18504# VPWR.t5798 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2636 VPWR.t5066 a_51868_9432# a_51780_9476# VPWR.t5065 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2637 VPWR.t5680 a_14796_26247# a_14708_26344# VPWR.t1936 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2638 a_30160_30301# a_29788_30345# VPWR.t1933 VPWR.t1932 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X2639 VPWR.t2679 a_26668_23544# a_26580_23588# VPWR.t2678 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2640 VGND.t1029 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN _245_.I1 VGND.t1028 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2641 VPWR.t6749 _474_.CLK.t38 _276_.A2 VPWR.t6748 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2642 VPWR.t5234 a_36636_1159# a_36548_1256# VPWR.t5233 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2643 a_3260_12568# a_3172_12612# VGND.t4900 VGND.t4899 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2644 VPWR.t5984 a_14796_23111# a_14708_23208# VPWR.t1972 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2645 VPWR.t5988 a_17932_24679# a_17844_24776# VPWR.t2127 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2646 VPWR.t943 a_52512_19715# a_52408_19759# VPWR.t942 pfet_06v0 ad=0.1044p pd=0.94u as=0.1791p ps=1.355u w=0.36u l=0.5u
X2647 a_39748_29480# _284_.ZN.t28 uo_out[1].t6 VPWR.t6517 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2648 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN VPWR.t2862 VPWR.t2861 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2649 VPWR.t2697 a_52316_2727# a_52228_2824# VPWR.t2696 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2650 a_22860_20408# a_22772_20452# VGND.t4902 VGND.t4901 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2651 a_60492_28248# a_60404_28292# VGND.t4904 VGND.t4903 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2652 a_27004_2727# a_26916_2824# VGND.t4803 VGND.t4802 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2653 a_56348_1592# a_56260_1636# VGND.t4805 VGND.t4804 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2654 a_22964_27967# a_21652_27591.t5 a_22620_27599# VPWR.t104 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X2655 VPWR.t3877 a_51644_1592# a_51556_1636# VPWR.t3876 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2656 VPWR.t2681 _383_.ZN a_48141_29480# VPWR.t2680 pfet_06v0 ad=0.5346p pd=3.31u as=0.37665p ps=1.835u w=1.215u l=0.5u
X2657 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I VGND.t1449 VGND.t1448 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2658 a_27004_21543# a_26916_21640# VGND.t4807 VGND.t4806 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2659 VPWR.t3402 _327_.A2 a_44276_20072# VPWR.t3401 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X2660 VPWR.t640 a_46044_2727# a_45956_2824# VPWR.t639 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2661 VPWR.t4308 a_59372_13703# a_59284_13800# VPWR.t4307 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2662 VPWR.t4967 a_63180_26680# a_63092_26724# VPWR.t4966 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2663 a_3708_29816# a_3620_29860# VGND.t4821 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2664 a_61164_13703# a_61076_13800# VGND.t4823 VGND.t4822 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2665 a_64748_23544# a_64660_23588# VGND.t4825 VGND.t4824 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2666 _332_.Z a_40244_18180# VGND.t878 VGND.t877 nfet_06v0 ad=0.341p pd=2.43u as=0.2424p ps=1.635u w=0.775u l=0.6u
X2667 VPWR.t2030 _287_.A2 a_33476_27912# VPWR.t2029 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2668 VPWR.t6308 a_49740_10567# a_49652_10664# VPWR.t6307 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2669 VPWR.t5088 a_59260_21976# a_59172_22020# VPWR.t5087 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2670 VPWR.t5090 a_25008_25597# a_24980_25273# VPWR.t5089 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X2671 a_18400_28733# a_18028_28777# VPWR.t2641 VPWR.t2640 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X2672 a_1468_19975# a_1380_20072# VGND.t4935 VGND.t2711 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2673 a_37324_28776# _334_.A1 _335_.ZN.t6 VGND.t2244 nfet_06v0 ad=0.1312p pd=1.14u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2674 VPWR.t4129 a_46716_10567# a_46628_10664# VPWR.t1419 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2675 a_36764_22512# _304_.A1.t8 a_36560_22512# VGND.t6318 nfet_06v0 ad=60.8f pd=0.7u as=79.8f ps=0.8u w=0.38u l=0.6u
X2676 a_51868_17272# a_51780_17316# VGND.t5848 VGND.t5847 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2677 a_59620_27208# _245_.Z VGND.t5828 VGND.t5827 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2678 _439_.ZN _438_.ZN VGND.t2513 VGND.t2512 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2679 a_57692_12568# a_57604_12612# VGND.t5852 VGND.t5851 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2680 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I VPWR.t2745 VPWR.t2744 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2681 a_5724_2727# a_5636_2824# VGND.t5854 VGND.t5853 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2682 VPWR.t6113 a_64412_6296# a_64324_6340# VPWR.t5306 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2683 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t5807 VGND.t5231 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2684 VPWR.t6916 a_42392_22825.t20 _452_.CLK.t6 VPWR.t6915 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2685 VGND.t6483 _287_.A1.t20 uo_out[5].t7 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2686 VPWR.t1750 a_36016_20893# a_36008_20569# VPWR.t1749 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X2687 VPWR.t4551 _330_.A2 a_38842_17316# VPWR.t4550 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X2688 VPWR.t6148 a_64412_3160# a_64324_3204# VPWR.t6147 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2689 a_37532_26680# a_37444_26724# VGND.t5887 VGND.t5886 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2690 VPWR.t6151 a_59820_12135# a_59732_12232# VPWR.t6150 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2691 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN VPWR.t2209 VPWR.t2208 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2692 a_48060_14136# a_47972_14180# VGND.t3876 VGND.t3875 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2693 a_22352_25987# a_22059_26399# VGND.t5616 VGND.t5615 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X2694 VGND.t4120 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN a_63721_28776# VGND.t4119 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2695 VPWR.t3415 a_50076_15704# a_49988_15748# VPWR.t3414 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2696 VPWR.t5906 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I VPWR.t3736 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2697 VPWR.t6837 clk.t5 a_44296_24393.t5 VPWR.t6836 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X2698 VGND.t6735 ui_in[4].t0 a_58063_30644# VGND.t45 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X2699 VPWR.t2047 a_37584_29123# a_37576_29535# VPWR.t2046 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X2700 VPWR.t4035 a_28796_21543# a_28708_21640# VPWR.t4034 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2701 VPWR.t3372 a_44864_27165# a_44856_26841# VPWR.t3371 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X2702 a_48060_11000# a_47972_11044# VGND.t5039 VGND.t5038 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2703 a_48272_25156.t10 clkbuf_1_0__f_clk.I.t43 VGND.t257 VGND.t256 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2704 a_3708_23544# a_3620_23588# VGND.t5040 VGND.t4407 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2705 _393_.A3 _324_.C.t17 a_50197_28776# VGND.t6507 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2706 a_55228_2727# a_55140_2824# VGND.t5041 VGND.t2753 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2707 VPWR.t5200 a_58588_1159# a_58500_1256# VPWR.t456 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2708 a_55116_22895# _478_.D a_54192_22851# VGND.t5813 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X2709 VPWR.t5390 a_3260_18840# a_3172_18884# VPWR.t1813 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2710 a_49448_20072# _417_.A2.t5 _417_.Z VPWR.t131 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2711 VPWR.t3860 a_62620_18407# a_62532_18504# VPWR.t3859 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2712 VPWR.t2372 a_5276_1159# a_5188_1256# VPWR.t2371 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2713 _419_.A4 _412_.A1 VGND.t3691 VGND.t3690 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X2714 VPWR.t4588 a_3260_15704# a_3172_15748# VPWR.t873 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2715 a_52452_24072# _424_.A2.t9 VPWR.t190 VPWR.t189 pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X2716 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN VGND.t4460 VGND.t4459 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2717 VPWR.t5396 a_20396_27815# a_20308_27912# VPWR.t5395 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2718 _301_.Z a_38340_21327# VPWR.t5147 VPWR.t5146 pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X2719 VPWR.t6654 _452_.CLK.t42 a_42596_27208.t0 VPWR.t6653 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2720 VGND.t5599 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN _267_.A1 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2721 a_65756_7864# a_65668_7908# VGND.t5601 VGND.t5020 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2722 _452_.CLK.t7 a_42392_22825.t21 VGND.t6603 VGND.t6602 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2723 a_57580_13703# a_57492_13800# VGND.t5603 VGND.t5602 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2724 VGND.t3122 hold2.Z a_42587_25940# VGND.t3121 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2725 _386_.ZN _404_.A1 VGND.t3675 VGND.t3674 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2726 VPWR.t3663 _296_.ZN a_39748_31048# VPWR.t3662 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2727 a_65756_4728# a_65668_4772# VGND.t967 VGND.t966 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2728 a_67324_15271# a_67236_15368# VGND.t969 VGND.t968 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2729 a_31036_21543# a_30948_21640# VGND.t971 VGND.t970 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2730 VPWR.t1004 a_19612_21543# a_19524_21640# VPWR.t1003 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2731 a_19052_20408# a_18964_20452# VGND.t975 VGND.t974 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2732 a_46984_23588# _397_.A1.t7 VGND.t11 VGND.t10 nfet_06v0 ad=0.126p pd=1.06u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2733 a_46352_22021# _421_.A1 _402_.ZN VPWR.t5997 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2734 VPWR.t3050 a_64972_10567# a_64884_10664# VPWR.t3049 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2735 VPWR.t1334 a_5388_26247# a_5300_26344# VPWR.t1333 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2736 a_49852_30951# a_49764_31048# VGND.t1096 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2737 a_10428_29383# a_10340_29480# VGND.t1098 VGND.t1097 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2738 a_24304_26795# a_23892_27208.t3 VPWR.t6339 VPWR.t6338 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2739 a_25962_29480# _349_.A4 _340_.ZN VPWR.t2559 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2740 VPWR.t2018 a_53772_10567# a_53684_10664# VPWR.t2017 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2741 a_27564_23544# a_27476_23588# VGND.t1103 VGND.t1102 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2742 a_66092_18407# a_66004_18504# VGND.t3918 VGND.t3917 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2743 VPWR.t2020 a_53996_18407# a_53908_18504# VPWR.t2019 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2744 VPWR.t4799 _474_.Q a_48964_20204# VPWR.t4798 pfet_06v0 ad=0.4005p pd=2.12u as=0.1456p ps=1.08u w=0.56u l=0.5u
X2745 VPWR.t4703 a_5388_23111# a_5300_23208# VPWR.t4702 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2746 VGND.t5883 a_63616_31128# _251_.A1.t6 VGND.t5880 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X2747 VGND.t1602 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t1601 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2748 VPWR.t3962 _427_.B1 a_53076_24776# VPWR.t3961 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2749 _250_.A2 _248_.B1 a_63313_28776# VGND.t1147 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2750 a_42896_18504# a_42484_18183.t2 VPWR.t7045 VPWR.t7044 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2751 a_63068_18407# a_62980_18504# VGND.t3920 VGND.t3919 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2752 VPWR.t4139 a_46492_15704# a_46404_15748# VPWR.t66 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2753 a_29788_30345# _370_.ZN a_29620_30345# VGND.t137 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X2754 VPWR.t2315 a_34620_1159# a_34532_1256# VPWR.t2314 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2755 vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t6058 VPWR.t6057 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2756 VPWR.t2316 a_2812_21543# a_2724_21640# VPWR.t1298 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2757 VPWR.t1756 a_21516_23544# a_21428_23588# VPWR.t1755 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2758 a_16252_30951# a_16164_31048# VGND.t2210 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2759 a_63292_14136# a_63204_14180# VGND.t2212 VGND.t2211 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2760 VPWR.t2322 a_63404_20408# a_63316_20452# VPWR.t2321 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2761 VGND.t3227 a_44864_27165# a_44816_27209# VGND.t3226 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X2762 VPWR.t5377 a_35292_15704# a_35204_15748# VPWR.t5376 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2763 _450_.D _330_.A1.t12 a_41776_20072# VPWR.t214 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2764 VGND.t6690 _251_.A1.t16 a_55956_25940# VGND.t6689 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2765 VPWR.t4968 a_3708_29816# a_3620_29860# VPWR.t4285 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2766 VPWR.t3854 a_63852_12135# a_63764_12232# VPWR.t3853 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2767 VPWR.t3800 a_34732_16839# a_34644_16936# VPWR.t3799 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2768 a_63292_11000# a_63204_11044# VGND.t3715 VGND.t3714 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2769 a_30364_1592# a_30276_1636# VGND.t3716 VGND.t3177 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2770 a_52092_14136# a_52004_14180# VGND.t3452 VGND.t3181 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2771 a_17140_26841# a_15828_27208.t3 a_16796_27209# VPWR.t6382 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X2772 a_60268_14136# a_60180_14180# VGND.t3454 VGND.t3453 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2773 a_49448_20072# a_48776_20204# VPWR.t3611 VPWR.t3610 pfet_06v0 ad=0.3172p pd=1.74u as=0.4005p ps=2.12u w=1.22u l=0.5u
X2774 VPWR.t4991 _302_.Z _324_.B.t14 VPWR.t4990 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2775 _422_.ZN _476_.Q a_52997_20936# VGND.t4163 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2776 VPWR.t3612 a_3708_26680# a_3620_26724# VPWR.t70 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2777 a_54332_1592# a_54244_1636# VGND.t3459 VGND.t3458 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2778 a_52092_11000# a_52004_11044# VGND.t2190 VGND.t2189 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2779 VPWR.t3700 a_20060_2727# a_19972_2824# VPWR.t3699 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2780 VPWR.t2757 a_65420_13703# a_65332_13800# VPWR.t2756 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2781 VPWR.t1935 a_31708_16839# a_31620_16936# VPWR.t1934 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2782 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I VPWR.t3973 VPWR.t3972 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2783 VPWR.t1931 a_2364_13703# a_2276_13800# VPWR.t693 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2784 VGND.t3210 input9.Z _268_.A1.t1 VGND.t3209 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2785 a_37968_31048# _285_.Z VPWR.t5932 VPWR.t5931 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2786 a_25340_29167# _340_.A2 VGND.t4732 VGND.t4731 nfet_06v0 ad=58.39999f pd=0.685u as=0.23405p ps=1.555u w=0.365u l=0.6u
X2787 VGND.t3378 a_33776_29123# _362_.B.t2 VGND.t3377 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2788 VGND.t6388 _355_.C.t9 _351_.ZN VGND.t6387 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X2789 a_1020_1592# a_932_1636# VGND.t2968 VGND.t2922 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2790 VPWR.t3247 a_54220_13703# a_54132_13800# VPWR.t3246 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2791 VPWR.t2059 a_34080_22461# a_34052_22137# VPWR.t2058 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X2792 _427_.A2 _417_.A2.t6 a_51332_24072# VGND.t130 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2793 a_51436_27208# _384_.A3.t12 VGND.t178 VGND.t177 nfet_06v0 ad=58.39999f pd=0.685u as=0.23405p ps=1.555u w=0.365u l=0.6u
X2794 VPWR.t5128 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN VPWR.t5127 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2795 VPWR.t4245 a_3708_7431# a_3620_7528# VPWR.t4244 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2796 a_48060_1592# a_47972_1636# VGND.t2970 VGND.t2969 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2797 a_43850_23588# a_43750_23544# a_43126_24119# VPWR.t4983 pfet_06v0 ad=61.19999f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2798 _351_.A2 _346_.A2 a_24900_27912# VPWR.t3635 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2799 VPWR.t2006 a_32828_2727# a_32740_2824# VPWR.t2005 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2800 VGND.t6692 _251_.A1.t17 _250_.B VGND.t6691 nfet_06v0 ad=0.22595p pd=1.45u as=0.21175p ps=1.41u w=0.465u l=0.6u
X2801 a_44856_26841# a_43008_26795# a_44571_26841# VPWR.t6008 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X2802 a_37576_29535# a_35728_29480# a_37291_29535# VPWR.t670 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X2803 a_62172_15704# a_62084_15748# VGND.t3663 VGND.t3662 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2804 a_42630_21236# a_42154_21236# VGND.t2381 VGND.t2380 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2805 a_63740_12568# a_63652_12612# VGND.t3665 VGND.t3664 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2806 VGND.t3789 a_35816_21192# _319_.A3 VGND.t3788 nfet_06v0 ad=0.23405p pd=1.555u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2807 a_52540_12568# a_52452_12612# VGND.t3667 VGND.t3666 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2808 VPWR.t6223 a_26556_2727# a_26468_2824# VPWR.t6222 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2809 VPWR.t3040 a_2812_4728# a_2724_4772# VPWR.t3039 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2810 a_62060_23111# a_61972_23208# VGND.t2891 VGND.t2890 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2811 a_27452_21543# a_27364_21640# VGND.t2893 VGND.t2892 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2812 VPWR.t5820 a_65756_7864# a_65668_7908# VPWR.t5819 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2813 VPWR.t2456 _264_.B a_42161_24776# VPWR.t2455 pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2814 a_25232_27165# a_24860_27209# VPWR.t5358 VPWR.t5357 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X2815 VGND.t610 a_23920_27555# a_23872_27599# VGND.t609 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X2816 VPWR.t3048 a_2812_12135# a_2724_12232# VPWR.t3047 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2817 _397_.Z a_46984_23588# VGND.t832 VGND.t831 nfet_06v0 ad=0.3608p pd=2.52u as=0.218p ps=1.52u w=0.82u l=0.6u
X2818 VPWR.t3707 a_2812_1592# a_2724_1636# VPWR.t76 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2819 VPWR.t5472 a_25884_1592# a_25796_1636# VPWR.t5471 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2820 a_43003_28409# a_41440_28363# a_42368_28733# VGND.t1454 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2821 a_18048_27209# a_15828_27208.t4 a_17803_26841# VGND.t6112 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2822 VPWR.t4176 a_62844_1159# a_62756_1256# VPWR.t4175 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2823 VPWR.t4147 a_49852_1592# a_49764_1636# VPWR.t4146 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2824 VPWR.t4178 a_14796_28248# a_14708_28292# VPWR.t4177 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2825 VPWR.t4180 a_23644_21543# a_23556_21640# VPWR.t4179 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2826 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I VGND.t6787 VGND.t6786 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2827 _245_.I1 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t1027 VGND.t1026 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2828 _403_.ZN _324_.C.t18 VPWR.t6799 VPWR pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2829 VGND.t3591 a_42796_23981# hold2.Z VGND.t3590 nfet_06v0 ad=0.28262p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2830 a_36544_24419# a_36172_24463# VGND.t5446 VGND.t5445 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X2831 VPWR.t5243 a_3708_17272# a_3620_17316# VPWR.t5242 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2832 a_39332_23588# _434_.ZN VPWR.t1289 VPWR.t1288 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2833 VPWR.t3601 a_14796_25112# a_14708_25156# VPWR.t3600 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2834 a_33500_18840# a_33412_18884# VGND.t3593 VGND.t3592 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2835 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I VGND.t6048 VGND.t6047 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2836 VGND.t922 a_52512_19715# a_52408_19759# VGND.t921 nfet_06v0 ad=0.2637p pd=1.825u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2837 a_53212_2727# a_53124_2824# VGND.t3599 VGND.t3598 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2838 VPWR.t6051 a_46268_9432# a_46180_9476# VPWR.t6050 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2839 VPWR.t4166 a_56572_1159# a_56484_1256# VPWR.t4165 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2840 a_33472_25641# a_32592_25227# a_33148_25641# VGND.t5691 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X2841 VPWR.t4168 a_3260_4295# a_3172_4392# VPWR.t4167 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2842 a_48060_10567# a_47972_10664# VGND.t4015 VGND.t2333 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2843 VPWR.t4174 a_44752_18147# a_44744_18559# VPWR.t4173 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X2844 VPWR.t2492 a_17932_23544# a_17844_23588# VPWR.t2491 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2845 VPWR.t5816 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN _267_.A1 VPWR.t5815 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2846 VPWR.t2280 a_3260_1159# a_3172_1256# VPWR.t2279 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2847 a_1020_26247# a_932_26344# VGND.t2176 VGND.t2175 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2848 a_30795_29977# a_28820_30344.t4 a_30160_30301# VPWR.t6366 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X2849 a_53300_23047# a_53744_22851.t3 a_53696_22895# VGND.t23 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X2850 a_31484_30951# a_31396_31048# VGND.t2180 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2851 VGND.t2779 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I VGND.t2778 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2852 VGND.t2046 _258_.ZN vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I VGND.t2045 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X2853 VPWR.t6851 _455_.Q.t6 _371_.A2 VPWR.t6850 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2854 a_41440_28363# a_41028_28776.t2 VPWR.t7097 VPWR.t7096 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2855 VPWR.t2232 a_17036_26247# a_16948_26344# VPWR.t2231 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2856 VGND.t6439 _402_.A1.t13 _383_.A2 VGND.t6438 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2857 VPWR.t2820 a_23084_21976# a_22996_22020# VPWR.t2819 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2858 a_1020_23111# a_932_23208# VGND.t2682 VGND.t2681 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2859 VPWR.t1870 a_22076_1592# a_21988_1636# VPWR.t1869 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2860 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN _248_.B1 VGND.t1146 VGND.t1145 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2861 a_2812_27815# a_2724_27912# VGND.t2684 VGND.t2683 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2862 _324_.C.t6 a_65072_29860# VGND.t1062 VGND.t1059 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X2863 VPWR.t3356 input9.Z _268_.A1.t0 VPWR.t3355 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2864 VPWR.t2836 a_17036_23111# a_16948_23208# VPWR.t415 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2865 VPWR.t5473 a_46044_1592# a_45956_1636# VPWR.t2235 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2866 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].I VPWR.t5202 VPWR.t1424 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2867 VPWR.t3483 _460_.Q _371_.A1.t5 VPWR.t3482 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2868 VPWR.t4635 a_51196_15271# a_51108_15368# VPWR.t4634 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2869 VPWR.t3741 a_26220_20408# a_26132_20452# VPWR.t3740 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2870 VPWR.t3743 a_3260_29383# a_3172_29480# VPWR.t3742 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2871 VGND.t5737 a_21424_25987# a_21376_26031# VGND.t5736 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X2872 VPWR.t4513 a_56348_12568# a_56260_12612# VPWR.t4512 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2873 VPWR.t3745 a_1468_5863# a_1380_5960# VPWR.t3744 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2874 a_25100_20408# a_25012_20452# VGND.t3605 VGND.t3604 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2875 VPWR.t2713 a_47612_13703# a_47524_13800# VPWR.t1044 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2876 VPWR.t2186 a_3260_26247# a_3172_26344# VPWR.t2185 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2877 a_29468_2727# a_29380_2824# VGND.t3127 VGND.t3126 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2878 VPWR.t530 a_1468_2727# a_1380_2824# VPWR.t529 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2879 a_51988_24776# _412_.A1 _412_.ZN VPWR.t3840 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2880 VPWR.t2741 a_3260_23111# a_3172_23208# VPWR.t421 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2881 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I VPWR.t3280 VPWR.t3279 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2882 clkload0.Z a_48384_26724# VPWR.t3006 VPWR.t3005 pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X2883 a_19035_28409# a_17060_28776.t5 a_18400_28733# VPWR.t6907 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X2884 a_44700_30951# a_44612_31048# VGND.t3132 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2885 a_13788_29816# a_13700_29860# VGND.t3133 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2886 a_41828_28777# a_41028_28776.t3 VGND.t6776 VGND.t6775 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2887 a_29736_27508# _350_.A2.t24 VGND.t6294 VGND.t6293 nfet_06v0 ad=98.39999f pd=1.06u as=0.2405p ps=1.52u w=0.82u l=0.6u
X2888 VPWR.t3788 a_59820_14136# a_59732_14180# VPWR.t3787 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2889 VPWR.t6656 _452_.CLK.t43 a_36996_18183.t0 VPWR.t6655 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2890 VPWR.t5097 a_55788_24679# a_55700_24776# VPWR.t4537 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2891 VPWR.t4873 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I VPWR.t4872 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2892 a_61948_9432# a_61860_9476# VGND.t3647 VGND.t3646 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2893 a_57132_17272# a_57044_17316# VGND.t3649 VGND.t3648 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2894 a_50732_23233# _395_.A2 a_50420_23233# VPWR.t5848 pfet_06v0 ad=0.2847p pd=1.615u as=0.58035p ps=2.155u w=1.095u l=0.5u
X2895 a_65308_17272# a_65220_17316# VGND.t3968 VGND.t3967 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2896 a_34080_22461# a_33708_22505# VGND.t3576 VGND.t3575 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X2897 VGND.t3969 a_12548_31048# uio_oe[3].t0 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2898 _350_.A2.t6 _337_.ZN a_30388_28776# VGND.t4979 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2899 a_42392_22825.t4 clkbuf_1_0__f_clk.I.t44 VPWR.t254 VPWR.t253 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X2900 VPWR.t3883 _241_.I0 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I VPWR.t3882 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X2901 VPWR.t1872 a_64412_15271# a_64324_15368# VPWR.t1871 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2902 VPWR.t4319 a_41340_15704# a_41252_15748# VPWR.t4318 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2903 a_51317_27508# _397_.A4 VGND.t1252 VGND.t1251 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2904 a_1020_16839# a_932_16936# VGND.t3971 VGND.t3970 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2905 a_67772_15271# a_67684_15368# VGND.t3922 VGND.t3921 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2906 a_25936_25597# a_25643_25273# VPWR.t4072 VPWR.t4071 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X2907 a_31484_21543# a_31396_21640# VGND.t3926 VGND.t3925 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2908 _270_.A2 a_58911_30644# VGND.t2788 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.28262p ps=1.87u w=0.82u l=0.6u
X2909 a_55676_9432# a_55588_9476# VGND.t3928 VGND.t3927 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2910 VPWR.t4080 a_53996_26680# a_53908_26724# VPWR.t4079 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2911 a_10876_29383# a_10788_29480# VGND.t3932 VGND.t3931 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2912 _371_.A2 _337_.A3.t8 a_27868_28776# VGND.t6140 nfet_06v0 ad=0.4161p pd=1.905u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2913 VPWR.t2759 a_9084_30951# a_8996_31048# VPWR.t2758 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2914 VPWR.t5971 a_52415_31220# a_52871_31198# VPWR.t5970 pfet_06v0 ad=0.379p pd=2.37u as=61.19999f ps=0.7u w=0.36u l=0.5u
X2915 a_2364_9432# a_2276_9476# VGND.t3846 VGND.t3845 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2916 a_45372_15271# a_45284_15368# VGND.t3847 VGND.t2887 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2917 a_53716_26399# _412_.ZN a_52848_25987# VPWR.t5256 pfet_06v0 ad=54f pd=0.66u as=0.1872p ps=1.4u w=0.36u l=0.5u
X2918 VPWR.t2761 a_35740_30951# a_35652_31048# VPWR.t2760 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2919 VPWR.t5938 a_62620_17272# a_62532_17316# VPWR.t5937 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2920 VGND.t5329 a_58687_31220# a_59163_30644# VGND.t45 nfet_06v0 ad=0.28262p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2921 VGND.t5882 a_63616_31128# _251_.A1.t5 VGND.t5880 nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X2922 a_34939_23705# a_33376_23659# a_34304_24029# VGND.t1813 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2923 _247_.ZN _243_.ZN a_59172_27912# VPWR.t4042 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2924 a_2364_6296# a_2276_6340# VGND.t3756 VGND.t3755 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2925 a_45372_12135# a_45284_12232# VGND.t3757 VGND.t3217 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2926 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I VPWR.t3991 VPWR.t3990 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2927 VPWR.t6473 _459_.CLK.t28 a_20084_26023.t0 VPWR.t6472 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2928 VPWR.t6018 a_51420_17272# a_51332_17316# VPWR.t6017 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2929 VPWR.t3358 a_35292_26247# a_35204_26344# VPWR.t3357 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2930 _250_.C _229_.I.t9 a_62148_29505# VPWR.t6873 pfet_06v0 ad=0.31207p pd=1.665u as=0.55297p ps=2.105u w=1.095u l=0.5u
X2931 a_18380_25112# a_18292_25156# VGND.t2653 VGND.t2652 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2932 VPWR.t2796 a_20396_26680# a_20308_26724# VPWR.t2795 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2933 VPWR.t2532 a_21964_23544# a_21876_23588# VPWR.t2531 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2934 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I VGND.t5517 VGND.t2171 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2935 a_60268_10567# a_60180_10664# VGND.t2657 VGND.t2656 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2936 VPWR.t2334 a_30812_2727# a_30724_2824# VPWR.t2333 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2937 VPWR.t2358 _334_.A1 _371_.A1.t1 VPWR.t2357 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2938 a_26548_24372# _336_.A2.t6 _352_.ZN VGND.t164 nfet_06v0 ad=0.2132p pd=1.34u as=0.4161p ps=1.905u w=0.82u l=0.6u
X2939 a_8636_29383# a_8548_29480# VGND.t2659 VGND.t2658 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2940 a_18380_21976# a_18292_22020# VGND.t2258 VGND.t2257 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2941 a_50280_19369# a_49936_19325.t3 a_49492_18840# VPWR.t121 pfet_06v0 ad=0.1791p pd=1.355u as=0.1665p ps=1.285u w=0.36u l=0.5u
X2942 VGND.t2521 _274_.A1 a_52756_29076# VGND.t2520 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2943 VGND.t6517 _325_.A1.t11 _226_.ZN VGND.t6516 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2944 VPWR.t1852 a_24092_23111# a_24004_23208# VPWR.t1851 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2945 a_25792_30301# a_25420_30345# VPWR.t5232 VPWR.t5231 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X2946 a_63628_16839# a_63540_16936# VGND.t2264 VGND.t2263 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2947 uo_out[1].t3 _284_.ZN.t29 VGND.t6245 VGND.t6244 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2948 a_22300_24679# a_22212_24776# VGND.t2266 VGND.t2265 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2949 a_34304_24029# a_33932_24073# VPWR.t528 VPWR.t527 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X2950 VGND.t6654 _459_.Q.t8 a_35108_28776# VGND.t6653 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2951 VPWR.t5091 a_1468_19975# a_1380_20072# VPWR.t2297 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2952 a_45820_13703# a_45732_13800# VGND.t3045 VGND.t3044 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2953 a_44744_18559# a_42896_18504# a_44459_18559# VPWR.t5974 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X2954 VPWR.t3209 a_4828_29383# a_4740_29480# VPWR.t3208 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2955 a_22300_21543# a_22212_21640# VGND.t3051 VGND.t3050 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2956 a_28572_1592# a_28484_1636# VGND.t3053 VGND.t3052 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2957 a_3708_15271# a_3620_15368# VGND.t3543 VGND.t3542 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2958 a_45232_25987# a_44784_25987.t4 a_45644_26399# VPWR.t177 pfet_06v0 ad=0.1872p pd=1.4u as=43.2f ps=0.6u w=0.36u l=0.5u
X2959 _272_.A2 _228_.ZN a_58116_30344# VGND.t71 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2960 a_5500_1592# a_5412_1636# VGND.t3545 VGND.t3544 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2961 a_33052_16839# a_32964_16936# VGND.t3547 VGND.t3546 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2962 VPWR.t2313 a_46156_16839# a_46068_16936# VPWR.t2312 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2963 a_56124_28248# a_56036_28292# VGND.t3549 VGND.t3548 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2964 VPWR.t3294 a_50524_9432# a_50436_9476# VPWR.t3293 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2965 a_3708_12135# a_3620_12232# VGND.t2730 VGND.t2729 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2966 VPWR.t6124 a_11324_1159# a_11236_1256# VPWR.t6123 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2967 a_48820_28292# _383_.A2 a_48596_28292# VPWR.t1056 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2968 a_31803_24831# a_30240_24776# a_31168_24419# VGND.t6049 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2969 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I VGND.t2734 VGND.t2733 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2970 _465_.D uio_out[5].t9 VGND.t6585 VGND.t102 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X2971 VPWR.t2924 a_67212_10567# a_67124_10664# VPWR.t2923 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2972 VGND.t6147 a_52064_19715.t6 a_52024_20083# VGND.t6146 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2973 VPWR.t1718 a_67436_18407# a_67348_18504# VPWR.t1717 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2974 VPWR.t2944 a_4156_10567# a_4068_10664# VPWR.t2943 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2975 VGND.t25 a_53744_22851.t4 a_55116_22895# VGND.t24 nfet_06v0 ad=0.1584p pd=1.6u as=43.2f ps=0.6u w=0.36u l=0.6u
X2976 VPWR.t4261 a_2812_20408# a_2724_20452# VPWR.t4260 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2977 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t1271 VPWR.t1270 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2978 VPWR.t2854 a_48060_18407# a_47972_18504# VPWR.t2853 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2979 VPWR.t1760 a_56012_10567# a_55924_10664# VPWR.t1759 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2980 VPWR.t4263 a_29020_1159# a_28932_1256# VPWR.t4262 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2981 a_51308_18407# a_51220_18504# VGND.t4101 VGND.t4100 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2982 a_65308_8999# a_65220_9096# VGND.t4102 VGND.t3309 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2983 a_39324_17272# a_39236_17316# VGND.t4104 VGND.t4103 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2984 VPWR.t1724 a_50300_1592# a_50212_1636# VPWR.t1723 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2985 a_33764_24073# a_32964_24072.t5 VGND.t154 VGND.t153 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2986 a_25124_28776# _455_.Q.t7 a_27460_28776# VGND.t6536 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2987 VPWR.t3512 a_31708_18840# a_31620_18884# VPWR.t3511 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2988 VGND.t874 _250_.ZN a_60276_29032# VGND.t873 nfet_06v0 ad=0.104p pd=0.92u as=0.14p ps=1.1u w=0.4u l=0.6u
X2989 a_65308_5863# a_65220_5960# VGND.t3362 VGND.t3096 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2990 VPWR.t1496 a_31708_15704# a_31620_15748# VPWR.t1495 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2991 VPWR.t3862 a_2364_12568# a_2276_12612# VPWR.t54 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2992 a_15244_26247# a_15156_26344# VGND.t3363 VGND.t660 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2993 clkload0.Z a_48384_26724# VGND.t2864 VGND.t2863 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X2994 a_33724_2727# a_33636_2824# VGND.t3660 VGND.t666 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2995 VPWR.t3407 a_3708_9432# a_3620_9476# VPWR.t3406 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2996 a_43380_20452# _452_.Q.t10 a_43156_20452# VPWR.t6954 pfet_06v0 ad=0.4599p pd=1.935u as=0.33945p ps=1.715u w=1.095u l=0.5u
X2997 a_36084_23208# _312_.ZN VPWR.t5540 VPWR.t5539 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2998 a_15244_23111# a_15156_23208# VGND.t3661 VGND.t2343 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2999 _480_.Q a_43296_28733# VGND.t6037 VGND.t6036 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3000 uo_out[1].t0 _284_.ZN.t30 a_40196_29480# VPWR.t6518 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3001 VPWR.t5894 a_52764_2727# a_52676_2824# VPWR.t5893 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3002 VPWR.t3786 a_13788_29816# a_13700_29860# VPWR.t3785 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3003 VPWR.t1703 a_32828_1592# a_32740_1636# VPWR.t1702 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3004 VGND.t1699 a_44786_24120# a_44906_24164# VGND.t1698 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X3005 VPWR.t3977 a_44812_17272# a_44724_17316# VPWR.t3976 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3006 a_43248_28777# a_41028_28776.t4 a_43003_28409# VGND.t6777 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3007 VPWR.t1862 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_62864_25156# VPWR.t1861 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X3008 a_56796_1592# a_56708_1636# VGND.t3759 VGND.t3758 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3009 VPWR.t1841 a_14908_30951# a_14820_31048# VPWR.t1840 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3010 VPWR.t2175 a_17484_26247# a_17396_26344# VPWR.t2174 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3011 a_61500_26247# a_61412_26344# VGND.t3761 VGND.t3760 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3012 VPWR.t3909 a_2812_14136# a_2724_14180# VPWR.t3908 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3013 VGND.t6207 _459_.CLK.t29 a_21652_27591.t1 VGND.t6206 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3014 VPWR.t3189 a_4156_8999# a_4068_9096# VPWR.t3188 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3015 a_48844_16839# a_48756_16936# VGND.t3807 VGND.t3806 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3016 VPWR.t3574 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I VPWR.t3573 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3017 VGND.t4858 _475_.Q _421_.B VGND.t4857 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X3018 VPWR.t2965 a_17484_23111# a_17396_23208# VPWR.t1901 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3019 VPWR.t3956 a_2812_11000# a_2724_11044# VPWR.t3955 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3020 VGND.t105 _294_.A2.t4 _290_.ZN VGND.t104 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X3021 a_16796_27209# _467_.D a_16672_26841# VPWR.t1023 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X3022 a_1468_29383# a_1380_29480# VGND.t3809 VGND.t3672 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3023 a_39780_22805# _441_.B VGND.t5090 VGND.t5089 nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3024 VPWR.t6475 _459_.CLK.t30 a_26916_25640.t0 VPWR.t6474 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3025 vgaringosc.workerclkbuff_notouch_.I.t2 _274_.ZN a_51665_30344# VGND.t199 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X3026 VPWR.t5683 a_33276_1159# a_33188_1256# VPWR.t4300 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3027 VPWR.t3627 a_56796_12568# a_56708_12612# VPWR.t3626 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3028 VGND.t6305 _447_.Q.t7 _319_.A2 VGND.t6304 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X3029 _301_.Z a_38340_21327# VGND.t4982 VGND.t4981 nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X3030 a_30628_24463# a_29828_24455.t4 VGND.t6118 VGND.t6117 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3031 VPWR.t5294 a_61388_16839# a_61300_16936# VPWR.t5293 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3032 a_62620_15271# a_62532_15368# VGND.t5486 VGND.t5485 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3033 a_21424_25987# a_21052_26031# VPWR.t1412 VPWR.t1411 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X3034 a_25867_26841# a_23892_27208.t4 a_25232_27165# VPWR.t6340 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X3035 VPWR.t2432 a_20060_24679# a_19972_24776# VPWR.t2431 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3036 VPWR.t2840 a_64860_6296# a_64772_6340# VPWR.t2839 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3037 VPWR.t2842 a_49292_12135# a_49204_12232# VPWR.t2841 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3038 VPWR.t5702 a_37360_19325# a_37352_19001# VPWR.t5701 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X3039 a_59260_23544# a_59172_23588# VGND.t2704 VGND.t2703 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3040 VGND.t1061 a_65072_29860# _324_.C.t5 VGND.t1059 nfet_06v0 ad=0.2002p pd=1.79u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3041 VPWR.t307 a_64860_3160# a_64772_3204# VPWR.t306 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3042 _241_.I0 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I VPWR.t3506 VPWR.t3505 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3043 a_40220_15271# a_40132_15368# VGND.t2706 VGND.t2705 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3044 a_61948_2727# a_61860_2824# VGND.t3235 VGND.t3234 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3045 VPWR.t3386 a_46268_12135# a_46180_12232# VPWR.t3385 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3046 a_56236_23544# a_56148_23588# VGND.t3238 VGND.t3237 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3047 a_57580_17272# a_57492_17316# VGND.t3240 VGND.t3239 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3048 a_65756_17272# a_65668_17316# VGND.t3242 VGND.t3241 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3049 a_59572_29076# _247_.ZN _258_.I VGND.t1811 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3050 a_36060_19369# _448_.D a_35936_19001# VPWR.t638 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X3051 a_49496_30345# a_49112_29885# a_48708_29816# VGND.t137 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3052 _258_.I _257_.B VPWR.t315 VPWR.t314 pfet_06v0 ad=0.4016p pd=1.94u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3053 _350_.A2.t12 _371_.A1.t15 a_30388_28776# VGND.t6235 nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3054 a_4156_19975# a_4068_20072# VGND.t2231 VGND.t1030 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3055 VPWR.t1728 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN VPWR.t1727 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3056 a_64412_7864# a_64324_7908# VGND.t2233 VGND.t2232 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3057 VGND.t5657 _441_.ZN _442_.ZN VGND.t5656 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3058 a_36524_18407# a_36436_18504# VGND.t2235 VGND.t2234 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3059 a_30812_19975# a_30724_20072# VGND.t2236 VGND.t1036 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3060 VPWR.t5902 a_17036_25112# a_16948_25156# VPWR.t5901 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3061 a_34700_28776# _459_.Q.t9 VGND.t6656 VGND.t6655 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3062 a_41788_15704# a_41700_15748# VGND.t2792 VGND.t2791 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3063 a_41440_23208# _260_.A1 a_41216_23208# VPWR.t3914 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3064 a_55312_22340# a_54824_22045# a_55744_22505# VGND.t3795 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X3065 a_55676_2727# a_55588_2824# VGND.t2794 VGND.t2793 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3066 a_64412_4728# a_64324_4772# VGND.t2796 VGND.t2795 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3067 VPWR.t388 a_53660_15271# a_53572_15368# VPWR.t387 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3068 VPWR.t6701 vgaringosc.workerclkbuff_notouch_.I.t7 a_41048_29816.t2 VPWR.t6700 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X3069 VPWR.t6423 _451_.Q.t4 a_38340_21327# VPWR.t6422 pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X3070 VPWR.t4341 a_30140_23111# a_30052_23208# VPWR.t4340 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3071 VPWR.t2903 a_3260_28248# a_3172_28292# VPWR.t2885 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3072 a_2364_2727# a_2276_2824# VGND.t2769 VGND.t347 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3073 a_32156_17272# a_32068_17316# VGND.t2771 VGND.t2770 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3074 VPWR.t2907 a_1468_4728# a_1380_4772# VPWR.t1459 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3075 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I VPWR.t2368 VPWR.t2367 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3076 _229_.I.t1 a_62532_30736# VGND.t2404 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X3077 vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN VPWR.t3113 VPWR.t3112 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3078 VPWR.t3109 a_47612_12568# a_47524_12612# VPWR.t1391 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3079 a_39781_24372# _431_.A3 a_39587_24372# VGND.t2058 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X3080 VPWR.t3498 a_3260_25112# a_3172_25156# VPWR.t3497 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3081 a_28432_29535# a_28000_29480# VPWR.t1930 VPWR.t1929 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X3082 VPWR.t1570 a_31260_15271# a_31172_15368# VPWR.t1569 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3083 VPWR.t1365 a_1468_1592# a_1380_1636# VPWR.t1364 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3084 vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN VPWR.t1367 VPWR.t1366 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3085 VPWR.t5904 a_52204_16839# a_52116_16936# VPWR.t5903 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3086 a_12892_1159# a_12804_1256# VGND.t2748 VGND.t2747 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3087 VPWR.t1267 _399_.ZN _427_.A2 VPWR.t1266 pfet_06v0 ad=0.2561p pd=1.505u as=0.4016p ps=1.94u w=0.985u l=0.5u
X3088 _319_.A2 _447_.Q.t8 a_37744_20452# VPWR.t6582 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X3089 a_61297_30300# _230_.I.t6 VGND.t6346 VGND.t1077 nfet_06v0 ad=93.59999f pd=0.88u as=0.2288p ps=1.58u w=0.36u l=0.6u
X3090 a_41804_19376# _327_.A2 a_41600_19376# VGND.t3249 nfet_06v0 ad=60.8f pd=0.7u as=79.8f ps=0.8u w=0.38u l=0.6u
X3091 VPWR.t5748 a_41004_16839# a_40916_16936# VPWR.t5747 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3092 VPWR.t1953 a_47164_30951# a_47076_31048# VPWR.t1952 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3093 VPWR.t2177 a_55788_23544# a_55700_23588# VPWR.t2176 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3094 a_33520_25597# a_33148_25641# VGND.t5891 VGND.t5890 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X3095 VPWR.t4696 _304_.B _281_.ZN.t3 VPWR.t4695 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3096 a_38325_22804# _447_.Q.t9 a_38131_22804# VGND.t6306 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X3097 _459_.Q.t0 a_32096_24419# VPWR.t2784 VPWR.t2783 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3098 VPWR.t4214 a_67548_6296# a_67460_6340# VPWR.t4213 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3099 a_35184_24073# a_32964_24072.t6 a_34939_23705# VGND.t155 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3100 VGND.t3520 a_19035_28409# a_19328_28733# VGND.t3519 nfet_06v0 ad=0.2608p pd=1.455u as=0.2119p ps=1.335u w=0.815u l=0.6u
X3101 VGND.t6390 _355_.C.t10 _459_.D VGND.t6389 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X3102 VPWR.t6723 _402_.A1.t14 _383_.A2 VPWR.t6722 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3103 VPWR.t6597 a_54864_22461.t4 a_54824_22045# VPWR.t6596 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3104 a_49740_29383# a_49652_29480# VGND.t4093 VGND.t4092 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3105 a_32604_15704# a_32516_15748# VGND.t4095 VGND.t4094 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3106 a_16028_29816# a_15940_29860# VGND.t4096 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3107 VPWR.t1176 a_67548_3160# a_67460_3204# VPWR.t1175 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3108 a_24080_25227# a_23668_25640.t3 VPWR.t7028 VPWR.t7027 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3109 a_1020_26680# a_932_26724# VGND.t5276 VGND.t4712 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3110 a_38576_22504# _447_.Q.t10 VPWR.t6584 VPWR.t6583 pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X3111 a_41099_26841# a_39124_27208.t4 a_40464_27165# VPWR.t221 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X3112 a_47524_22021# _474_.Q _421_.B VPWR.t4797 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3113 a_3708_4295# a_3620_4392# VGND.t5281 VGND.t4938 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3114 a_5388_13703# a_5300_13800# VGND.t5283 VGND.t5282 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3115 VPWR.t5469 a_59260_26680# a_59172_26724# VPWR.t5468 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3116 a_34292_28776# _460_.Q a_34084_28776# VGND.t3334 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3117 VGND.t2032 a_36432_19325# a_36384_19369# VGND.t2031 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X3118 VGND.t6272 a_48272_25156.t27 _474_.CLK.t13 VGND.t6271 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3119 a_11548_1592# a_11460_1636# VGND.t5071 VGND.t5070 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3120 _287_.A1.t5 a_38472_30169# VGND.t4814 VGND.t1059 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3121 VPWR.t1671 a_67660_10567# a_67572_10664# VPWR.t1670 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3122 VGND.t2942 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN VGND.t2941 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3123 VPWR.t1673 a_67884_18407# a_67796_18504# VPWR.t1672 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3124 VPWR.t3216 a_5388_8999# a_5300_9096# VPWR.t3215 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3125 VPWR.t7015 _251_.A1.t18 _228_.ZN VPWR.t7014 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3126 VGND.t4056 _336_.A1 _355_.B VGND.t4055 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X3127 a_35516_1592# a_35428_1636# VGND.t5073 VGND.t5072 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3128 a_47600_27912# _404_.A1 a_47376_27912# VPWR.t3825 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3129 VPWR.t3441 a_30812_1592# a_30724_1636# VPWR.t1114 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3130 vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN VPWR.t2858 VPWR.t2857 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3131 VGND.t6508 _324_.C.t19 a_51988_24072# VGND.t186 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3132 VPWR.t5767 a_56460_10567# a_56372_10664# VPWR.t5766 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3133 a_51532_10567# a_51444_10664# VGND.t5319 VGND.t5318 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3134 VPWR.t6328 a_56684_18407# a_56596_18504# VPWR.t6327 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3135 _451_.Q.t0 a_39264_18147# VPWR.t6265 VPWR.t6264 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3136 a_51756_18407# a_51668_18504# VGND.t5321 VGND.t5320 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3137 a_54432_31128# ui_in[7].t2 VGND.t7 VGND.t6 nfet_06v0 ad=0.2662p pd=2.09u as=0.2662p ps=2.09u w=0.605u l=0.6u
X3138 VPWR.t5735 a_25212_2727# a_25124_2824# VPWR.t5734 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3139 a_54780_1592# a_54692_1636# VGND.t5287 VGND.t440 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3140 VPWR.t6634 _230_.I.t7 _243_.B2 VPWR.t6633 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3141 a_19716_29977# a_18404_30344.t3 a_19372_30345# VPWR.t137 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X3142 uio_out[5].t1 a_20672_30301# VPWR.t5017 VPWR.t5016 pfet_06v0 ad=0.4392p pd=1.94u as=0.38575p ps=1.92u w=1.22u l=0.5u
X3143 VPWR.t2341 a_64412_7864# a_64324_7908# VPWR.t2340 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3144 VPWR.t1414 a_21068_25112# a_20980_25156# VPWR.t1413 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3145 a_18264_29480# uio_out[7].t10 _379_.Z VPWR.t6896 pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3146 VPWR.t1805 a_24540_1592# a_24452_1636# VPWR.t1804 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3147 VPWR.t1807 a_49180_15704# a_49092_15748# VPWR.t1806 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3148 hold2.I hold1.Z a_42161_24776# VPWR.t3569 pfet_06v0 ad=0.3159p pd=1.735u as=0.32805p ps=1.755u w=1.215u l=0.5u
X3149 a_21404_1159# a_21316_1256# VGND.t5291 VGND.t5290 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3150 VPWR.t4609 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN VPWR.t4608 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3151 a_15692_26247# a_15604_26344# VGND.t5058 VGND.t4828 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3152 a_23868_26247# a_23780_26344# VGND.t5060 VGND.t5059 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3153 VPWR.t3236 a_50384_19204# a_50280_19369# VPWR.t3235 pfet_06v0 ad=0.1044p pd=0.94u as=0.1791p ps=1.355u w=0.36u l=0.5u
X3154 a_52064_19715.t1 _474_.CLK.t39 VGND.t6453 VGND.t6452 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3155 a_26427_29977# a_24452_30344.t5 a_25792_30301# VPWR.t160 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X3156 VPWR.t2494 a_62844_12568# a_62756_12612# VPWR.t2493 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3157 VPWR.t1961 a_20508_23111# a_20420_23208# VPWR.t1960 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3158 _459_.Q.t1 a_32096_24419# VGND.t2643 VGND.t2642 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3159 a_15692_23111# a_15604_23208# VGND.t5063 VGND.t5062 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3160 VGND.t6669 _352_.A2.t23 a_31116_26020# VGND.t6668 nfet_06v0 ad=0.2424p pd=1.635u as=79.8f ps=0.8u w=0.38u l=0.6u
X3161 a_43664_29535# a_43232_29480# VPWR.t806 VPWR.t805 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X3162 a_3708_28248# a_3620_28292# VGND.t3502 VGND.t3501 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3163 _249_.A2 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN VGND.t1459 VGND.t71 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3164 VPWR.t5760 a_37420_16839# a_37332_16936# VPWR.t5759 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3165 a_37408_18504# a_36996_18183.t6 VGND.t6632 VGND.t6631 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3166 VPWR.t2627 a_51644_12568# a_51556_12612# VPWR.t2626 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3167 a_4940_18407# a_4852_18504# VGND.t3504 VGND.t3503 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3168 a_56804_30344# _258_.I _274_.A2 VGND.t325 nfet_06v0 ad=85.2f pd=0.95u as=0.3124p ps=2.3u w=0.71u l=0.6u
X3169 _455_.Q.t0 a_22352_25987# VPWR.t4007 VPWR.t4006 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3170 VPWR.t6687 a_41048_29816.t11 _459_.CLK.t5 VPWR.t6686 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3171 a_1916_18407# a_1828_18504# VGND.t2850 VGND.t2849 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3172 _475_.D _421_.B VGND.t3042 VGND.t3041 nfet_06v0 ad=0.21175p pd=1.41u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3173 VPWR.t6971 _459_.Q.t10 _371_.A3 VPWR.t6970 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3174 _454_.Q a_23920_27555# VPWR.t613 VPWR.t612 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3175 _284_.B _397_.A2.t9 a_47636_25940# VGND.t6723 nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3176 VPWR.t3939 a_52988_9432# a_52900_9476# VPWR.t3938 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3177 a_10428_2727# a_10340_2824# VGND.t2852 VGND.t2851 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3178 VPWR.t2989 a_13788_1159# a_13700_1256# VPWR.t389 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3179 a_45396_25156# _304_.B _284_.ZN.t13 VPWR.t4694 pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X3180 _247_.B _245_.Z a_59828_26724# VPWR.t6087 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3181 VGND.t5793 a_19328_28733# uio_out[6].t5 VGND.t5792 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X3182 a_44786_24120# hold2.I VGND.t2416 VGND.t2415 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3183 VGND.t6403 a_41048_29816.t12 _459_.CLK.t13 VGND.t6400 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3184 VPWR.t133 _417_.A2.t7 a_49034_21640# VPWR.t132 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X3185 a_53660_2727# a_53572_2824# VGND.t4500 VGND.t4499 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3186 VGND.t3739 _241_.I0 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I VGND.t3738 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3187 a_2812_3160# a_2724_3204# VGND.t4501 VGND.t4200 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3188 a_44302_23588# a_44162_24120# VPWR.t4979 VPWR.t4978 pfet_06v0 ad=61.19999f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X3189 VGND.t6694 _251_.A1.t19 a_56404_27208# VGND.t6693 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3190 a_19204_30345# a_18404_30344.t4 VGND.t138 VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3191 _452_.CLK.t8 a_42392_22825.t22 VPWR.t6918 VPWR.t6917 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3192 a_53260_26399# a_52744_26031# VPWR.t5791 VPWR.t5790 pfet_06v0 ad=43.2f pd=0.6u as=0.1044p ps=0.94u w=0.36u l=0.5u
X3193 a_28124_2727# a_28036_2824# VGND.t5580 VGND.t3947 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3194 a_6844_29816# a_6756_29860# VGND.t5581 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3195 _473_.Q a_47552_19715# VGND.t1828 VGND.t1827 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3196 VPWR.t3682 a_23196_2727# a_23108_2824# VPWR.t3681 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3197 VPWR.t5797 a_37532_21543# a_37444_21640# VPWR.t5796 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3198 a_3708_18840# a_3620_18884# VGND.t5584 VGND.t4127 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3199 VPWR.t5854 a_47164_2727# a_47076_2824# VPWR.t5853 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3200 _400_.ZN _402_.A1.t15 VPWR.t6725 VPWR.t6724 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3201 a_56684_23544# a_56596_23588# VGND.t5586 VGND.t5585 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3202 VPWR.t1878 a_27228_1592# a_27140_1636# VPWR.t1877 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3203 a_4156_1592# a_4068_1636# VGND.t5587 VGND.t4129 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3204 a_52316_27815# a_52228_27912# VGND.t5589 VGND.t5588 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3205 VPWR.t5808 a_38816_27555# a_38808_27967# VPWR.t5807 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X3206 VPWR.t1477 a_17484_25112# a_17396_25156# VPWR.t1476 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3207 VPWR.t2717 a_46492_1592# a_46404_1636# VPWR.t2716 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3208 _272_.B1 _474_.CLK.t40 VGND.t6454 VGND.t102 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X3209 a_60604_9432# a_60516_9476# VGND.t5595 VGND.t5594 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3210 VPWR.t2753 a_61836_23544# a_61748_23588# VPWR.t2752 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3211 VGND.t6255 _362_.B.t11 _362_.ZN VGND.t6254 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X3212 a_56964_26724# a_56404_27208# a_56836_27208# VGND.t5530 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X3213 VPWR.t4259 a_16028_29816# a_15940_29860# VPWR.t4258 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3214 a_33948_18407# a_33860_18504# VGND.t5565 VGND.t5441 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3215 _242_.Z a_56516_26344# VGND.t332 VGND.t331 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3216 VPWR.t5779 a_27228_26680# a_27140_26724# VPWR.t4994 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3217 _234_.ZN _436_.B VPWR.t5870 VPWR.t5869 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3218 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I _249_.A2 VPWR.t1531 VPWR.t1530 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3219 a_23084_23544# a_22996_23588# VGND.t5569 VGND.t5568 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3220 VPWR.t5785 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I VPWR.t5784 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3221 _421_.A1 _324_.B.t26 VGND.t6417 VGND.t6416 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3222 a_54332_9432# a_54244_9476# VGND.t5575 VGND.t5574 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3223 a_33492_25273# a_32180_25640.t5 a_33148_25641# VPWR.t39 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X3224 a_59372_14136# a_59284_14180# VGND.t1519 VGND.t1518 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3225 VPWR.t2710 a_61388_15704# a_61300_15748# VPWR.t2709 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3226 VPWR.t2712 a_39548_15704# a_39460_15748# VPWR.t2711 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3227 VPWR.t3419 a_52652_16839# a_52564_16936# VPWR.t3418 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3228 a_1020_9432# a_932_9476# VGND.t5576 VGND.t3890 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3229 VPWR.t2790 a_5948_1592# a_5860_1636# VPWR.t2789 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3230 VPWR.t5942 a_65084_15271# a_64996_15368# VPWR.t5941 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3231 a_3260_13703# a_3172_13800# VGND.t5577 VGND.t4899 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3232 a_56348_14136# a_56260_14180# VGND.t1066 VGND.t1065 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3233 a_48060_9432# a_47972_9476# VGND.t2334 VGND.t2333 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3234 VPWR.t2461 a_46268_14136# a_46180_14180# VPWR.t393 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3235 VPWR.t3822 a_41452_16839# a_41364_16936# VPWR.t3821 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3236 a_1020_6296# a_932_6340# VGND.t353 VGND.t352 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3237 a_47552_19715# a_47259_20127# VGND.t2338 VGND.t2337 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X3238 VPWR.t44 _363_.Z.t4 a_33140_29860# VPWR.t43 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3239 a_56348_11000# a_56260_11044# VGND.t5075 VGND.t5074 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3240 VPWR.t2465 a_46268_11000# a_46180_11044# VPWR.t2464 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3241 VPWR.t4707 a_59036_12568# a_58948_12612# VPWR.t4706 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3242 a_15244_26680# a_15156_26724# VGND.t2342 VGND.t2341 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3243 a_42368_28733# a_41996_28777# VPWR.t2980 VPWR.t2979 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X3244 a_67772_24679# a_67684_24776# VGND.t5026 VGND.t5025 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3245 VGND.t180 _384_.A3.t13 a_51240_23340# VGND.t179 nfet_06v0 ad=93.59999f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X3246 VGND.t1922 a_37472_24419# a_37424_24463# VGND.t1921 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X3247 a_25212_1159# a_25124_1256# VGND.t5497 VGND.t5496 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3248 a_33724_1159# a_33636_1256# VGND.t1719 VGND.t1718 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3249 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I VPWR.t1770 VPWR.t1769 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3250 VPWR.t5960 a_49628_17272# a_49540_17316# VPWR.t5959 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3251 VGND.t474 _358_.A3 _459_.D VGND.t473 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3252 a_36300_23544# a_36212_23588# VGND.t5032 VGND.t5031 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3253 a_3708_30951# a_3620_31048# VGND.t5033 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3254 a_30388_28776# _337_.ZN _350_.A2.t5 VGND.t4978 nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X3255 a_67772_21543# a_67684_21640# VGND.t5222 VGND.t5221 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3256 VPWR.t6034 a_35008_22461# a_35000_22137# VPWR.t6033 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X3257 VPWR.t4676 a_54432_31128# _304_.B VPWR.t4675 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3258 a_42778_21812# a_42154_21236# a_42630_21236# VGND.t2379 nfet_06v0 ad=0.369p pd=2.77u as=43.2f ps=0.6u w=0.36u l=0.6u
X3259 a_53548_24679# a_53460_24776# VGND.t5224 VGND.t5223 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3260 VPWR.t5351 a_22188_30951# a_22100_31048# VPWR.t5350 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3261 a_55228_15704# a_55140_15748# VGND.t5226 VGND.t5225 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3262 VPWR.t3167 a_2812_16839# a_2724_16936# VPWR.t3166 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3263 _249_.A2 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN VPWR.t1525 VPWR.t1524 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3264 a_34155_25273# a_32592_25227# a_33520_25597# VGND.t5690 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3265 VGND.t2819 a_43936_27165# a_43888_27209# VGND.t2818 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X3266 VPWR.t1924 a_47552_19715# a_47544_20127# VPWR.t1923 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X3267 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I VPWR.t509 VPWR.t508 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3268 VGND.t4910 a_24952_29032# _343_.A2 VGND.t4909 nfet_06v0 ad=0.23405p pd=1.555u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3269 a_44028_15704# a_43940_15748# VGND.t4189 VGND.t4188 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3270 a_65868_13703# a_65780_13800# VGND.t4191 VGND.t4190 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3271 _392_.A2 _384_.ZN VPWR.t3181 VPWR.t3180 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3272 VPWR.t1217 _248_.B1 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t1216 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3273 VGND.t6273 a_48272_25156.t28 _474_.CLK.t14 VGND.t2353 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3274 a_54668_13703# a_54580_13800# VGND.t4195 VGND.t4194 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3275 a_62620_18840# a_62532_18884# VGND.t5268 VGND.t4739 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3276 _260_.A1 _327_.A2 VPWR.t3400 VPWR.t3397 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3277 VGND.t2262 a_25792_30301# a_25744_30345# VGND.t137 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X3278 a_51980_10567# a_51892_10664# VGND.t5270 VGND.t5269 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3279 _294_.ZN.t0 _294_.A2.t5 VGND.t107 VGND.t106 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X3280 _358_.A3 a_30724_26020# VGND.t1039 VGND.t1038 nfet_06v0 ad=0.341p pd=2.43u as=0.2424p ps=1.635u w=0.775u l=0.6u
X3281 a_37067_19001# a_35504_18955# a_36432_19325# VGND.t1262 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3282 a_16240_26795# a_15828_27208.t5 VPWR.t6384 VPWR.t6383 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3283 uio_out[5].t0 a_20672_30301# VPWR.t5015 VPWR.t5014 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3284 a_62404_25640# _245_.I1 VGND.t5230 VGND.t5229 nfet_06v0 ad=98.39999f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3285 a_48060_12135# a_47972_12232# VGND.t5271 VGND.t5038 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3286 _436_.ZN _435_.ZN a_40357_24776# VPWR.t4830 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3287 _362_.ZN _460_.Q a_32836_27208# VGND.t3333 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3288 a_66204_1159# a_66116_1256# VGND.t4406 VGND.t4405 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3289 a_3708_24679# a_3620_24776# VGND.t4408 VGND.t4407 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3290 _313_.ZN _312_.ZN VGND.t5345 VGND.t5344 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X3291 VGND.t1521 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I VGND.t1520 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3292 _474_.CLK.t15 a_48272_25156.t29 VPWR.t6559 VPWR.t6558 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3293 VGND.t4813 a_38472_30169# _287_.A1.t4 VGND.t1059 nfet_06v0 ad=0.23432p pd=1.94u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3294 VPWR.t1803 a_50972_9432# a_50884_9476# VPWR.t1802 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3295 a_53300_23047# a_53704_23219# a_53648_23263# VPWR.t3985 pfet_06v0 ad=0.1665p pd=1.285u as=50.4f ps=0.64u w=0.36u l=0.5u
X3296 VPWR.t6714 _324_.B.t27 a_48321_23208# VPWR.t6713 pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3297 VPWR.t4556 a_11772_1159# a_11684_1256# VPWR.t4555 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3298 a_3708_21543# a_3620_21640# VGND.t4629 VGND.t2883 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3299 VPWR.t1396 a_20956_23111# a_20868_23208# VPWR.t1395 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3300 VPWR.t4438 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t4437 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3301 VGND.t213 _330_.A1.t13 _443_.D VGND.t212 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X3302 VPWR.t5795 a_6844_29816# a_6756_29860# VPWR.t5794 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3303 a_49152_30301.t0 _474_.CLK.t41 VPWR.t6751 VPWR.t6750 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3304 uio_out[6].t1 a_19328_28733# VPWR.t6045 VPWR.t6044 pfet_06v0 ad=0.4392p pd=1.94u as=0.38575p ps=1.92u w=1.22u l=0.5u
X3305 VPWR.t4782 a_35740_1159# a_35652_1256# VPWR.t4781 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3306 VPWR.t2002 a_37384_19624# _325_.A2.t0 VPWR.t2001 pfet_06v0 ad=0.40575p pd=2.055u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3307 VPWR.t1408 a_13004_30951# a_12916_31048# VPWR.t1407 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3308 a_61724_1592# a_61636_1636# VGND.t4633 VGND.t4632 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3309 a_2364_20408# a_2276_20452# VGND.t3849 VGND.t640 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3310 a_25252_30345# a_24452_30344.t6 VGND.t157 VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3311 VPWR.t2935 a_51420_2727# a_51332_2824# VPWR.t2934 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3312 VPWR.t2339 a_4156_19975# a_4068_20072# VPWR.t2338 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3313 VPWR.t5180 a_7516_29383# a_7428_29480# VPWR.t5179 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3314 VPWR.t2345 a_30812_19975# a_30724_20072# VPWR.t2344 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3315 a_65756_8999# a_65668_9096# VGND.t5021 VGND.t5020 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3316 _352_.A2.t7 _371_.A2 VGND.t3433 VGND.t3432 nfet_06v0 ad=0.1326p pd=1.03u as=0.2244p ps=1.9u w=0.51u l=0.6u
X3317 VPWR.t2141 a_56684_17272# a_56596_17316# VPWR.t2140 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3318 a_20853_30644# uio_out[6].t10 VGND.t6590 VGND.t34 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3319 a_65756_5863# a_65668_5960# VGND.t5022 VGND.t966 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3320 _352_.ZN _336_.A2.t7 a_26756_24801# VPWR.t171 pfet_06v0 ad=0.31207p pd=1.665u as=0.55297p ps=2.105u w=1.095u l=0.5u
X3321 VPWR.t6194 a_62508_13703# a_62420_13800# VPWR.t6193 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3322 VPWR.t5109 a_2364_21976# a_2276_22020# VPWR.t641 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3323 VGND.t259 clkbuf_1_0__f_clk.I.t45 a_42392_22825.t10 VGND.t258 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3324 VPWR.t1321 vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t1320 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3325 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _275_.A2 VGND.t2628 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3326 _452_.CLK.t9 a_42392_22825.t23 VPWR.t6920 VPWR.t6919 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3327 a_59708_23111# a_59620_23208# VGND.t4956 VGND.t4955 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3328 VPWR.t2155 a_27676_2727# a_27588_2824# VPWR.t2154 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3329 VPWR.t5115 vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN VPWR.t5114 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3330 a_2364_14136# a_2276_14180# VGND.t743 VGND.t742 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3331 _300_.A2 _448_.Q.t6 VPWR.t6887 VPWR.t6886 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3332 a_36116_29167# a_35316_29159.t2 VGND.t6738 VGND.t6737 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3333 VGND.t6362 _452_.CLK.t44 a_45508_20936.t1 VGND.t6361 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3334 a_47733_29098# _386_.ZN VGND.t1784 VGND.t1783 nfet_06v0 ad=85.2f pd=0.95u as=0.3124p ps=2.3u w=0.71u l=0.6u
X3335 a_2364_11000# a_2276_11044# VGND.t5614 VGND.t1049 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3336 _231_.I vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN VGND.t542 VGND.t541 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3337 a_37532_1159# a_37444_1256# VGND.t5259 VGND.t5258 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3338 VPWR.t1784 a_5052_12568# a_4964_12612# VPWR.t1783 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3339 a_29020_1159# a_28932_1256# VGND.t4099 VGND.t4098 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3340 a_52764_27815# a_52676_27912# VGND.t5261 VGND.t5260 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3341 a_59948_30352# _256_.A2.t2 a_59744_30352# VGND.t3682 nfet_06v0 ad=60.8f pd=0.7u as=79.8f ps=0.8u w=0.38u l=0.6u
X3342 VPWR.t5445 a_67996_21976# a_67908_22020# VPWR.t5444 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3343 VPWR.t7095 _256_.A2.t3 a_59332_29816# VPWR.t7094 pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X3344 VGND.t1447 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN VGND.t1446 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3345 a_30364_2727# a_30276_2824# VGND.t3178 VGND.t3177 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3346 VPWR.t3330 a_38428_1159# a_38340_1256# VPWR.t3329 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3347 a_52092_15271# a_52004_15368# VGND.t3182 VGND.t3181 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3348 a_47544_20127# a_45696_20072# a_47259_20127# VPWR.t2597 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X3349 a_53280_26031# a_52744_26031# VGND.t5579 VGND.t5578 nfet_06v0 ad=43.2f pd=0.6u as=0.2637p ps=1.825u w=0.36u l=0.6u
X3350 a_56816_26724# _241_.I0 VPWR.t3881 VPWR.t3880 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3351 a_59372_10567# a_59284_10664# VGND.t3184 VGND.t3183 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3352 VPWR.t3335 a_27676_26680# a_27588_26724# VPWR.t361 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3353 a_38428_15271# a_38340_15368# VGND.t5006 VGND.t5005 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3354 _478_.D _398_.C a_52852_24372# VGND.t3155 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3355 VPWR.t5169 a_40780_27815# a_40692_27912# VPWR.t5168 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3356 a_54332_2727# a_54244_2824# VGND.t5009 VGND.t3458 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3357 VPWR.t3141 a_40038_28720# uo_out[7].t1 VPWR.t3140 pfet_06v0 ad=0.4941p pd=2.03u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3358 vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t2276 VGND.t2275 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3359 a_60268_12135# a_60180_12232# VGND.t5011 VGND.t5010 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3360 VGND.t5994 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN VGND.t5993 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3361 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I VGND.t5015 VGND.t5014 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3362 VPWR.t5139 _337_.ZN a_31068_28292# VPWR.t5138 pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X3363 _371_.A3 _223_.I a_31031_27208# VGND.t6792 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X3364 VPWR.t2870 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN VPWR.t2869 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3365 VPWR.t3075 a_17148_29383# a_17060_29480# VPWR.t3074 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3366 a_1020_2727# a_932_2824# VGND.t2923 VGND.t2922 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3367 a_2812_12568# a_2724_12612# VGND.t2925 VGND.t2924 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3368 VPWR.t2053 a_39996_15704# a_39908_15748# VPWR.t2052 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3369 VGND.t5725 _412_.B2 a_51332_24372# VGND.t130 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3370 VPWR.t2055 a_53436_1592# a_53348_1636# VPWR.t2054 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3371 a_52964_29480# _268_.A1.t4 VPWR.t6737 VPWR.t6736 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3372 VPWR.t6229 a_1468_24679# a_1380_24776# VPWR.t4417 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3373 a_48060_2727# a_47972_2824# VGND.t3174 VGND.t2969 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3374 VPWR.t5936 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN VPWR.t5935 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3375 a_56796_14136# a_56708_14180# VGND.t1806 VGND.t1805 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3376 VPWR.t1713 a_28348_23111# a_28260_23208# VPWR.t1712 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3377 VGND.t2332 _264_.B hold2.I VGND.t2331 nfet_06v0 ad=0.23975p pd=1.475u as=0.1469p ps=1.085u w=0.565u l=0.6u
X3378 a_57276_27208# _251_.A1.t20 a_56964_26724# VGND.t6695 nfet_06v0 ad=98.39999f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3379 a_47689_25156# _279_.Z VPWR.t5588 VPWR.t5587 pfet_06v0 ad=0.1469p pd=1.085u as=0.38705p ps=2.08u w=0.565u l=0.5u
X3380 a_67861_31220# a_67741_30600# a_67117_30600# VPWR.t3323 pfet_06v0 ad=61.19999f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3381 a_60401_30300# _237_.A1 a_60793_29860# VPWR.t1130 pfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.5u
X3382 VPWR.t109 _294_.A2.t6 a_30778_31048# VPWR.t108 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X3383 a_56796_11000# a_56708_11044# VGND.t1819 VGND.t1818 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3384 a_28903_24776# _352_.A2.t24 _355_.ZN VPWR.t6990 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3385 a_4156_29383# a_4068_29480# VGND.t3287 VGND.t483 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3386 VPWR.t4862 a_59484_12568# a_59396_12612# VPWR.t4861 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3387 a_64860_7864# a_64772_7908# VGND.t3289 VGND.t3288 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3388 VGND.t6633 a_49152_30301.t4 a_49112_29885# VGND.t139 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3389 VPWR.t1429 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN VPWR.t1428 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3390 a_47525_29480# _384_.ZN _393_.A1 VPWR.t3179 pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3391 a_51428_23340# _384_.A1 a_51240_23340# VPWR.t938 pfet_06v0 ad=0.196p pd=1.26u as=0.2464p ps=2u w=0.56u l=0.5u
X3392 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t2358 VGND.t71 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3393 VGND.t6527 clk.t6 a_44296_24393.t6 VGND.t6526 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3394 VPWR.t1782 a_58924_13703# a_58836_13800# VPWR.t1781 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3395 VPWR.t2157 a_64076_16839# a_63988_16936# VPWR.t2156 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3396 VPWR.t3435 a_62732_26680# a_62644_26724# VPWR.t3434 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3397 a_60716_13703# a_60628_13800# VGND.t5918 VGND.t5917 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3398 a_64860_4728# a_64772_4772# VGND.t5919 VGND.t4604 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3399 _470_.Q a_44864_27165# VGND.t3225 VGND.t3224 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3400 a_38304_20072# _319_.A3 VPWR.t2707 VPWR.t2706 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3401 a_53648_23263# a_52920_22760# VPWR.t1293 VPWR.t1292 pfet_06v0 ad=50.4f pd=0.64u as=0.23p ps=1.54u w=0.36u l=0.5u
X3402 VPWR.t6183 a_23308_20408# a_23220_20452# VPWR.t6182 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3403 _243_.ZN _243_.A1 a_58228_27912# VPWR.t6037 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3404 a_7516_2727# a_7428_2824# VGND.t5923 VGND.t5922 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3405 a_32132_27912# _287_.A2 VPWR.t2028 VPWR.t2027 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X3406 VPWR.t6186 a_66204_6296# a_66116_6340# VPWR.t1208 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3407 a_53996_24679# a_53908_24776# VGND.t5869 VGND.t5868 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3408 _284_.ZN.t6 hold2.I VPWR.t2544 VPWR.t2543 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3409 VGND.t3 a_59332_29816# _267_.A2 VGND.t2 nfet_06v0 ad=0.2424p pd=1.635u as=0.341p ps=2.43u w=0.775u l=0.6u
X3410 VPWR.t5983 a_66204_3160# a_66116_3204# VPWR.t5244 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3411 _402_.B _324_.C.t20 VPWR.t6801 VPWR.t6800 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3412 VPWR.t5292 a_63404_23111# a_63316_23208# VPWR.t5291 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3413 VPWR.t5 a_59332_29816# _267_.A2 VPWR.t4 pfet_06v0 ad=0.4268p pd=2.175u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3414 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN VGND.t1313 VGND.t1312 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3415 a_33500_19975# a_33412_20072# VGND.t5874 VGND.t3592 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3416 a_50724_24908# _381_.A2.t4 a_50464_24908# VPWR.t6981 pfet_06v0 ad=0.1736p pd=1.18u as=0.224p ps=1.36u w=0.56u l=0.5u
X3417 a_44476_15704# a_44388_15748# VGND.t5876 VGND.t5875 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3418 VGND.t1141 _290_.ZN uo_out[5].t2 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X3419 a_67861_30644# a_67741_30600# a_67117_30600# VGND.t45 nfet_06v0 ad=43.2f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3420 _379_.Z uio_out[7].t11 a_18472_29076# VGND.t6584 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3421 VPWR.t3177 a_59932_11000# a_59844_11044# VPWR.t3176 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3422 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t1049 VPWR.t1048 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3423 VGND.t4458 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN VGND.t4457 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3424 _475_.D _421_.A1 a_47271_21640# VPWR pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X3425 _370_.B _334_.A1 a_32240_31048# VPWR.t2356 pfet_06v0 ad=0.3159p pd=1.735u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3426 a_47612_14136# a_47524_14180# VGND.t1541 VGND.t1540 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3427 VPWR.t5733 a_1468_15271# a_1380_15368# VPWR.t1241 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3428 _390_.ZN _395_.A2 VGND.t5623 VGND.t5622 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X3429 VPWR.t6839 clk.t7 a_44296_24393.t7 VPWR.t6838 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X3430 a_1468_3160# a_1380_3204# VGND.t3021 VGND.t501 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3431 a_10204_1592# a_10116_1636# VGND.t3365 VGND.t3364 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3432 a_40444_1159# a_40356_1256# VGND.t3367 VGND.t3366 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3433 _230_.I.t0 a_61860_30736# VPWR.t5653 VPWR.t5652 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X3434 a_56796_9432# a_56708_9476# VGND.t3369 VGND.t3368 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3435 a_47612_11000# a_47524_11044# VGND.t4369 VGND.t1524 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3436 VPWR.t3524 a_67996_6296# a_67908_6340# VPWR.t3523 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3437 VPWR.t3526 a_7068_1159# a_6980_1256# VPWR.t3525 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3438 VPWR.t5708 a_27172_24328# _352_.ZN VPWR.t5707 pfet_06v0 ad=0.34437p pd=1.895u as=0.31207p ps=1.665u w=1.095u l=0.5u
X3439 a_16588_20408# a_16500_20452# VGND.t1006 VGND.t1005 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3440 VPWR.t4230 a_67996_3160# a_67908_3204# VPWR.t1432 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3441 _335_.ZN.t14 _362_.B.t12 VPWR.t6534 VPWR.t6533 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3442 _474_.CLK.t16 a_48272_25156.t30 VPWR.t6561 VPWR.t6560 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3443 VPWR.t3233 a_2812_18840# a_2724_18884# VPWR.t365 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3444 a_43003_28409# a_41028_28776.t5 a_42368_28733# VPWR.t7098 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X3445 VPWR.t1660 a_24652_30951# a_24564_31048# VPWR.t1659 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3446 a_67548_7864# a_67460_7908# VGND.t3079 VGND.t3078 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3447 VPWR.t1568 a_2812_15704# a_2724_15748# VPWR.t1567 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3448 VPWR.t2446 a_13452_30951# a_13364_31048# VPWR.t2445 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3449 a_18028_28777# _378_.ZN a_17860_28777# VGND.t3302 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X3450 VPWR.t5346 a_2812_7431# a_2724_7528# VPWR.t5345 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3451 vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t1317 VPWR.t1316 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3452 a_46316_29977# a_45800_30345# VPWR.t5258 VPWR.t5257 pfet_06v0 ad=43.2f pd=0.6u as=0.1044p ps=0.94u w=0.36u l=0.5u
X3453 VPWR.t3487 a_31932_2727# a_31844_2824# VPWR.t3486 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3454 a_67548_4728# a_67460_4772# VGND.t4588 VGND.t4290 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3455 a_25008_25597# a_24636_25641# VGND.t4590 VGND.t4589 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X3456 a_11996_1592# a_11908_1636# VGND.t4592 VGND.t4591 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3457 a_49852_1159# a_49764_1256# VGND.t4594 VGND.t4593 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3458 VPWR.t4693 _304_.B a_50176_26724# VPWR.t4692 pfet_06v0 ad=0.389p pd=2.02u as=0.224p ps=1.36u w=0.56u l=0.5u
X3459 a_33612_24679# a_33524_24776# VGND.t4596 VGND.t4595 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3460 a_26668_21976# a_26580_22020# VGND.t413 VGND.t412 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3461 VPWR.t4749 a_16588_21976# a_16500_22020# VPWR.t893 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3462 a_35964_1592# a_35876_1636# VGND.t4599 VGND.t4598 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3463 VPWR.t4471 a_7964_29383# a_7876_29480# VPWR.t4470 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3464 VGND.t4326 _311_.Z _313_.ZN VGND.t4325 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3465 VPWR.t2955 _352_.ZN a_26746_26344# VPWR.t2954 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X3466 a_59932_1592# a_59844_1636# VGND.t4328 VGND.t4327 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3467 a_35616_24776# a_35204_24455.t3 VPWR.t6397 VPWR.t6396 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3468 VGND.t6419 _324_.B.t28 _399_.ZN VGND.t6418 nfet_06v0 ad=0.23975p pd=1.475u as=0.1469p ps=1.085u w=0.565u l=0.6u
X3469 VPWR.t3759 a_25660_2727# a_25572_2824# VPWR.t3758 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3470 a_44364_16839# a_44276_16936# VGND.t4330 VGND.t4329 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3471 VPWR.t3761 a_49292_16839# a_49204_16936# VPWR.t3760 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3472 VPWR.t4480 vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I VPWR.t4479 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3473 VPWR.t3763 a_57468_16839# a_57380_16936# VPWR.t3762 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3474 VPWR.t3370 a_16140_24679# a_16052_24776# VPWR.t3369 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3475 VPWR.t3433 a_64860_7864# a_64772_7908# VPWR.t3432 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3476 a_18604_20408# a_18516_20452# VGND.t1391 VGND.t1390 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3477 _284_.ZN.t17 _284_.B VPWR.t5593 VPWR.t5592 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X3478 VPWR.t2430 a_62956_13703# a_62868_13800# VPWR.t2429 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3479 a_54420_21976# a_54824_22045# a_54768_22137# VPWR.t3944 pfet_06v0 ad=0.1665p pd=1.285u as=50.4f ps=0.64u w=0.36u l=0.5u
X3480 a_68108_13703# a_68020_13800# VGND.t5000 VGND.t4999 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3481 VPWR.t5165 a_55004_21543# a_54916_21640# VPWR.t5164 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3482 VPWR.t6226 a_12444_1159# a_12356_1256# VPWR.t549 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3483 _330_.ZN _330_.A1.t14 VGND.t215 VGND.t214 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X3484 a_45036_28248# a_44948_28292# VGND.t5436 VGND.t5435 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3485 a_65420_10567# a_65332_10664# VGND.t5004 VGND.t5003 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3486 VPWR.t2919 a_46156_25112# a_46068_25156# VPWR.t2918 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3487 a_2364_10567# a_2276_10664# VGND.t4486 VGND.t3845 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3488 a_35818_29860# _460_.Q _288_.ZN.t0 VPWR.t3481 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3489 VGND.t2915 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I VGND.t2914 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3490 a_54220_10567# a_54132_10664# VGND.t4488 VGND.t4487 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3491 a_11772_1159# a_11684_1256# VGND.t4410 VGND.t4409 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3492 a_54444_18407# a_54356_18504# VGND.t4490 VGND.t4489 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3493 VPWR.t4648 a_29804_21976# a_29716_22020# VPWR.t4647 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3494 VPWR.t1830 a_45372_9432# a_45284_9476# VPWR.t1829 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3495 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN VPWR.t1726 VPWR.t1725 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3496 a_24988_24679# a_24900_24776# VGND.t4165 VGND.t4164 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3497 a_62844_14136# a_62756_14180# VGND.t5432 VGND.t5431 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3498 VPWR.t1967 a_34844_15704# a_34756_15748# VPWR.t1966 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3499 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t2482 VPWR.t2481 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3500 a_24988_21543# a_24900_21640# VGND.t4167 VGND.t4166 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3501 a_58140_26680# a_58052_26724# VGND.t4169 VGND.t4168 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3502 a_63616_31128# ui_in[0].t1 VPWR.t7053 VPWR.t7052 pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X3503 a_50076_17272# a_49988_17316# VGND.t4171 VGND.t4170 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3504 a_62844_11000# a_62756_11044# VGND.t785 VGND.t784 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3505 VPWR.t5290 a_4940_13703# a_4852_13800# VPWR.t5289 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3506 a_51644_14136# a_51556_14180# VGND.t4741 VGND.t4302 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3507 a_10876_2727# a_10788_2824# VGND.t4173 VGND.t4172 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3508 VPWR.t4216 a_21180_1592# a_21092_1636# VPWR.t4215 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3509 VPWR.t2201 a_65532_12568# a_65444_12612# VPWR.t2200 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3510 a_26556_23111# a_26468_23208# VGND.t5206 VGND.t5205 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3511 VPWR.t6922 a_42392_22825.t24 _452_.CLK.t10 VPWR.t6921 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3512 VPWR.t1534 a_35516_15271# a_35428_15368# VPWR.t1533 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3513 a_51644_11000# a_51556_11044# VGND.t5408 VGND.t5407 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3514 VPWR.t1291 a_1916_13703# a_1828_13800# VPWR.t1290 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3515 a_38876_15271# a_38788_15368# VGND.t5208 VGND.t5207 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3516 a_36148_21976# _301_.A1 a_36764_22512# VGND.t3202 nfet_06v0 ad=0.1672p pd=1.64u as=60.8f ps=0.7u w=0.38u l=0.6u
X3517 a_64188_27815# a_64100_27912# VGND.t5210 VGND.t5209 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3518 a_28124_30600# a_28124_30600# VPWR.t5387 VPWR.t5386 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3519 VPWR.t5284 a_65084_30951# a_64996_31048# VPWR.t5283 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3520 _350_.A2.t13 _371_.A1.t16 a_31516_28292# VPWR.t6511 pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X3521 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN VGND.t5495 VGND.t5494 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3522 a_28572_2727# a_28484_2824# VGND.t4177 VGND.t3052 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3523 VPWR.t4347 a_4604_4728# a_4516_4772# VPWR.t4346 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3524 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I VGND.t5689 VGND.t5688 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3525 a_3260_17272# a_3172_17316# VGND.t4180 VGND.t1722 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3526 VPWR.t3234 a_67548_7864# a_67460_7908# VPWR.t1401 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3527 a_38842_17316# _330_.A1.t15 _330_.ZN VPWR.t215 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3528 VPWR.t5758 a_28796_23111# a_28708_23208# VPWR.t5757 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3529 a_9308_1592# a_9220_1636# VGND.t4182 VGND.t4181 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3530 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I VGND.t5404 VGND.t5403 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3531 _362_.ZN _358_.A3 a_32628_26725# VPWR.t474 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3532 VPWR.t6011 a_4604_1592# a_4516_1636# VPWR.t6010 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3533 VPWR.t6009 a_27676_1592# a_27588_1636# VPWR.t5972 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3534 a_54420_21976# a_54864_22461.t5 a_54816_22505# VGND.t6311 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X3535 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t6246 VPWR.t6245 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3536 a_44252_1159# a_44164_1256# VGND.t4986 VGND.t4985 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3537 a_52764_1159# a_52676_1256# VGND.t1259 VGND.t1258 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3538 a_38772_28292# _437_.A1.t10 a_38584_28292# VPWR.t6861 pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X3539 a_50524_15704# a_50436_15748# VGND.t4988 VGND.t4987 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3540 a_43784_19369# a_43440_19325.t4 a_42996_18840# VPWR.t6463 pfet_06v0 ad=0.1791p pd=1.355u as=0.1665p ps=1.285u w=0.36u l=0.5u
X3541 a_30778_31048# _459_.Q.t11 _287_.A2 VPWR.t6972 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3542 VPWR.t4102 a_64636_1159# a_64548_1256# VPWR.t1097 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3543 a_61612_23111# a_61524_23208# VGND.t4990 VGND.t4989 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3544 VPWR.t1427 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN VPWR.t1426 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3545 a_63952_29480# _230_.I.t8 _250_.B VPWR.t6635 pfet_06v0 ad=0.5346p pd=3.31u as=0.37665p ps=1.835u w=1.215u l=0.5u
X3546 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I VGND.t3645 VGND.t3644 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3547 VPWR.t5156 _473_.Q _417_.A2.t1 VPWR.t5155 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3548 a_63952_29480# _251_.A1.t21 a_63336_29480# VPWR.t7016 pfet_06v0 ad=0.3402p pd=1.775u as=0.37665p ps=1.835u w=1.215u l=0.5u
X3549 VGND.t6364 _452_.CLK.t45 a_33748_20936.t1 VGND.t6363 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3550 _452_.CLK.t11 a_42392_22825.t25 VPWR.t6924 VPWR.t6923 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3551 VPWR.t1479 a_44160_29123# a_44132_29535# VPWR.t1478 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X3552 VGND.t1144 _248_.B1 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t1143 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3553 VPWR.t5476 _243_.B2 a_58656_27912# VPWR.t5475 pfet_06v0 ad=0.6588p pd=3.52u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3554 VPWR.t5373 a_23756_20408# a_23668_20452# VPWR.t5372 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3555 a_32580_27912# _287_.A1.t21 uo_out[6].t6 VPWR.t6784 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3556 a_54780_9432# a_54692_9476# VGND.t5202 VGND.t5201 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3557 a_37472_24419# a_37179_24831# VGND.t1590 VGND.t1589 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X3558 VPWR.t7106 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN VPWR.t7105 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3559 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I VGND.t5915 VGND.t5914 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3560 VPWR.t1265 _399_.ZN a_46580_23588# VPWR.t1264 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3561 VPWR.t1037 a_63852_23111# a_63764_23208# VPWR.t1036 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3562 a_49152_30301.t1 _474_.CLK.t42 VGND.t6455 VGND.t139 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3563 a_51532_12135# a_51444_12232# VGND.t4726 VGND.t4725 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3564 a_35740_25112# a_35652_25156# VGND.t4727 VGND.t1991 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3565 VPWR.t5178 a_2364_27815# a_2276_27912# VPWR.t2642 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3566 a_47612_10567# a_47524_10664# VGND.t4728 VGND.t1287 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3567 a_45564_21236# _324_.C.t21 _424_.A2.t4 VGND.t6509 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3568 VGND.t5791 a_19328_28733# a_19280_28777# VGND.t5790 nfet_06v0 ad=0.2333p pd=1.555u as=43.2f ps=0.6u w=0.36u l=0.6u
X3569 a_22352_25987# a_22059_26399# VPWR.t5836 VPWR.t5835 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X3570 VPWR.t3491 a_1468_23544# a_1380_23588# VPWR.t425 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3571 VPWR.t3193 a_19612_26247# a_19524_26344# VPWR.t3192 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3572 a_34256_24073# a_33376_23659# a_33932_24073# VGND.t1812 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X3573 a_46492_17272# a_46404_17316# VGND.t5249 VGND.t5248 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3574 a_48060_30951# a_47972_31048# VGND.t5250 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3575 a_6620_29383# a_6532_29480# VGND.t5252 VGND.t5251 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3576 a_23920_27555# a_23627_27967# VPWR.t2520 VPWR.t2519 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X3577 a_54768_22137# a_54040_22366# VPWR.t3254 VPWR.t3253 pfet_06v0 ad=50.4f pd=0.64u as=0.23p ps=1.54u w=0.36u l=0.5u
X3578 VPWR.t3922 a_19612_23111# a_19524_23208# VPWR.t3921 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3579 a_21516_25112# a_21428_25156# VGND.t5254 VGND.t5253 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3580 VPWR.t5436 a_22636_21976# a_22548_22020# VPWR.t5435 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3581 a_35292_17272# a_35204_17316# VGND.t4427 VGND.t4426 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3582 a_40464_27165# a_40092_27209# VPWR.t526 VPWR.t525 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X3583 VPWR.t3250 a_66540_16839# a_66452_16936# VPWR.t3249 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3584 VGND.t5055 _246_.B2 a_59620_27208# VGND.t5054 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3585 VGND.t3266 a_62564_29032# a_61940_29076# VGND.t3265 nfet_06v0 ad=0.218p pd=1.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3586 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN VGND.t3912 VGND.t3911 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3587 a_21516_21976# a_21428_22020# VGND.t5325 VGND.t5324 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3588 a_50412_16839# a_50324_16936# VGND.t4429 VGND.t4428 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3589 VGND.t588 a_42392_19243# _325_.A1.t3 VGND.t587 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3590 VPWR.t3027 a_50748_15271# a_50660_15368# VPWR.t3026 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3591 VPWR.t1608 a_2812_29383# a_2724_29480# VPWR.t1607 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3592 a_46268_12568# a_46180_12612# VGND.t4430 VGND.t381 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3593 VPWR.t30 _284_.A2.t4 a_45396_25156# VPWR.t29 pfet_06v0 ad=0.4818p pd=3.07u as=0.4599p ps=1.935u w=1.095u l=0.5u
X3594 a_30588_23111# a_30500_23208# VGND.t4787 VGND.t4786 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3595 VPWR.t329 a_1020_21543# a_932_21640# VPWR.t328 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3596 a_7964_1159# a_7876_1256# VGND.t5945 VGND.t5944 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3597 a_36284_29167# _462_.D a_36116_29167# VGND.t3410 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X3598 VPWR.t3029 a_2812_26247# a_2724_26344# VPWR.t3028 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3599 a_15580_1159# a_15492_1256# VGND.t4791 VGND.t4790 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3600 a_59036_11000# a_58948_11044# VGND.t4659 VGND.t4658 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3601 VPWR.t4941 a_62060_12135# a_61972_12232# VPWR.t4940 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3602 VPWR.t3100 a_2812_23111# a_2724_23208# VPWR.t3099 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3603 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN VPWR.t1516 VPWR.t1515 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3604 a_46940_15704# a_46852_15748# VGND.t4795 VGND.t4794 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3605 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN VGND.t2862 VGND.t2861 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3606 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t2908 VGND.t2907 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3607 a_35740_15704# a_35652_15748# VGND.t4915 VGND.t4914 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3608 VPWR.t2514 a_2364_18407# a_2276_18504# VPWR.t2513 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3609 clkbuf_1_0__f_clk.I.t27 a_44296_24393.t25 VGND.t275 VGND.t274 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X3610 a_56236_24679# a_56148_24776# VGND.t4916 VGND.t3237 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3611 VPWR.t5075 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN VPWR.t5074 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3612 a_4156_9432# a_4068_9476# VGND.t4921 VGND.t1641 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3613 VGND.t6574 _448_.Q.t7 a_43819_24372# VGND.t6573 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3614 a_64412_8999# a_64324_9096# VGND.t4922 VGND.t2232 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3615 a_53744_22851.t1 _474_.CLK.t43 VGND.t6457 VGND.t6456 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3616 a_24952_29032# _349_.A4 a_25340_29167# VGND.t2436 nfet_06v0 ad=0.1606p pd=1.61u as=58.39999f ps=0.685u w=0.365u l=0.6u
X3617 a_4156_6296# a_4068_6340# VGND.t5152 VGND.t730 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3618 VPWR.t6249 a_55452_21543# a_55364_21640# VPWR.t6248 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3619 VPWR.t2658 _274_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I VPWR.t2657 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3620 a_64412_5863# a_64324_5960# VGND.t5133 VGND.t2795 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3621 a_45156_21236# _324_.B.t29 VGND.t6421 VGND.t6420 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3622 VGND.t6275 a_48272_25156.t31 _474_.CLK.t17 VGND.t6274 nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3623 a_42908_1592# a_42820_1636# VGND.t5134 VGND.t4639 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3624 VPWR.t2228 a_24392_28248# _346_.A2 VPWR.t2227 pfet_06v0 ad=0.40575p pd=2.055u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3625 a_45484_28248# a_45396_28292# VGND.t4072 VGND.t4071 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3626 VGND.t6605 a_42392_22825.t26 _452_.CLK.t12 VGND.t6604 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3627 a_44924_15271# a_44836_15368# VGND.t5136 VGND.t5135 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3628 _336_.A1 a_29184_25597# VPWR.t4204 VPWR.t4203 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3629 a_21404_23111# a_21316_23208# VGND.t5138 VGND.t5137 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3630 a_16252_29383# a_16164_29480# VGND.t5235 VGND.t5234 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3631 VPWR.t2726 a_2812_9432# a_2724_9476# VPWR.t2725 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3632 a_2364_29816# a_2276_29860# VGND.t5236 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3633 VPWR.t4223 _470_.Q _411_.A2.t5 VPWR.t4222 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3634 VPWR.t5419 a_1020_12135# a_932_12232# VPWR.t4583 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3635 a_48060_1159# a_47972_1256# VGND.t5547 VGND.t5546 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3636 a_56572_1159# a_56484_1256# VGND.t4013 VGND.t4012 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3637 a_54892_18407# a_54804_18504# VGND.t5239 VGND.t5238 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3638 VPWR.t3732 a_42796_23981# hold2.Z VPWR.t3731 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3639 a_44282_24164# a_44162_24120# VGND.t4838 VGND.t4837 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3640 a_23084_28248# a_22996_28292# VGND.t492 VGND.t491 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3641 VPWR.t2122 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN VPWR.t2121 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3642 a_47860_21640# _421_.A1 _416_.A2 VPWR.t5996 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3643 VPWR.t2126 vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I VPWR.t2125 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3644 a_17932_25112# a_17844_25156# VGND.t2024 VGND.t2023 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3645 _436_.B a_41392_27165# VPWR.t820 VPWR.t819 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3646 VGND.t6313 a_54864_22461.t6 a_56236_22505# VGND.t6312 nfet_06v0 ad=0.1584p pd=1.6u as=43.2f ps=0.6u w=0.36u l=0.6u
X3647 VPWR.t532 a_55900_1592# a_55812_1636# VPWR.t531 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3648 a_22496_27967# a_22064_27912# VPWR.t3412 VPWR.t3411 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X3649 VPWR.t1917 a_12444_29383# a_12356_29480# VPWR.t1916 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3650 a_17932_21976# a_17844_22020# VGND.t3412 VGND.t3411 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3651 VPWR.t347 a_45372_10567# a_45284_10664# VPWR.t346 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3652 VGND.t2732 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN VGND.t2731 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3653 VGND.t277 a_44296_24393.t26 clkbuf_1_0__f_clk.I.t26 VGND.t276 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3654 a_48776_20204# _417_.A2.t8 VGND.t132 VGND.t131 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3655 _274_.ZN _268_.A1.t5 a_52756_29076# VGND.t6442 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3656 VPWR.t6889 _448_.Q.t8 _441_.A2 VPWR.t6888 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3657 VPWR.t4759 a_65980_12568# a_65892_12612# VPWR.t4758 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3658 VPWR.t2386 a_23644_23111# a_23556_23208# VPWR.t2385 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3659 VPWR.t1939 a_52316_9432# a_52228_9476# VPWR.t1938 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3660 VPWR.t2389 a_3260_8999# a_3172_9096# VPWR.t647 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3661 VPWR.t3935 a_35816_21192# _319_.A3 VPWR.t3934 pfet_06v0 ad=0.40575p pd=2.055u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3662 VPWR.t732 a_16140_23544# a_16052_23588# VPWR.t731 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3663 VPWR.t2847 a_35964_15271# a_35876_15368# VPWR.t2846 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3664 a_5052_20408# a_4964_20452# VGND.t3963 VGND.t3962 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3665 VPWR.t4311 a_64188_14136# a_64100_14180# VPWR.t4310 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3666 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN VGND.t2913 VGND.t2912 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3667 VPWR.t2167 _431_.A3 a_38852_25156# VPWR.t2166 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3668 uo_out[4].t5 _287_.A1.t22 VGND.t6484 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X3669 a_32604_16839# a_32516_16936# VGND.t4149 VGND.t4094 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3670 VGND.t1351 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN VGND.t1350 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3671 VPWR.t4855 a_32380_1159# a_32292_1256# VPWR.t574 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3672 a_2364_1159# a_2276_1256# VGND.t636 VGND.t635 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3673 VPWR.t1180 a_45708_16839# a_45620_16936# VPWR.t576 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3674 a_48272_25156.t5 clkbuf_1_0__f_clk.I.t46 VPWR.t256 VPWR.t255 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X3675 VPWR.t4857 a_64188_11000# a_64100_11044# VPWR.t4856 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3676 VPWR.t6134 a_33500_19975# a_33412_20072# VPWR.t6133 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3677 a_49068_20408# _475_.Q a_49856_20936# VGND.t4856 nfet_06v0 ad=0.1848p pd=1.72u as=67.2f ps=0.74u w=0.42u l=0.6u
X3678 VPWR.t1789 a_44786_24120# a_44906_23588# VPWR.t1788 pfet_06v0 ad=0.1116p pd=0.98u as=61.19999f ps=0.7u w=0.36u l=0.5u
X3679 a_36420_28776# _334_.A1 _335_.ZN.t4 VGND.t2243 nfet_06v0 ad=0.1312p pd=1.14u as=0.4161p ps=1.905u w=0.82u l=0.6u
X3680 a_1020_27815# a_932_27912# VGND.t4713 VGND.t4712 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3681 a_29856_29123# a_29563_29535# VPWR.t5052 VPWR.t5051 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X3682 _444_.D _311_.A2.t8 VGND.t6107 VGND.t6106 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3683 VGND.t182 _384_.A3.t14 _384_.ZN VGND.t181 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3684 a_2364_23544# a_2276_23588# VGND.t4760 VGND.t619 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3685 a_51220_22504# _474_.Q VGND.t4655 VGND.t4654 nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3686 VPWR.t2777 a_67548_17272# a_67460_17316# VPWR.t2776 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3687 uo_out[6].t2 _287_.A2 VGND.t1930 VGND.t1929 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X3688 a_50704_27912# _424_.B1.t11 _409_.ZN VPWR.t6618 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3689 a_52092_1592# a_52004_1636# VGND.t4762 VGND.t4761 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3690 VPWR.t4915 a_52428_12135# a_52340_12232# VPWR.t4914 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3691 a_50972_15704# a_50884_15748# VGND.t4766 VGND.t4765 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3692 VPWR.t4493 a_5052_21976# a_4964_22020# VPWR.t4492 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3693 VPWR.t1027 a_3708_10567# a_3620_10664# VPWR.t1026 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3694 VGND.t161 a_41088_17757.t5 a_41048_17341# VGND.t160 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3695 VPWR.t4953 a_60828_2727# a_60740_2824# VPWR.t4952 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3696 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t2280 VGND.t2279 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3697 VPWR.t4957 a_47612_18407# a_47524_18504# VPWR.t4956 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3698 VGND.t1966 a_38616_24328# _311_.A2.t1 VGND.t1965 nfet_06v0 ad=0.23405p pd=1.555u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3699 VPWR.t2294 a_18268_30951# a_18180_31048# VPWR.t2293 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3700 a_23196_29816# a_23108_29860# VGND.t4345 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3701 VPWR.t634 a_16588_27815# a_16500_27912# VPWR.t633 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3702 VPWR.t6115 a_1468_7431# a_1380_7528# VPWR.t6114 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3703 vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN VGND.t5030 VGND.t5029 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3704 a_51332_24372# _424_.A2.t10 _412_.ZN VGND.t186 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3705 _397_.A4 _402_.A1.t16 VPWR.t6727 VPWR.t6726 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3706 _358_.A3 a_30724_26020# VPWR.t1084 VPWR.t1083 pfet_06v0 ad=0.5346p pd=3.31u as=0.4268p ps=2.175u w=1.215u l=0.5u
X3707 a_54780_2727# a_54692_2824# VGND.t441 VGND.t440 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3708 a_5052_14136# a_4964_14180# VGND.t3320 VGND.t3319 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3709 a_43246_23610# a_43126_24119# VPWR.t3362 VPWR.t3361 pfet_06v0 ad=61.19999f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X3710 VPWR.t2699 a_1916_12568# a_1828_12612# VPWR.t2698 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3711 a_55208_22505# a_54824_22045# a_54420_21976# VGND.t3794 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3712 VPWR.t455 a_9532_1159# a_9444_1256# VPWR.t454 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3713 a_58588_1592# a_58500_1636# VGND.t445 VGND.t444 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3714 a_5052_11000# a_4964_11044# VGND.t4042 VGND.t4041 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3715 VPWR.t1780 a_53884_1592# a_53796_1636# VPWR.t1779 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3716 VPWR.t459 a_55004_14136# a_54916_14180# VPWR.t458 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3717 a_59397_26344# _251_.A1.t22 _252_.ZN VPWR.t7017 pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3718 a_51980_12135# a_51892_12232# VGND.t669 VGND.t668 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3719 VPWR.t6673 _355_.C.t11 a_20250_31048# VPWR.t6672 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X3720 VPWR.t678 a_65308_4295# a_65220_4392# VPWR.t677 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3721 VPWR.t933 a_28256_25597# a_28228_25273# VPWR.t932 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X3722 VPWR.t680 a_55004_11000# a_54916_11044# VPWR.t679 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3723 VGND.t453 a_36544_24419# a_36496_24463# VGND.t452 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X3724 VPWR.t2835 a_1468_30951# a_1380_31048# VPWR.t2834 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3725 _450_.D _327_.Z VGND.t5367 VGND.t5366 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X3726 VPWR.t901 a_62844_27815# a_62756_27912# VPWR.t900 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3727 a_50188_13703# a_50100_13800# VGND.t675 VGND.t674 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3728 a_58364_25112# a_58276_25156# VGND.t677 VGND.t676 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3729 VPWR.t2149 a_24196_31048# a_24196_31048# VPWR.t2148 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3730 VPWR.t339 a_15244_21543# a_15156_21640# VPWR.t338 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3731 a_41228_27815# a_41140_27912# VGND.t5306 VGND.t5305 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3732 a_21964_25112# a_21876_25156# VGND.t5308 VGND.t5307 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3733 VPWR.t5500 a_59036_1159# a_58948_1256# VPWR.t762 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3734 a_21964_21976# a_21876_22020# VGND.t1636 VGND.t1635 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3735 a_7964_2727# a_7876_2824# VGND.t5312 VGND.t5311 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3736 a_50860_16839# a_50772_16936# VGND.t5314 VGND.t5313 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3737 VPWR.t2948 a_31372_23544# a_31284_23588# VPWR.t2947 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3738 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I _274_.A1 VGND.t2519 VGND.t2518 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3739 VPWR.t5506 a_66652_6296# a_66564_6340# VPWR.t5505 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3740 VPWR.t164 a_41088_17757.t6 a_41048_17341# VPWR.t163 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3741 VPWR.t6016 a_43888_19204# a_43784_19369# VPWR.t6015 pfet_06v0 ad=0.1044p pd=0.94u as=0.1791p ps=1.355u w=0.36u l=0.5u
X3742 VPWR.t4977 a_4156_24679# a_4068_24776# VPWR.t557 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3743 uo_out[5].t6 _287_.A1.t23 VGND.t6485 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X3744 a_4940_7431# a_4852_7528# VGND.t5140 VGND.t5139 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3745 _436_.ZN _433_.ZN a_40565_24394# VGND.t568 nfet_06v0 ad=0.21175p pd=1.41u as=85.2f ps=0.95u w=0.71u l=0.6u
X3746 VPWR.t1506 a_20172_23544# a_20084_23588# VPWR.t1505 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3747 a_53212_29816# _268_.A1.t6 a_54000_30344# VGND.t3612 nfet_06v0 ad=0.1848p pd=1.72u as=67.2f ps=0.74u w=0.42u l=0.6u
X3748 VPWR.t5316 a_62060_20408# a_61972_20452# VPWR.t5315 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3749 VPWR.t2510 a_66652_3160# a_66564_3204# VPWR.t2509 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3750 a_23084_30951# a_22996_31048# VGND.t5143 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3751 a_59484_11000# a_59396_11044# VGND.t3994 VGND.t3993 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3752 VPWR.t5418 a_2364_29816# a_2276_29860# VPWR.t2663 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3753 a_49180_9432# a_49092_9476# VGND.t5145 VGND.t5144 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3754 VPWR.t26 a_53744_22851.t5 a_53704_23219# VPWR.t25 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3755 _452_.D _330_.A1.t16 VGND.t217 VGND.t216 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3756 _231_.ZN _231_.I VGND.t5903 VGND.t5902 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3757 a_2812_4295# a_2724_4392# VGND.t4201 VGND.t4200 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3758 a_63404_13703# a_63316_13800# VGND.t4203 VGND.t4202 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3759 VPWR.t4370 a_2364_26680# a_2276_26724# VPWR.t4369 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3760 a_66204_7864# a_66116_7908# VGND.t4206 VGND.t863 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3761 a_57468_2727# a_57380_2824# VGND.t4208 VGND.t4207 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3762 a_66204_4728# a_66116_4772# VGND.t1257 VGND.t833 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3763 a_10652_1592# a_10564_1636# VGND.t4210 VGND.t4209 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3764 a_3708_19975# a_3620_20072# VGND.t4128 VGND.t4127 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3765 _434_.ZN _304_.A1.t9 VPWR.t6605 VPWR.t6604 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3766 a_4156_2727# a_4068_2824# VGND.t4130 VGND.t4129 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3767 a_34620_1592# a_34532_1636# VGND.t4132 VGND.t4131 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3768 _302_.Z a_38576_22504# VGND.t5606 VGND.t5605 nfet_06v0 ad=0.3586p pd=2.51u as=0.226p ps=1.515u w=0.815u l=0.6u
X3769 _342_.ZN _343_.A2 VGND.t1183 VGND.t1182 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X3770 a_59932_12568# a_59844_12612# VGND.t4134 VGND.t4133 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3771 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I VPWR.t1602 VPWR.t1601 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3772 VPWR.t4299 a_63516_18840# a_63428_18884# VPWR.t1989 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3773 a_40244_18180# _452_.Q.t11 VPWR.t6956 VPWR.t6955 pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X3774 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN VGND.t3282 VGND.t3281 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3775 a_50420_23233# _395_.A1 _399_.A1 VPWR.t907 pfet_06v0 ad=0.58035p pd=2.155u as=0.4012p ps=1.85u w=1.095u l=0.5u
X3776 VGND.t1956 a_34080_22461# a_34032_22505# VGND.t1955 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X3777 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t1319 VPWR.t1318 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3778 VPWR.t2572 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN VPWR.t2571 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3779 a_6172_1159# a_6084_1256# VGND.t5935 VGND.t5934 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3780 VPWR.t5259 a_63516_15704# a_63428_15748# VPWR.t1611 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3781 VPWR.t6198 a_2812_28248# a_2724_28292# VPWR.t2822 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3782 VPWR.t6405 _337_.A3.t9 _371_.A2 VPWR.t6404 pfet_06v0 ad=0.4056p pd=1.805u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3783 VGND.t6607 a_42392_22825.t27 _452_.CLK.t13 VGND.t6606 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3784 a_25100_30951# a_25012_31048# VGND.t5937 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3785 a_67996_7864# a_67908_7908# VGND.t5939 VGND.t5938 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3786 a_31708_17272# a_31620_17316# VGND.t5940 VGND.t5649 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3787 VPWR.t3995 a_1020_20408# a_932_20452# VPWR.t3540 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3788 VPWR.t6232 a_4156_15271# a_4068_15368# VPWR.t2117 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3789 VPWR.t1481 a_52316_15704# a_52228_15748# VPWR.t1480 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3790 a_21852_23111# a_21764_23208# VGND.t3842 VGND.t3841 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3791 a_54000_30344# _268_.A2.t2 a_53796_30344# VGND.t3612 nfet_06v0 ad=67.2f pd=0.74u as=88.2f ps=0.84u w=0.42u l=0.6u
X3792 VPWR.t6999 _335_.ZN.t23 _350_.A2.t17 VPWR.t6998 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3793 VPWR.t1359 a_2812_25112# a_2724_25156# VPWR.t1358 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3794 VPWR.t5004 _475_.Q a_47524_22021# VPWR.t5003 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3795 VGND.t6725 _397_.A2.t10 _386_.ZN VGND.t6724 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3796 VPWR.t2131 a_30812_15271# a_30724_15368# VPWR.t1543 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3797 VPWR.t4106 a_44340_26183# a_43736_25896# VPWR.t4105 pfet_06v0 ad=0.23p pd=1.54u as=0.352p ps=2.48u w=0.8u l=0.5u
X3798 a_67996_4728# a_67908_4772# VGND.t3492 VGND.t3491 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3799 VPWR.t6477 _459_.CLK.t31 a_21652_27591.t0 VPWR.t6476 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3800 a_59372_12135# a_59284_12232# VGND.t3844 VGND.t3843 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3801 a_56348_15271# a_56260_15368# VGND.t5296 VGND.t1065 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3802 VPWR.t5549 a_46716_30951# a_46628_31048# VPWR.t5548 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3803 VPWR.t1219 a_12892_29383# a_12804_29480# VPWR.t1218 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3804 a_36960_27912# a_36548_27591.t3 VPWR.t6614 VPWR.t6613 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3805 VPWR.t6064 vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t6063 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3806 VPWR.t6309 a_2364_17272# a_2276_17316# VPWR.t5711 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3807 VPWR.t304 _424_.A1 _395_.A3 VPWR.t303 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3808 VPWR.t5493 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN VPWR.t5492 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3809 VGND.t279 a_44296_24393.t27 clkbuf_1_0__f_clk.I.t25 VGND.t278 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3810 VPWR.t4495 a_23196_29816# a_23108_29860# VPWR.t4494 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3811 VGND.t4496 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN VGND.t4495 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3812 VPWR.t6822 _325_.A1.t12 _226_.ZN VPWR.t6821 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3813 a_40416_18885# _327_.Z _331_.ZN VPWR.t5571 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3814 a_15244_27815# a_15156_27912# VGND.t4476 VGND.t2341 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3815 _251_.A1.t4 a_63616_31128# VGND.t5881 VGND.t5880 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X3816 _275_.A2 _268_.A2.t3 VGND.t6745 VGND.t6744 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X3817 a_34304_24029# a_33932_24073# VGND.t530 VGND.t529 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X3818 a_16588_23544# a_16500_23588# VGND.t4477 VGND.t1165 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3819 VPWR.t6974 _459_.Q.t12 _335_.ZN.t17 VPWR.t6973 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3820 _352_.ZN _352_.A2.t25 a_26548_24372# VGND.t6670 nfet_06v0 ad=0.4161p pd=1.905u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3821 VPWR.t2882 a_12892_1159# a_12804_1256# VPWR.t1551 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3822 VGND.t2179 a_53300_23047# a_52920_22760# VGND.t2178 nfet_06v0 ad=0.142p pd=1.14u as=0.176p ps=1.68u w=0.4u l=0.6u
X3823 a_29356_21976# a_29268_22020# VGND.t5363 VGND.t5362 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3824 VPWR.t4633 a_19276_21976# a_19188_22020# VPWR.t4632 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3825 a_24636_25641# _457_.D a_24512_25273# VPWR.t2956 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X3826 a_52988_26680# a_52900_26724# VGND.t4835 VGND.t4834 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3827 VGND.t1349 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN VGND.t1348 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3828 a_58252_16839# a_58164_16936# VGND.t4481 VGND.t4480 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3829 a_50197_28776# _392_.A2 VGND.t4193 VGND.t4192 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3830 a_59820_13703# a_59732_13800# VGND.t4615 VGND.t4614 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3831 a_63292_1159# a_63204_1256# VGND.t4617 VGND.t4616 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3832 VPWR.t4773 a_1020_14136# a_932_14180# VPWR.t2109 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3833 _417_.A2.t2 _473_.Q a_46389_21236# VGND.t4996 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3834 a_56388_25940# vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I VGND.t4284 VGND.t4283 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3835 VPWR.t6332 _288_.ZN.t6 a_37844_29860# VPWR.t6331 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3836 a_54332_20408# a_54244_20452# VGND.t3257 VGND.t3256 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3837 VGND.t1656 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I VGND.t1655 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3838 a_37308_1592# a_37220_1636# VGND.t4620 VGND.t4619 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3839 a_47052_16839# a_46964_16936# VGND.t4622 VGND.t4621 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3840 a_19948_26680# a_19860_26724# VGND.t1095 VGND.t350 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3841 VPWR.t5543 a_47388_15271# a_47300_15368# VPWR.t1559 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3842 VGND.t4653 _474_.Q a_48776_20204# VGND.t4652 nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3843 a_52756_29076# _268_.A2.t4 _274_.ZN VGND.t6746 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3844 a_60276_29032# _238_.I VGND.t2133 VGND.t2132 nfet_06v0 ad=0.176p pd=1.68u as=0.104p ps=0.92u w=0.4u l=0.6u
X3845 VPWR.t4520 a_1020_11000# a_932_11044# VPWR.t3594 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3846 a_21600_26725# _346_.ZN VPWR.t4522 VPWR.t4521 pfet_06v0 ad=0.44955p pd=1.955u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3847 uo_out[6].t10 _287_.A1.t24 VGND.t6487 VGND.t6486 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X3848 a_61500_27815# a_61412_27912# VGND.t4377 VGND.t4376 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3849 VPWR.t4934 a_67996_17272# a_67908_17316# VPWR.t4933 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3850 VPWR.t4947 a_27004_2727# a_26916_2824# VPWR.t4946 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3851 VPWR.t4526 a_52876_12135# a_52788_12232# VPWR.t4525 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3852 a_52352_26031# a_51576_25896# VGND.t2158 VGND.t2157 nfet_06v0 ad=43.2f pd=0.6u as=0.142p ps=1.14u w=0.36u l=0.6u
X3853 VPWR.t4371 a_66204_7864# a_66116_7908# VPWR.t1615 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3854 a_3260_1592# a_3172_1636# VGND.t4734 VGND.t1171 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3855 VPWR.t5746 a_26332_1592# a_26244_1636# VPWR.t5745 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3856 VPWR.t4887 a_30028_20408# a_29940_20452# VPWR.t4886 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3857 a_51332_24072# _384_.A3.t15 _427_.A2 VGND.t183 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3858 a_29804_23544# a_29716_23588# VGND.t4738 VGND.t4737 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3859 a_62620_19975# a_62532_20072# VGND.t4740 VGND.t4739 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3860 VPWR.t4691 _304_.B _435_.A3 VPWR.t4690 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3861 VPWR.t6853 _455_.Q.t8 _371_.A2 VPWR.t6852 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3862 _437_.A1.t1 a_38816_27555# VGND.t5593 VGND.t5592 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3863 a_48321_23208# _399_.A2 _399_.ZN VPWR.t1473 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3864 a_44786_24120# hold2.I VPWR.t2542 VPWR.t2541 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3865 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I VPWR.t3073 VPWR.t3072 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3866 a_56828_25940# _251_.A1.t23 a_56516_26344# VGND.t6696 nfet_06v0 ad=98.39999f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3867 a_30160_30301# a_29788_30345# VGND.t1841 VGND.t137 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X3868 a_53592_30344# _267_.A2 VGND.t3613 VGND.t3612 nfet_06v0 ad=88.2f pd=0.84u as=0.226p ps=1.515u w=0.42u l=0.6u
X3869 a_57132_18407# a_57044_18504# VGND.t5153 VGND.t3648 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3870 VPWR.t3394 a_34396_17272# a_34308_17316# VPWR.t3393 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3871 a_65308_18407# a_65220_18504# VGND.t5154 VGND.t3967 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3872 VPWR.t5327 a_62508_21976# a_62420_22020# VPWR.t5326 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3873 a_42587_25940# _324_.C.t22 _265_.ZN VGND.t6510 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3874 a_38506_26724# _437_.A1.t11 _443_.D VPWR.t6862 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3875 VPWR.t5554 a_48732_15704# a_48644_15748# VPWR.t4852 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3876 a_40220_19975# a_40132_20072# VGND.t5157 VGND.t5156 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3877 a_35552_27216# _358_.A3 VGND.t472 VGND.t471 nfet_06v0 ad=79.8f pd=0.8u as=0.2424p ps=1.635u w=0.38u l=0.6u
X3878 VPWR.t5330 a_57020_1159# a_56932_1256# VPWR.t5329 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3879 a_65532_14136# a_65444_14180# VGND.t3617 VGND.t3616 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3880 VPWR.t1650 a_37532_15704# a_37444_15748# VPWR.t1649 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3881 VPWR.t6112 a_5724_2727# a_5636_2824# VPWR.t6111 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3882 VPWR.t4919 a_55452_14136# a_55364_14180# VPWR.t4918 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3883 VGND.t324 _258_.I _258_.ZN VGND.t323 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3884 _261_.ZN _301_.A1 a_40004_22020# VPWR.t3349 pfet_06v0 ad=0.4016p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3885 VPWR.t6202 a_67996_7864# a_67908_7908# VPWR.t6201 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3886 a_65532_11000# a_65444_11044# VGND.t3799 VGND.t3798 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3887 VPWR.t4921 a_55452_11000# a_55364_11044# VPWR.t4920 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3888 a_9756_1592# a_9668_1636# VGND.t4773 VGND.t4772 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3889 a_54624_22895# a_54088_22895# VGND.t2800 VGND.t2799 nfet_06v0 ad=43.2f pd=0.6u as=0.2637p ps=1.825u w=0.36u l=0.6u
X3890 a_48988_26369# _397_.A1.t8 _284_.B VPWR.t16 pfet_06v0 ad=0.33945p pd=1.715u as=0.2847p ps=1.615u w=1.095u l=0.5u
X3891 a_62148_29505# _230_.I.t9 VPWR.t6637 VPWR.t6636 pfet_06v0 ad=0.55297p pd=2.105u as=0.4818p ps=3.07u w=1.095u l=0.5u
X3892 a_29244_23111# a_29156_23208# VGND.t4381 VGND.t4380 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3893 vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN VGND.t5414 VGND.t5413 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3894 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN VGND.t5873 VGND.t5872 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3895 VPWR.t5547 a_15692_21543# a_15604_21640# VPWR.t5546 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3896 a_39924_27209# a_39124_27208.t5 VGND.t228 VGND.t227 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3897 a_34084_28776# _460_.Q a_34700_28776# VGND.t3332 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3898 a_2364_7431# a_2276_7528# VGND.t4386 VGND.t3755 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3899 VPWR.t4534 a_39548_1159# a_39460_1256# VPWR.t2103 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3900 a_31484_2727# a_31396_2824# VGND.t4390 VGND.t4389 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3901 a_55788_25112# a_55700_25156# VGND.t4392 VGND.t4391 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3902 VPWR.t4355 a_1468_9432# a_1380_9476# VPWR.t2564 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3903 VPWR.t1772 a_60828_1592# a_60740_1636# VPWR.t1771 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3904 a_64220_29098# _249_.A2 VGND.t1465 VGND.t1464 nfet_06v0 ad=85.2f pd=0.95u as=0.22595p ps=1.45u w=0.71u l=0.6u
X3905 a_23920_27555# a_23627_27967# VGND.t2393 VGND.t2392 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X3906 a_43156_20452# _304_.A1.t10 _304_.ZN.t4 VPWR.t6606 pfet_06v0 ad=0.33945p pd=1.715u as=0.2847p ps=1.615u w=1.095u l=0.5u
X3907 a_4604_3160# a_4516_3204# VGND.t4214 VGND.t4213 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3908 VPWR.t5199 a_55228_2727# a_55140_2824# VPWR.t5198 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3909 VPWR.t3004 a_48384_26724# clkload0.Z VPWR.t3003 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3910 a_50032_30345# a_49496_30345# VGND.t860 VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=0.2637p ps=1.825u w=0.36u l=0.6u
X3911 a_59932_9432# a_59844_9476# VGND.t4216 VGND.t4215 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3912 a_44948_25156# _284_.A2.t5 VPWR.t32 VPWR.t31 pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X3913 a_64412_15704# a_64324_15748# VGND.t4218 VGND.t4217 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3914 VPWR.t1536 a_65196_23544# a_65108_23588# VPWR.t1535 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3915 a_53212_15704# a_53124_15748# VGND.t4220 VGND.t4219 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3916 a_53212_29816# _268_.A2.t5 VPWR.t7063 VPWR.t7062 pfet_06v0 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X3917 a_54088_22895# a_53704_23219# a_53300_23047# VGND.t3828 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3918 VPWR.t258 clkbuf_1_0__f_clk.I.t47 a_42392_22825.t3 VPWR.t257 pfet_06v0 ad=0.3608p pd=2.52u as=0.2542p ps=1.44u w=0.82u l=0.5u
X3919 VPWR.t4843 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN VPWR.t4842 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3920 a_64300_23111# a_64212_23208# VGND.t4695 VGND.t4694 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3921 a_41188_18840# _325_.A1.t13 a_41804_19376# VGND.t6518 nfet_06v0 ad=0.1672p pd=1.64u as=60.8f ps=0.7u w=0.38u l=0.6u
X3922 a_62284_16839# a_62196_16936# VGND.t4697 VGND.t4696 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3923 a_37744_20452# _317_.A2 VPWR.t2576 VPWR.t2575 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3924 a_63852_13703# a_63764_13800# VGND.t4699 VGND.t4698 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3925 VPWR.t6012 a_61276_1159# a_61188_1256# VPWR.t2099 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3926 a_40332_21543# a_40244_21640# VGND.t4701 VGND.t4700 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3927 VGND.t2517 _274_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I VGND.t2516 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3928 VPWR.t1592 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_56720_26344# VPWR.t1591 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X3929 VGND.t2242 _334_.A1 a_35216_27533# VGND.t2241 nfet_06v0 ad=0.218p pd=1.52u as=57.59999f ps=0.68u w=0.36u l=0.6u
X3930 a_2364_15271# a_2276_15368# VGND.t1040 VGND.t742 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3931 a_33764_27208# _460_.Q VGND.t3331 VGND.t3330 nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3932 VPWR.t1088 a_15244_20408# a_15156_20452# VPWR.t1087 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3933 a_65420_12135# a_65332_12232# VGND.t1044 VGND.t1043 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3934 a_8636_2727# a_8548_2824# VGND.t1046 VGND.t1045 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3935 a_50196_22805# _218_.ZN VGND.t3631 VGND.t3630 nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3936 a_56124_9432# a_56036_9476# VGND.t1048 VGND.t1047 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3937 a_2364_12135# a_2276_12232# VGND.t1050 VGND.t1049 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3938 _305_.A2 a_41488_24072# VPWR.t5629 VPWR.t5628 pfet_06v0 ad=0.5368p pd=3.32u as=0.395p ps=2.02u w=1.22u l=0.5u
X3939 _287_.A1.t3 a_38472_30169# VPWR.t4965 VPWR.t4964 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3940 a_43452_18191# _450_.D a_43328_18559# VPWR.t3852 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X3941 VPWR.t59 a_63964_18840# a_63876_18884# VPWR.t58 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3942 a_54220_12135# a_54132_12232# VGND.t52 VGND.t51 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3943 _495_.I _304_.B a_41708_30644# VGND.t34 nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3944 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN VPWR.t3067 VPWR.t3066 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3945 _416_.A2 _421_.A1 a_48068_21236# VGND.t5746 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3946 _378_.I _346_.B a_21287_29076# VGND.t401 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X3947 VPWR.t4484 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN VPWR.t4483 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3948 VGND.t3061 _378_.I _378_.ZN VGND.t3060 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3949 VPWR.t5878 a_63964_15704# a_63876_15748# VPWR.t5274 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3950 VPWR.t5879 a_4156_23544# a_4068_23588# VPWR.t1445 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3951 a_22636_23544# a_22548_23588# VGND.t54 VGND.t53 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3952 VPWR.t4065 a_66092_18407# a_66004_18504# VPWR.t4064 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3953 VPWR.t335 a_56516_26344# _242_.Z VPWR.t334 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X3954 a_49180_17272# a_49092_17316# VGND.t5160 VGND.t5159 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3955 a_36608_29167# a_35728_29480# a_36284_29167# VGND.t662 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X3956 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I VGND.t316 VGND.t315 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3957 VPWR.t5892 a_52764_15704# a_52676_15748# VPWR.t5891 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3958 a_29184_25597# a_28891_25273# VPWR.t463 VPWR.t462 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X3959 a_58924_14136# a_58836_14180# VGND.t5082 VGND.t5081 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3960 VPWR.t3684 a_41116_26247# a_41028_26344# VPWR.t3683 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3961 _390_.ZN _395_.A1 a_51968_26724# VPWR.t906 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X3962 VPWR.t4067 a_63068_18407# a_62980_18504# VPWR.t4066 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3963 VPWR.t5336 a_25324_21976# a_25236_22020# VPWR.t5335 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3964 VGND.t6658 _459_.Q.t13 a_34292_28776# VGND.t6657 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3965 a_41216_23208# _452_.Q.t12 a_41012_23208# VPWR.t6957 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3966 VGND.t4896 a_48708_29816# a_48104_30219# VGND.t2052 nfet_06v0 ad=0.142p pd=1.14u as=0.176p ps=1.68u w=0.4u l=0.6u
X3967 a_2812_13703# a_2724_13800# VGND.t4504 VGND.t2924 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3968 VGND.t3566 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I VGND.t3565 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3969 _360_.ZN _358_.A3 a_33188_25940# VGND.t470 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3970 VPWR.t3792 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t3791 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3971 VPWR.t4662 a_50300_20408# a_50212_20452# VPWR.t4661 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3972 a_53100_16839# a_53012_16936# VGND.t4508 VGND.t4507 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3973 a_60916_29612# _250_.ZN a_60656_29612# VPWR.t897 pfet_06v0 ad=0.1736p pd=1.18u as=0.224p ps=1.36u w=0.56u l=0.5u
X3974 VGND.t1193 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t1192 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3975 a_56796_15271# a_56708_15368# VGND.t4509 VGND.t1805 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3976 a_33276_23111# a_33188_23208# VGND.t4511 VGND.t4510 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3977 VPWR.t5570 _327_.Z a_39268_18840# VPWR.t5569 pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X3978 VPWR.t3648 a_42236_15271# a_42148_15368# VPWR.t423 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3979 VPWR.t4654 a_61052_12568# a_60964_12612# VPWR.t4653 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3980 a_64860_8999# a_64772_9096# VGND.t4600 VGND.t3288 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3981 a_15692_27815# a_15604_27912# VGND.t4602 VGND.t4601 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3982 a_53212_29816# _267_.A2 VPWR.t3751 VPWR.t3750 pfet_06v0 ad=0.156p pd=1.12u as=0.395p ps=2.02u w=0.6u l=0.5u
X3983 _373_.A2 _371_.ZN VGND.t5613 VGND.t102 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X3984 a_29020_1592# a_28932_1636# VGND.t4603 VGND.t595 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3985 VGND.t426 a_33520_25597# a_33472_25641# VGND.t425 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X3986 a_64860_5863# a_64772_5960# VGND.t4605 VGND.t4604 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3987 a_17904_28409# a_17472_28363# VPWR.t2639 VPWR.t2638 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X3988 a_54780_20408# a_54692_20452# VGND.t5373 VGND.t5372 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3989 _462_.D _359_.B.t8 a_36288_31048# VPWR.t6771 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X3990 a_41572_20072# _327_.Z VPWR.t5568 VPWR.t5567 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3991 a_37396_29860# _288_.ZN.t7 VPWR.t6334 VPWR.t6333 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3992 VPWR.t4540 a_61500_14136# a_61412_14180# VPWR.t4539 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3993 a_33724_21543# a_33636_21640# VGND.t4396 VGND.t4395 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3994 vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN VGND.t4257 VGND.t4256 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3995 _294_.ZN.t1 _223_.I a_32144_26724# VPWR.t7111 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X3996 VPWR.t4603 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].I VPWR.t4602 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3997 a_35516_28776# _459_.Q.t14 VGND.t6660 VGND.t6659 nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3998 VPWR.t3098 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN VPWR.t3097 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3999 VPWR.t4544 a_61500_11000# a_61412_11044# VPWR.t4543 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4000 VPWR.t4546 a_50300_14136# a_50212_14180# VPWR.t4545 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4001 vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN VGND.t4494 VGND.t4493 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4002 VPWR.t4547 a_43804_1159# a_43716_1256# VPWR.t2409 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4003 VPWR.t4501 a_30476_20408# a_30388_20452# VPWR.t4500 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4004 a_7740_1592# a_7652_1636# VGND.t4355 VGND.t4354 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4005 a_58116_30344# _270_.A2 _272_.A2 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4006 VPWR.t4505 a_50300_11000# a_50212_11044# VPWR.t4504 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4007 VPWR.t5413 _245_.I1 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t5412 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4008 VPWR.t260 clkbuf_1_0__f_clk.I.t48 a_48272_25156.t4 VPWR.t259 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X4009 _362_.B.t0 a_33776_29123# VPWR.t3534 VPWR.t3533 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4010 a_1468_4295# a_1380_4392# VGND.t502 VGND.t501 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4011 a_5052_29816# a_4964_29860# VGND.t4358 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4012 VGND.t6742 a_45456_30301.t2 a_45416_29885# VGND.t139 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X4013 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I VGND.t4362 VGND.t4361 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4014 a_47612_12135# a_47524_12232# VGND.t1525 VGND.t1524 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4015 a_36412_15271# a_36324_15368# VGND.t4775 VGND.t4774 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4016 a_57580_18407# a_57492_18504# VGND.t4776 VGND.t3239 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4017 _245_.Z a_61836_25515# VGND.t2466 VGND.t2465 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4018 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I VPWR.t7104 VPWR.t7103 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4019 VPWR.t5441 a_37532_1159# a_37444_1256# VPWR.t5440 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4020 a_49044_28292# _381_.Z a_48820_28292# VPWR.t3949 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4021 VGND.t6097 a_52400_25987.t4 a_52360_26355# VGND.t6096 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X4022 VPWR.t491 a_37532_26247# a_37444_26344# VPWR.t490 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4023 a_38644_19368# _451_.Q.t5 _330_.A2 VGND.t6148 nfet_06v0 ad=0.2132p pd=1.34u as=0.4161p ps=1.905u w=0.82u l=0.6u
X4024 a_32048_24463# a_29828_24455.t5 a_31803_24831# VGND.t6119 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4025 a_19388_1159# a_19300_1256# VGND.t4778 VGND.t4777 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4026 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN VGND.t1654 VGND.t1653 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4027 a_62508_10567# a_62420_10664# VGND.t4780 VGND.t4779 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4028 VGND.t6391 _355_.C.t12 _465_.D VGND.t102 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4029 a_65980_14136# a_65892_14180# VGND.t1687 VGND.t726 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4030 VPWR.t3739 a_53212_2727# a_53124_2824# VPWR.t3738 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4031 VPWR.t3768 a_37980_15704# a_37892_15748# VPWR.t3767 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4032 VPWR.t3502 a_15132_29383# a_15044_29480# VPWR.t3501 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4033 VPWR.t1834 a_38336_18147# a_38308_18559# VPWR.t1833 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X4034 a_33276_1592# a_33188_1636# VGND.t4136 VGND.t735 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4035 _250_.A2 _230_.I.t10 a_63105_28293# VPWR.t6638 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4036 VPWR.t4170 a_48060_10567# a_47972_10664# VPWR.t4169 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4037 a_35180_18407# a_35092_18504# VGND.t4138 VGND.t4137 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4038 _427_.B2 _281_.A1 VGND.t3146 VGND.t3145 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X4039 _261_.ZN _325_.A1.t14 VPWR.t6824 VPWR.t6823 pfet_06v0 ad=0.44325p pd=2.87u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4040 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I VPWR.t1683 VPWR.t1682 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4041 a_65980_11000# a_65892_11044# VGND.t5648 VGND.t5647 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4042 VPWR.t2476 a_49852_15271# a_49764_15368# VPWR.t2475 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4043 a_67548_8999# a_67460_9096# VGND.t4139 VGND.t3078 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4044 a_57244_1592# a_57156_1636# VGND.t4286 VGND.t4285 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4045 a_1916_20408# a_1828_20452# VGND.t1315 VGND.t1314 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4046 a_30672_24831# a_30240_24776# VPWR.t6318 VPWR.t6317 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X4047 VPWR.t3165 a_52540_1592# a_52452_1636# VPWR.t3164 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4048 a_27868_28776# _455_.Q.t9 a_25124_28776# VGND.t6537 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4049 a_29692_23111# a_29604_23208# VGND.t4288 VGND.t4287 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4050 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN VPWR.t5905 VPWR.t3734 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4051 a_32156_18407# a_32068_18504# VGND.t4289 VGND.t2770 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4052 VPWR.t3298 _281_.A1 _281_.ZN.t0 VPWR.t3297 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X4053 a_67548_5863# a_67460_5960# VGND.t4291 VGND.t4290 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4054 VPWR.t4293 a_3708_19975# a_3620_20072# VPWR.t3033 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4055 a_64188_12568# a_64100_12612# VGND.t4293 VGND.t4292 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4056 VGND.t2435 _349_.A4 a_26148_28776# VGND.t2434 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4057 VGND.t3018 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN VGND.t3017 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4058 VPWR.t282 a_44296_24393.t28 clkbuf_1_0__f_clk.I.t8 VPWR.t281 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4059 VGND.t540 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN _231_.I VGND.t539 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4060 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I VGND.t4282 VGND.t4281 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4061 a_59932_2727# a_59844_2824# VGND.t4468 VGND.t4327 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4062 a_67548_18840# a_67460_18884# VGND.t1185 VGND.t1184 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4063 VPWR.t5841 a_66316_12135# a_66228_12232# VPWR.t5840 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4064 a_64860_15704# a_64772_15748# VGND.t4470 VGND.t4469 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4065 a_48172_18840# a_48084_18884# VGND.t3233 VGND.t3232 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4066 a_5052_23544# a_4964_23588# VGND.t4472 VGND.t4471 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4067 VPWR.t6658 _452_.CLK.t46 a_33748_20936.t0 VPWR.t6657 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4068 vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN VGND.t2476 VGND.t2475 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4069 VPWR.t4629 a_1916_21976# a_1828_22020# VPWR.t3288 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4070 _284_.ZN.t15 _304_.B a_44028_25156# VPWR.t4689 pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
X4071 a_6620_2727# a_6532_2824# VGND.t4577 VGND.t4576 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4072 VPWR.t3276 a_29468_2727# a_29380_2824# VPWR.t3275 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4073 VPWR.t4735 a_9980_1159# a_9892_1256# VPWR.t4734 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4074 VPWR.t4352 a_55116_12135# a_55028_12232# VPWR.t4351 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4075 a_53660_15704# a_53572_15748# VGND.t4581 VGND.t4580 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4076 VPWR.t4158 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I VPWR.t4157 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4077 a_24392_28248# _343_.A2 VPWR.t1257 VPWR.t1256 pfet_06v0 ad=0.156p pd=1.12u as=0.40575p ps=2.055u w=0.6u l=0.5u
X4078 VPWR.t5993 a_65756_4295# a_65668_4392# VPWR.t997 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4079 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN VPWR.t903 VPWR.t902 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4080 VGND.t2274 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t2273 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4081 VPWR.t4738 a_41788_1159# a_41700_1256# VPWR.t4737 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4082 a_22064_27912# a_21652_27591.t6 VGND.t101 VGND.t100 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4083 VPWR.t5762 a_65756_1159# a_65668_1256# VPWR.t5761 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4084 a_40780_21543# a_40692_21640# VGND.t4109 VGND.t4108 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4085 a_1916_14136# a_1828_14180# VGND.t4154 VGND.t4153 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4086 a_31260_15704# a_31172_15748# VGND.t4111 VGND.t4110 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4087 a_56572_29383# a_56484_29480# VGND.t4113 VGND.t4112 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4088 a_37868_16839# a_37780_16936# VGND.t4115 VGND.t4114 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4089 a_59828_26724# _246_.B2 VPWR.t5213 VPWR.t5212 pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X4090 uio_out[6].t4 a_19328_28733# VGND.t5789 VGND.t5788 nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X4091 a_1916_11000# a_1828_11044# VGND.t1709 VGND.t1708 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4092 _441_.ZN _303_.ZN a_39780_22805# VGND.t2813 nfet_06v0 ad=0.4137p pd=1.9u as=0.2119p ps=1.335u w=0.815u l=0.6u
X4093 a_18816_29931# a_18404_30344.t5 VPWR.t139 VPWR.t138 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X4094 VPWR.t7102 a_4604_12568# a_4516_12612# VPWR.t7101 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4095 VPWR.t4277 a_15692_20408# a_15604_20452# VPWR.t4276 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4096 a_56124_2727# a_56036_2824# VGND.t4299 VGND.t4298 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4097 VPWR.t4068 a_1020_16839# a_932_16936# VPWR.t1061 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4098 VPWR.t4487 a_59484_1159# a_59396_1256# VPWR.t1065 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4099 a_55004_12568# a_54916_12612# VGND.t4301 VGND.t4300 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4100 VPWR.t7100 a_49068_20408# _419_.Z VPWR.t4798 pfet_06v0 ad=0.395p pd=2.02u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4101 VPWR.t1029 a_7180_30951# a_7092_31048# VPWR.t1028 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4102 VGND.t2357 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4103 a_51644_15271# a_51556_15368# VGND.t4303 VGND.t4302 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4104 VPWR.t6197 a_6172_1159# a_6084_1256# VPWR.t6196 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4105 VPWR.t2887 a_55228_1592# a_55140_1636# VPWR.t2685 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4106 VGND.t3101 a_54040_22366# _281_.A1 VGND.t3100 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4107 a_58924_10567# a_58836_10664# VGND.t4305 VGND.t4304 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4108 VPWR.t6117 a_4156_30951# a_4068_31048# VPWR.t6116 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4109 VPWR.t2162 a_45012_29816# a_44632_30206# VPWR.t2161 pfet_06v0 ad=0.23p pd=1.54u as=0.352p ps=2.48u w=0.8u l=0.5u
X4110 a_24960_25641# a_24080_25227# a_24636_25641# VGND.t4264 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X4111 VPWR.t7038 _397_.A2.t11 _395_.A1 VPWR.t7037 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4112 a_37516_27599# _443_.D a_37348_27599# VGND.t3879 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X4113 VPWR.t3721 a_4940_5863# a_4852_5960# VPWR.t3720 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4114 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN VGND.t4693 VGND.t4692 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4115 a_67436_19975# a_67348_20072# VGND.t4675 VGND.t4674 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4116 VPWR.t5093 a_41564_26247# a_41476_26344# VPWR.t5092 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4117 VPWR.t4826 a_25772_21976# a_25684_22020# VPWR.t4825 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4118 a_66652_7864# a_66564_7908# VGND.t4678 VGND.t577 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4119 VPWR.t3147 a_43132_27815# a_43044_27912# VPWR.t3146 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4120 _439_.ZN _325_.A1.t15 a_41440_23208# VPWR.t6825 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4121 a_56348_30951# a_56260_31048# VGND.t4679 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4122 VPWR.t135 _417_.A2.t9 a_51892_23340# VPWR.t134 pfet_06v0 ad=0.389p pd=2.02u as=0.1736p ps=1.18u w=0.56u l=0.5u
X4123 VGND.t6366 _452_.CLK.t47 a_32740_22504.t1 VGND.t6365 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X4124 a_33932_24073# _313_.ZN a_33764_24073# VGND.t1000 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X4125 VPWR.t324 _258_.I _258_.ZN VPWR.t323 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4126 VPWR.t2798 a_60268_10567# a_60180_10664# VPWR.t2797 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4127 a_66652_4728# a_66564_4772# VGND.t2472 VGND.t2471 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4128 VGND.t1311 vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN VGND.t1310 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4129 VPWR.t6425 _451_.Q.t6 a_41642_25156# VPWR.t6424 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X4130 a_45148_30951# a_45060_31048# VGND.t4123 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4131 a_3708_29383# a_3620_29480# VGND.t4124 VGND.t3501 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4132 VPWR.t4076 _270_.A2 a_58340_29860# VPWR.t4075 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4133 VPWR.t4891 a_62620_19975# a_62532_20072# VPWR.t4890 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4134 a_44500_22020# _304_.B _324_.B.t10 VPWR.t4688 pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X4135 VPWR.t5064 a_42684_15271# a_42596_15368# VPWR.t5030 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4136 _316_.A3 _301_.A1 a_37296_22020# VPWR.t3348 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X4137 a_62284_26680# a_62196_26724# VGND.t3005 VGND.t3004 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4138 VPWR.t5063 a_24952_29032# _343_.A2 VPWR.t5062 pfet_06v0 ad=0.40575p pd=2.055u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4139 VGND.t2121 a_24392_28248# _346_.A2 VGND.t2120 nfet_06v0 ad=0.23405p pd=1.555u as=0.3586p ps=2.51u w=0.815u l=0.6u
X4140 VPWR.t2383 a_63628_16839# a_63540_16936# VPWR.t2382 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4141 a_2364_28248# a_2276_28292# VGND.t2507 VGND.t1823 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4142 VPWR.t3203 a_22300_24679# a_22212_24776# VPWR.t3202 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4143 VPWR.t4507 a_5052_29816# a_4964_29860# VPWR.t4506 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4144 a_19248_29977# a_18816_29931# VPWR.t6098 VPWR.t6097 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X4145 VPWR.t5614 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN VPWR.t5613 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4146 VPWR.t2920 a_55340_25112# a_55252_25156# VPWR.t1609 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4147 VPWR.t4905 a_5052_26680# a_4964_26724# VPWR.t4904 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4148 VPWR.t5328 a_40220_19975# a_40132_20072# VPWR.t486 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4149 a_24736_26841# a_24304_26795# VPWR.t1157 VPWR.t1156 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X4150 VPWR.t3697 a_33052_16839# a_32964_16936# VPWR.t3696 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4151 a_50792_26344# a_50120_26476# VPWR.t2478 VPWR.t2477 pfet_06v0 ad=0.3172p pd=1.74u as=0.4005p ps=2.12u w=1.22u l=0.5u
X4152 VPWR.t524 _407_.A1 _407_.ZN VPWR.t523 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4153 VPWR.t1914 a_48508_12135# a_48420_12232# VPWR.t580 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4154 a_45128_26031# a_44784_25987.t5 a_44340_26183# VPWR.t178 pfet_06v0 ad=0.1791p pd=1.355u as=0.1665p ps=1.285u w=0.36u l=0.5u
X4155 a_36288_31048# _365_.ZN VPWR.t3560 VPWR.t3559 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4156 a_42084_24072# _260_.A1 a_41880_24072# VGND.t3773 nfet_06v0 ad=88.2f pd=0.84u as=88.2f ps=0.84u w=0.42u l=0.6u
X4157 a_58588_9432# a_58500_9476# VGND.t1988 VGND.t1987 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4158 VPWR.t5756 a_63068_17272# a_62980_17316# VPWR.t5755 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4159 VPWR.t1390 vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN VPWR.t1389 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4160 VPWR.t2090 a_66204_18840# a_66116_18884# VPWR.t2089 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4161 a_38131_22804# _448_.Q.t9 VGND.t6576 VGND.t6575 nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4162 a_35740_26247# a_35652_26344# VGND.t1992 VGND.t1991 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4163 _459_.D _358_.A2 VGND.t4689 VGND.t4688 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X4164 a_25792_30301# a_25420_30345# VGND.t5076 VGND.t137 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X4165 a_31260_1592# a_31172_1636# VGND.t1994 VGND.t1993 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4166 VPWR.t6156 a_55900_15271# a_55812_15368# VPWR.t6155 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4167 VGND.t6404 a_41048_29816.t13 _459_.CLK.t12 VGND.t6400 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4168 a_25740_28776# _349_.A4 VGND.t2433 VGND.t2432 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4169 a_47047_21640# _416_.A1.t8 VPWR.t202 VPWR pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4170 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN VGND.t3423 VGND.t3422 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4171 VPWR.t6231 a_66204_15704# a_66116_15748# VPWR.t6230 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4172 VPWR.t1590 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t1589 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4173 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN VGND.t3749 VGND.t3748 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4174 VGND.t6698 _251_.A1.t24 _228_.ZN VGND.t6697 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X4175 VPWR.t4265 a_51308_18407# a_51220_18504# VPWR.t4264 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4176 _379_.A2 uio_out[5].t10 a_20853_30644# VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4177 a_24540_23111# a_24452_23208# VGND.t4234 VGND.t4233 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4178 VPWR.t3427 a_33500_15271# a_33412_15368# VPWR.t1346 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4179 a_36860_15271# a_36772_15368# VGND.t4236 VGND.t4235 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4180 a_49292_13703# a_49204_13800# VGND.t4238 VGND.t4237 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4181 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I VGND.t5667 VGND.t5666 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4182 a_2364_18840# a_2276_18884# VGND.t3848 VGND.t557 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4183 VPWR.t3171 a_37980_26247# a_37892_26344# VPWR.t3170 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4184 _350_.A2.t18 _335_.ZN.t24 VPWR.t7001 VPWR.t7000 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4185 VPWR.t3812 a_33724_2727# a_33636_2824# VPWR.t3811 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4186 _474_.CLK.t18 a_48272_25156.t32 VGND.t6277 VGND.t6276 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X4187 a_13788_1592# a_13700_1636# VGND.t378 VGND.t377 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4188 a_34404_31048# _287_.A1.t25 uo_out[5].t4 VPWR.t6785 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4189 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I VGND.t4349 VGND.t4348 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4190 a_48384_26724# _474_.CLK.t44 VPWR.t6753 VPWR.t6752 pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X4191 a_62956_10567# a_62868_10664# VGND.t380 VGND.t379 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4192 a_46268_13703# a_46180_13800# VGND.t382 VGND.t381 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4193 VPWR.t3065 a_49404_30951# a_49316_31048# VPWR.t3064 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4194 VPWR.t3843 a_15580_29383# a_15492_29480# VPWR.t78 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4195 a_37756_1592# a_37668_1636# VGND.t384 VGND.t383 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4196 _386_.ZN _397_.A2.t12 a_47600_27912# VPWR.t7039 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4197 VPWR.t1746 a_5052_17272# a_4964_17316# VPWR.t1745 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4198 VPWR.t4094 _247_.B a_59172_27912# VPWR.t4093 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X4199 VPWR.t398 a_37084_26680# a_36996_26724# VPWR.t397 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4200 VPWR.t1043 a_20508_1159# a_20420_1256# VPWR.t1042 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4201 a_19276_23544# a_19188_23588# VGND.t4797 VGND.t4796 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4202 a_36656_29123# a_36284_29167# VGND.t4789 VGND.t4788 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X4203 VPWR.t4827 a_66652_7864# a_66564_7908# VPWR.t2731 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4204 VPWR.t779 a_27004_30951# a_26916_31048# VPWR.t778 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4205 a_28054_30196# _359_.B.t9 VPWR.t6773 VPWR.t6772 pfet_06v0 ad=0.5368p pd=3.32u as=0.4941p ps=2.03u w=1.22u l=0.5u
X4206 VPWR.t1255 _343_.A2 a_23834_28292# VPWR.t614 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X4207 VPWR.t6091 a_26780_1592# a_26692_1636# VPWR.t6090 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4208 VGND.t2154 a_51956_26183# a_51576_25896# VGND.t2153 nfet_06v0 ad=0.142p pd=1.14u as=0.176p ps=1.68u w=0.4u l=0.6u
X4209 VPWR.t117 _411_.A2.t10 a_47802_26724# VPWR.t116 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X4210 a_43804_1159# a_43716_1256# VGND.t4401 VGND.t4400 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4211 VPWR.t1498 a_53436_9432# a_53348_9476# VPWR.t1497 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4212 VPWR.t4945 a_63740_1159# a_63652_1256# VPWR.t1282 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4213 VPWR.t3954 a_48844_16839# a_48756_16936# VPWR.t3953 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4214 VPWR.t4015 a_35088_20893# a_35060_20569# VPWR.t4014 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X4215 VPWR.t5637 a_24428_23544# a_24340_23588# VPWR.t5636 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4216 VPWR.t284 a_44296_24393.t29 clkbuf_1_0__f_clk.I.t7 VPWR.t283 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4217 a_43916_16839# a_43828_16936# VGND.t4432 VGND.t4431 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4218 VPWR.t4579 a_66316_20408# a_66228_20452# VPWR.t4578 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4219 a_19164_30951# a_19076_31048# VGND.t4435 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4220 VPWR.t4582 a_14236_1159# a_14148_1256# VPWR.t1284 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4221 a_1020_12568# a_932_12612# VGND.t4438 VGND.t2006 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4222 VGND.t13 _397_.A1.t9 a_50120_26476# VGND.t12 nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4223 a_67996_18840# a_67908_18884# VGND.t3708 VGND.t3707 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4224 a_31820_20408# a_31732_20452# VGND.t5482 VGND.t5481 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4225 a_1020_7431# a_932_7528# VGND.t4439 VGND.t352 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4226 VPWR.t4587 a_21740_20408# a_21652_20452# VPWR.t4586 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4227 VPWR.t1008 a_66764_12135# a_66676_12232# VPWR.t1007 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4228 a_4940_10567# a_4852_10664# VGND.t4637 VGND.t4636 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4229 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN VPWR.t1404 VPWR.t1403 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4230 VPWR.t5280 a_47164_9432# a_47076_9476# VPWR.t5279 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4231 VPWR.t5631 a_55564_12135# a_55476_12232# VPWR.t5630 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4232 VPWR.t1791 a_37532_25112# a_37444_25156# VPWR.t1790 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4233 _311_.Z a_34980_22895# VGND.t3065 VGND.t3064 nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X4234 a_1916_10567# a_1828_10664# VGND.t4638 VGND.t3339 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4235 a_42908_2727# a_42820_2824# VGND.t4640 VGND.t4639 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4236 a_25332_28776# _454_.Q a_25124_28776# VGND.t3939 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4237 VPWR.t3232 a_57132_13703# a_57044_13800# VPWR.t3231 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4238 VGND.t2603 a_51620_19911# a_51240_19624# VGND.t2602 nfet_06v0 ad=0.142p pd=1.14u as=0.176p ps=1.68u w=0.4u l=0.6u
X4239 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I VGND.t4334 VGND.t4333 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4240 a_45820_18407# a_45732_18504# VGND.t4642 VGND.t4641 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4241 a_34396_18840# a_34308_18884# VGND.t3889 VGND.t3888 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4242 VPWR.t5538 a_48284_17272# a_48196_17316# VPWR.t5537 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4243 VGND.t5493 vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN VGND.t5492 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4244 a_2364_30951# a_2276_31048# VGND.t4742 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4245 VPWR.t3384 a_61948_2727# a_61860_2824# VPWR.t3383 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4246 VPWR.t4895 a_31820_21976# a_31732_22020# VPWR.t4894 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4247 VGND.t5475 a_35232_24029# a_35184_24073# VGND.t5474 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X4248 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN VGND.t3016 VGND.t3015 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4249 VPWR.t2442 a_37084_17272# a_36996_17316# VPWR.t2441 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4250 a_36636_2727# a_36548_2824# VGND.t4746 VGND.t4745 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4251 VPWR.t4899 a_39996_1159# a_39908_1256# VPWR.t4898 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4252 VGND.t5402 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN VGND.t5401 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4253 VPWR.t6287 _260_.A2 _260_.ZN VPWR.t6286 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4254 VPWR.t4901 a_20620_21976# a_20532_22020# VPWR.t4900 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4255 a_17932_26247# a_17844_26344# VGND.t4751 VGND.t2023 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4256 VPWR.t2343 a_36524_18407# a_36436_18504# VPWR.t2342 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4257 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN VGND.t5610 VGND.t5609 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4258 a_55452_12568# a_55364_12612# VGND.t4445 VGND.t4444 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4259 a_49600_30180# a_49152_30301.t5 a_50012_29977# VPWR.t6946 pfet_06v0 ad=0.1872p pd=1.4u as=43.2f ps=0.6u w=0.36u l=0.5u
X4260 VPWR.t2928 a_55676_2727# a_55588_2824# VPWR.t2927 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4261 a_17932_23111# a_17844_23208# VGND.t4446 VGND.t3411 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4262 VPWR.t3105 a_2364_5863# a_2276_5960# VPWR.t3104 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4263 a_19164_24679# a_19076_24776# VGND.t4448 VGND.t4447 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4264 VPWR.t6926 a_42392_22825.t28 _452_.CLK.t14 VPWR.t6925 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4265 VGND.t3643 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t3642 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4266 VPWR.t4595 a_58140_11000# a_58052_11044# VPWR.t4594 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4267 VPWR.t2904 a_2364_2727# a_2276_2824# VPWR.t1539 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4268 a_19164_21543# a_19076_21640# VGND.t4452 VGND.t4451 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4269 _349_.A4 a_26720_30301# VPWR.t4400 VPWR.t4399 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4270 VPWR.t3832 a_29468_1592# a_29380_1636# VPWR.t2690 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4271 a_6396_1592# a_6308_1636# VGND.t4244 VGND.t4243 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4272 a_67884_19975# a_67796_20072# VGND.t4246 VGND.t4245 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4273 VPWR.t3123 a_26556_21543# a_26468_21640# VPWR.t3122 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4274 a_16588_28248# a_16500_28292# VGND.t2077 VGND.t2076 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4275 _285_.Z _402_.A1.t17 a_39256_28292# VPWR.t6728 pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4276 a_63068_15271# a_62980_15368# VGND.t4248 VGND.t4247 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4277 VGND.t5913 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN VGND.t5912 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4278 a_62844_9432# a_62756_9476# VGND.t4250 VGND.t4249 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4279 VGND.t6699 _251_.A1.t25 _272_.B1 VGND.t102 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4280 VPWR.t3749 a_43580_27815# a_43492_27912# VPWR.t3748 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4281 a_2812_17272# a_2724_17316# VGND.t4251 VGND.t354 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4282 _284_.ZN.t10 _304_.B a_42168_25640.t6 VGND.t4536 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4283 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t6062 VPWR.t6061 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4284 VPWR.t617 a_36188_1159# a_36100_1256# VPWR.t616 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4285 uo_out[5].t10 _287_.A1.t26 a_33956_31048# VPWR.t6786 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4286 a_67100_15704# a_67012_15748# VGND.t618 VGND.t617 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4287 a_2364_24679# a_2276_24776# VGND.t620 VGND.t619 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4288 VGND.t330 a_56516_26344# _242_.Z VGND.t329 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4289 a_45596_30951# a_45508_31048# VGND.t621 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4290 VPWR.t624 a_1020_18840# a_932_18884# VPWR.t68 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4291 _475_.Q a_47776_20893# VPWR.t1908 VPWR.t1907 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4292 a_49172_27508# _470_.Q a_48988_27508# VGND.t4066 nfet_06v0 ad=0.1148p pd=1.1u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4293 a_37296_22020# _311_.Z VPWR.t4474 VPWR.t4473 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4294 VPWR.t1626 a_42368_28733# a_42340_28409# VPWR.t1625 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X4295 a_2364_21543# a_2276_21640# VGND.t641 VGND.t640 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4296 VPWR.t1104 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I VPWR.t1103 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4297 a_37584_29123# a_37291_29535# VPWR.t672 VPWR.t671 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X4298 _386_.A4 _383_.A2 VPWR.t1055 VPWR.t1054 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X4299 VPWR.t4194 a_1020_15704# a_932_15748# VPWR.t3340 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4300 VPWR.t4834 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t4833 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4301 VPWR.t4021 a_51196_1592# a_51108_1636# VPWR.t4020 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4302 VGND.t2480 vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN VGND.t2479 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4303 a_3260_9432# a_3172_9476# VGND.t647 VGND.t646 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4304 VGND.t5265 _323_.A3 _448_.D VGND.t5264 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X4305 VGND.t3910 vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN VGND.t3909 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4306 a_50068_27508# _407_.A1 _409_.ZN VGND.t525 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4307 a_3260_6296# a_3172_6340# VGND.t2621 VGND.t362 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4308 hold2.I _264_.B VGND.t2330 VGND.t2329 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X4309 VPWR.t3979 a_4940_27815# a_4852_27912# VPWR.t3978 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4310 VGND.t5672 _272_.A2 a_56804_30344# VGND.t325 nfet_06v0 ad=0.22595p pd=1.45u as=85.2f ps=0.95u w=0.71u l=0.6u
X4311 VPWR.t3702 a_6172_29383# a_6084_29480# VPWR.t3701 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4312 a_36148_21976# _301_.A1 VPWR.t3347 VPWR.t3346 pfet_06v0 ad=0.2354p pd=1.95u as=0.1391p ps=1.055u w=0.535u l=0.5u
X4313 a_41188_18840# _325_.A1.t16 VPWR.t6827 VPWR.t6826 pfet_06v0 ad=0.2354p pd=1.95u as=0.1391p ps=1.055u w=0.535u l=0.5u
X4314 a_28012_20408# a_27924_20452# VGND.t3091 VGND.t3090 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4315 VPWR.t3270 a_1916_27815# a_1828_27912# VPWR.t3269 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4316 a_58588_2727# a_58500_2824# VGND.t624 VGND.t444 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4317 VPWR.t5282 a_19724_25112# a_19636_25156# VPWR.t5281 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4318 a_39100_1159# a_39012_1256# VGND.t626 VGND.t625 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4319 a_47612_1159# a_47524_1256# VGND.t628 VGND.t627 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4320 VPWR.t4970 a_61164_13703# a_61076_13800# VPWR.t4969 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4321 VPWR.t632 a_66652_18840# a_66564_18884# VPWR.t631 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4322 a_32476_28776# _335_.ZN.t25 a_30388_28776# VGND.t835 nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4323 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I VGND.t1510 VGND.t1509 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4324 a_26672_30345# a_24452_30344.t7 a_26427_29977# VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4325 a_5276_2727# a_5188_2824# VGND.t632 VGND.t631 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4326 VGND.t2860 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN VGND.t2859 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4327 a_47612_30951# a_47524_31048# VGND.t5124 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4328 _355_.C.t1 a_28054_30196# VPWR.t890 VPWR.t889 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4329 VPWR.t3088 a_66652_15704# a_66564_15748# VPWR.t3087 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4330 VPWR.t5510 a_51532_10567# a_51444_10664# VPWR.t5509 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4331 a_25324_23544# a_25236_23588# VGND.t5126 VGND.t5125 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4332 VPWR.t5512 a_51756_18407# a_51668_18504# VPWR.t5511 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4333 VGND.t2906 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN VGND.t2905 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4334 _304_.B a_54432_31128# VPWR.t4674 VPWR.t4673 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4335 a_34844_17272# a_34756_17316# VGND.t5128 VGND.t5127 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4336 VGND.t2963 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN VGND.t2962 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4337 _433_.ZN _452_.Q.t13 VGND.t6640 VGND.t3771 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X4338 a_48308_23588# _474_.Q _399_.A2 VPWR.t4796 pfet_06v0 ad=0.3078p pd=1.68u as=0.2964p ps=1.66u w=1.14u l=0.5u
X4339 VPWR.t5952 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN VPWR.t5951 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4340 VGND.t5129 a_15460_31048# uio_oe[1].t0 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4341 a_34396_24679# a_34308_24776# VGND.t4551 VGND.t4550 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4342 VPWR.t4711 a_28012_21976# a_27924_22020# VPWR.t4710 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4343 VPWR.t1000 a_67324_15271# a_67236_15368# VPWR.t999 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4344 a_19372_30345# _465_.D a_19204_30345# VGND.t137 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X4345 a_29856_29123# a_29563_29535# VGND.t4898 VGND.t4897 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X4346 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I VGND.t4971 VGND.t4970 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4347 VPWR.t4713 a_33052_18840# a_32964_18884# VPWR.t4712 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4348 VPWR.t5649 a_51420_9432# a_51332_9476# VPWR.t5648 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4349 a_23196_24679# a_23108_24776# VGND.t4556 VGND.t4555 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4350 VPWR.t4716 a_48508_14136# a_48420_14180# VPWR.t1224 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4351 a_34396_21543# a_34308_21640# VGND.t4560 VGND.t4559 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4352 _474_.CLK.t19 a_48272_25156.t33 VGND.t6278 VGND.t18 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X4353 a_61052_14136# a_60964_14180# VGND.t2109 VGND.t2108 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4354 _397_.A2.t3 a_48104_30219# VGND.t2314 VGND.t71 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4355 VPWR.t3197 a_33052_15704# a_32964_15748# VPWR.t1968 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4356 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I VGND.t945 VGND.t944 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4357 VPWR.t1152 a_49852_30951# a_49764_31048# VPWR.t1151 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4358 VPWR.t4726 a_48508_11000# a_48420_11044# VPWR.t4725 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4359 a_23196_21543# a_23108_21640# VGND.t4569 VGND.t4568 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4360 a_13788_29383# a_13700_29480# VGND.t4571 VGND.t4570 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4361 a_1916_1159# a_1828_1256# VGND.t4573 VGND.t4572 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4362 VPWR.t945 a_61612_12135# a_61524_12232# VPWR.t944 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4363 a_61052_11000# a_60964_11044# VGND.t5803 VGND.t5802 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4364 a_36544_24419# a_36172_24463# VPWR.t5643 VPWR.t5642 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X4365 a_48284_15271# a_48196_15368# VGND.t4575 VGND.t4574 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4366 VGND.t6791 _223_.I _294_.ZN.t2 VGND.t6790 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4367 VPWR.t3651 a_4940_18407# a_4852_18504# VPWR.t3650 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4368 a_47172_27912# _386_.A4 VPWR.t646 VPWR.t645 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4369 VPWR.t3847 a_30588_21543# a_30500_21640# VPWR.t3846 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4370 _300_.ZN _300_.A2 VPWR.t959 VPWR.t958 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X4371 a_26556_27815# a_26468_27912# VGND.t862 VGND.t861 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4372 VGND.t6458 _474_.CLK.t45 _276_.A2 VGND.t3209 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X4373 _250_.B _230_.I.t11 a_64220_29098# VGND.t6347 nfet_06v0 ad=0.3124p pd=2.3u as=85.2f ps=0.95u w=0.71u l=0.6u
X4374 VPWR.t3632 a_45232_25987# a_45128_26031# VPWR.t3631 pfet_06v0 ad=0.1044p pd=0.94u as=0.1791p ps=1.355u w=0.36u l=0.5u
X4375 a_66204_8999# a_66116_9096# VGND.t864 VGND.t863 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4376 VPWR.t180 uio_in[0].t1 a_51791_30644# VPWR.t179 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4377 VPWR.t2986 a_1916_18407# a_1828_18504# VPWR.t2896 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4378 a_38876_19975# a_38788_20072# VGND.t866 VGND.t865 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4379 _393_.A3 _392_.A2 VPWR.t4360 VPWR.t4359 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X4380 a_18816_29931# a_18404_30344.t6 VGND.t140 VGND.t139 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4381 VPWR.t3061 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN VPWR.t3060 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4382 _264_.B _261_.ZN a_40468_25157# VPWR.t3568 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4383 VPWR.t6563 a_48272_25156.t34 _474_.CLK.t20 VPWR.t6562 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4384 VPWR.t2318 a_16252_30951# a_16164_31048# VPWR.t2317 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4385 a_66204_5863# a_66116_5960# VGND.t834 VGND.t833 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4386 a_46252_19759# _416_.ZN a_46128_20127# VPWR.t1113 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X4387 VPWR.t3645 a_24876_23544# a_24788_23588# VPWR.t3644 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4388 VGND.t392 a_18096_27165# uio_out[7].t6 VGND.t391 nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X4389 VPWR.t4809 a_66764_20408# a_66676_20452# VPWR.t4808 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4390 VPWR.t2988 a_10428_2727# a_10340_2824# VPWR.t2987 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4391 a_34620_2727# a_34532_2824# VGND.t4662 VGND.t4131 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4392 VPWR.t3925 a_4604_9432# a_4516_9476# VPWR.t3924 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4393 VPWR.t4813 a_37980_1159# a_37892_1256# VPWR.t4812 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4394 a_61500_12568# a_61412_12612# VGND.t4666 VGND.t4665 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4395 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN VPWR.t4841 VPWR.t4840 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4396 VPWR.t434 a_30160_30301# a_30132_29977# VPWR.t433 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X4397 a_18940_1159# a_18852_1256# VGND.t4668 VGND.t4667 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4398 VGND.t4995 _473_.Q _416_.A2 VGND.t4994 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X4399 VPWR.t4824 a_67436_19975# a_67348_20072# VPWR.t4823 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4400 VGND.t6280 a_48272_25156.t35 _474_.CLK.t21 VGND.t6279 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X4401 VPWR.t4658 a_53660_2727# a_53572_2824# VPWR.t4657 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4402 a_50300_12568# a_50212_12612# VGND.t4462 VGND.t4461 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4403 VPWR.t674 a_33724_1592# a_33636_1636# VPWR.t673 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4404 VPWR.t5822 a_57580_13703# a_57492_13800# VPWR.t5821 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4405 VPWR.t4617 a_33164_20408# a_33076_20452# VPWR.t4616 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4406 VPWR.t5793 a_28124_2727# a_28036_2824# VPWR.t5792 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4407 a_57692_1592# a_57604_1636# VGND.t4466 VGND.t4465 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4408 a_1916_29816# a_1828_29860# VGND.t4467 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4409 VPWR.t3490 _267_.ZN a_52292_29480# VPWR.t3489 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4410 a_40004_22020# _447_.Q.t11 VPWR.t6586 VPWR.t6585 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X4411 _399_.ZN _324_.B.t30 VGND.t6423 VGND.t6422 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X4412 VGND.t3689 _412_.A1 a_49764_26724# VGND.t3688 nfet_06v0 ad=0.104p pd=0.92u as=0.176p ps=1.68u w=0.4u l=0.6u
X4413 a_21044_27508# _346_.A2 _346_.ZN VGND.t3484 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4414 VPWR.t2496 a_64412_4295# a_64324_4392# VPWR.t2495 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4415 a_22636_28248# a_22548_28292# VGND.t2618 VGND.t2617 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4416 VPWR.t3520 a_40444_1159# a_40356_1256# VPWR.t3519 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4417 a_50524_1159# a_50436_1256# VGND.t4259 VGND.t4258 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4418 VPWR.t1489 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN VPWR.t1488 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4419 a_48580_27508# _470_.Q a_48376_27508# VGND.t4065 nfet_06v0 ad=0.1312p pd=1.14u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4420 VGND.t5745 _421_.A1 a_46620_22504# VGND.t248 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4421 VPWR.t3557 a_21404_21543# a_21316_21640# VPWR.t3556 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4422 a_1468_25112# a_1380_25156# VGND.t4260 VGND.t650 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4423 a_5388_18407# a_5300_18504# VGND.t4262 VGND.t4261 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4424 a_42392_22825.t9 clkbuf_1_0__f_clk.I.t49 VGND.t261 VGND.t260 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4425 a_1468_21976# a_1380_22020# VGND.t4609 VGND.t416 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4426 VPWR.t3042 a_62060_23111# a_61972_23208# VPWR.t3041 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4427 a_29804_30951# a_29716_31048# VGND.t1160 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4428 VPWR.t6689 a_41048_29816.t14 _459_.CLK.t4 VPWR.t6688 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4429 VPWR.t3426 a_34172_1159# a_34084_1256# VPWR.t912 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4430 _384_.A3.t4 _476_.Q VPWR.t4325 VPWR.t4324 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4431 a_36612_20072# _330_.A1.t17 _448_.D VPWR.t216 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4432 a_62396_26247# a_62308_26344# VGND.t1162 VGND.t1161 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4433 VPWR.t1887 a_18400_28733# a_18372_28409# VPWR.t1886 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X4434 VPWR.t5778 a_33948_18407# a_33860_18504# VPWR.t2941 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4435 VPWR.t1236 a_58140_1159# a_58052_1256# VPWR.t914 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4436 VGND.t949 _435_.A3 _264_.B VGND.t948 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X4437 a_4604_20408# a_4516_20452# VGND.t2647 VGND.t2646 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4438 VPWR.t6536 _362_.B.t13 _335_.ZN.t13 VPWR.t6535 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4439 VGND.t770 _252_.B _252_.ZN VGND.t769 nfet_06v0 ad=0.1209p pd=0.985u as=0.21175p ps=1.41u w=0.465u l=0.6u
X4440 a_42168_22504# _304_.B _324_.B.t9 VGND.t4535 nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X4441 a_16588_24679# a_16500_24776# VGND.t1166 VGND.t1165 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4442 _245_.I1 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t1068 VPWR.t1067 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4443 VPWR.t6479 _459_.CLK.t32 a_27588_29159.t0 VPWR.t6478 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4444 VGND.t6425 _324_.B.t31 a_45564_21236# VGND.t6424 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4445 a_16588_21543# a_16500_21640# VGND.t1079 VGND.t1005 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4446 a_44296_24393.t8 clk.t8 VGND.t6529 VGND.t6528 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4447 a_59932_1159# a_59844_1256# VGND.t2425 VGND.t2424 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4448 a_32836_27208# _358_.A3 VGND.t469 VGND.t468 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4449 a_62844_2727# a_62756_2824# VGND.t2533 VGND.t2532 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4450 a_1916_23544# a_1828_23588# VGND.t2534 VGND.t2281 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4451 VPWR.t3770 a_58924_17272# a_58836_17316# VPWR.t3769 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4452 VPWR.t5513 a_1020_29383# a_932_29480# VPWR.t86 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4453 a_19948_27815# a_19860_27912# VGND.t351 VGND.t350 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4454 a_52400_25987.t0 _474_.CLK.t46 VPWR.t6755 VPWR.t6754 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X4455 VPWR.t3808 a_54108_12568# a_54020_12612# VPWR.t3807 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4456 a_61836_25515# _251_.A1.t26 a_62404_25640# VGND.t6700 nfet_06v0 ad=0.2132p pd=1.34u as=98.39999f ps=1.06u w=0.82u l=0.6u
X4457 VPWR.t2672 a_4604_21976# a_4516_22020# VPWR.t2671 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4458 a_56572_2727# a_56484_2824# VGND.t1168 VGND.t1167 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4459 VPWR.t2282 a_1020_26247# a_932_26344# VPWR.t2281 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4460 VPWR.t5186 a_67772_24679# a_67684_24776# VPWR.t5185 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4461 VPWR.t2288 a_31484_30951# a_31396_31048# VPWR.t2287 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4462 VPWR.t2401 vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I VPWR.t2400 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4463 a_1468_15704# a_1380_15748# VGND.t1170 VGND.t1169 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4464 VPWR.t2821 a_1020_23111# a_932_23208# VPWR.t1899 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4465 a_3260_2727# a_3172_2824# VGND.t1172 VGND.t1171 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4466 a_51332_24372# _424_.B1.t12 VGND.t6335 VGND.t183 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4467 VPWR.t1582 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t1581 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4468 VGND.t335 a_59955_30600# _237_.A1 VGND.t34 nfet_06v0 ad=0.28262p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4469 VPWR.t1915 a_2364_4728# a_2276_4772# VPWR.t383 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4470 VPWR.t6959 _452_.Q.t14 a_42154_21236# VPWR.t6958 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4471 a_11548_29816# a_11460_29860# VGND.t1173 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4472 a_4604_14136# a_4516_14180# VGND.t2607 VGND.t2606 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4473 a_5724_1159# a_5636_1256# VGND.t2115 VGND.t2114 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4474 _452_.CLK.t15 a_42392_22825.t29 VGND.t6609 VGND.t6608 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X4475 VPWR.t5405 a_53548_24679# a_53460_24776# VPWR.t5404 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4476 VPWR.t357 a_2364_1592# a_2276_1636# VPWR.t356 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4477 a_21852_1159# a_21764_1256# VGND.t5488 VGND.t5487 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4478 a_13340_1159# a_13252_1256# VGND.t5490 VGND.t5489 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4479 a_25420_30345# _342_.ZN a_25252_30345# VGND.t137 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X4480 a_38575_24072# _439_.ZN VGND.t5850 VGND.t5849 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4481 VGND.t1113 a_48529_22460# _279_.Z VGND.t1112 nfet_06v0 ad=0.2288p pd=1.58u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4482 a_4604_11000# a_4516_11044# VGND.t4364 VGND.t4363 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4483 VPWR.t2063 a_62396_1159# a_62308_1256# VPWR.t2062 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4484 a_28460_20408# a_28372_20452# VGND.t4368 VGND.t4367 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4485 VPWR.t2165 _431_.A3 _441_.A3 VPWR.t2164 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4486 a_65532_15271# a_65444_15368# VGND.t5491 VGND.t3616 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4487 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN VPWR.t3096 VPWR.t3095 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4488 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I _274_.A1 VPWR.t2656 VPWR.t2655 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4489 VGND.t1295 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I VGND.t1294 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4490 a_33148_25641# _460_.D a_32980_25641# VGND.t5817 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X4491 _337_.A3.t0 a_26160_27165# VPWR.t949 VPWR.t948 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4492 a_63336_29480# vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN VPWR.t4871 VPWR.t4870 pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4493 a_58656_27912# _242_.Z _243_.ZN VPWR.t2508 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4494 VPWR.t3282 a_44700_30951# a_44612_31048# VPWR.t3281 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4495 a_9308_29816# a_9220_29860# VGND.t431 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4496 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN _245_.I1 VPWR.t5411 VPWR.t5410 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4497 a_57916_25112# a_57828_25156# VGND.t433 VGND.t432 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4498 VGND.t3073 a_40264_30320# _294_.A2.t1 VGND.t3072 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X4499 a_57244_9432# a_57156_9476# VGND.t435 VGND.t434 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4500 VPWR.t5450 a_51980_10567# a_51892_10664# VPWR.t5449 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4501 a_25772_23544# a_25684_23588# VGND.t437 VGND.t436 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4502 a_43132_15271# a_43044_15368# VGND.t439 VGND.t438 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4503 a_62508_12135# a_62420_12232# VGND.t5381 VGND.t5380 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4504 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN VGND.t2478 VGND.t2477 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4505 _245_.Z a_61836_25515# VPWR.t2596 VPWR.t2595 pfet_06v0 ad=0.3477p pd=1.79u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4506 VPWR.t5992 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN VPWR.t5991 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4507 VPWR.t4124 a_12548_31048# a_12548_31048# VPWR.t4123 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4508 VPWR.t3615 a_28460_21976# a_28372_22020# VPWR.t3614 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4509 VPWR.t4955 a_30924_23544# a_30836_23588# VPWR.t4954 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4510 a_50084_24328# _398_.C a_50724_24908# VPWR.t3310 pfet_06v0 ad=0.2464p pd=2u as=0.1736p ps=1.18u w=0.56u l=0.5u
X4511 VPWR.t4070 a_67772_15271# a_67684_15368# VPWR.t4069 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4512 VPWR.t4554 a_3708_24679# a_3620_24776# VPWR.t1139 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4513 a_24980_25273# a_23668_25640.t4 a_24636_25641# VPWR.t7029 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X4514 uo_out[5].t1 _290_.ZN VGND.t1140 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4515 _270_.A2 a_58911_30644# VPWR.t2922 VPWR.t2921 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X4516 VPWR.t5424 a_49896_18909# a_51252_19001# VPWR.t5423 pfet_06v0 ad=0.4554p pd=3.25u as=54f ps=0.66u w=0.36u l=0.5u
X4517 a_16140_25112# a_16052_25156# VGND.t3462 VGND.t2294 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4518 VPWR.t3618 a_48956_14136# a_48868_14180# VPWR.t3617 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4519 VPWR.t3619 a_16700_1159# a_16612_1256# VPWR.t1145 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4520 a_37384_19624# _319_.A3 VPWR.t2705 VPWR.t2704 pfet_06v0 ad=0.156p pd=1.12u as=0.40575p ps=2.055u w=0.6u l=0.5u
X4521 VPWR.t3621 a_61612_20408# a_61524_20452# VPWR.t3620 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4522 a_14460_30951# a_14372_31048# VGND.t545 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4523 a_36284_29167# _462_.D a_36160_29535# VPWR.t3561 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X4524 a_43564_27209# _470_.D a_43440_26841# VPWR.t5514 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X4525 a_22636_30951# a_22548_31048# VGND.t546 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4526 a_16140_21976# a_16052_22020# VGND.t3213 VGND.t2300 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4527 VPWR.t548 a_48956_11000# a_48868_11044# VPWR.t547 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4528 VPWR.t4620 a_1916_29816# a_1828_29860# VPWR.t1999 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4529 VPWR.t4002 a_45372_15271# a_45284_15368# VPWR.t1147 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4530 a_12444_1592# a_12356_1636# VGND.t550 VGND.t549 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4531 a_62404_25156# _245_.I1 VPWR.t5409 VPWR.t5408 pfet_06v0 ad=0.4758p pd=2u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4532 a_54332_1159# a_54244_1256# VGND.t2809 VGND.t2808 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4533 a_62844_1159# a_62756_1256# VGND.t4021 VGND.t4020 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4534 a_5052_28248# a_4964_28292# VGND.t1750 VGND.t1749 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4535 _274_.A2 _268_.A2.t6 VGND.t6747 VGND.t325 nfet_06v0 ad=0.21175p pd=1.41u as=0.22595p ps=1.45u w=0.465u l=0.6u
X4536 VPWR.t963 a_1916_26680# a_1828_26724# VPWR.t962 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4537 a_36412_1592# a_36324_1636# VGND.t1721 VGND.t1720 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4538 a_37888_27555# a_37516_27599# VGND.t891 VGND.t890 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X4539 _389_.ZN _381_.Z VGND.t3803 VGND.t3802 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4540 a_47252_18884# _416_.A2 a_47028_18884# VPWR.t6290 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4541 _402_.ZN _402_.B VGND.t3125 VGND.t3124 nfet_06v0 ad=0.2569p pd=1.56u as=0.2244p ps=1.9u w=0.51u l=0.6u
X4542 a_24692_27209# a_23892_27208.t5 VGND.t6068 VGND.t6067 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4543 a_3260_18407# a_3172_18504# VGND.t1723 VGND.t1722 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4544 VGND.t1610 _495_.I a_41160_29083# VGND.t1609 nfet_06v0 ad=0.2662p pd=2.09u as=0.51425p ps=2.91u w=0.605u l=0.6u
X4545 a_63068_18840# a_62980_18884# VGND.t1569 VGND.t1022 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4546 a_39669_21236# _448_.Q.t10 a_39475_21236# VGND.t6577 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X4547 a_63721_28776# _230_.I.t12 _250_.A2 VGND.t6348 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X4548 VPWR.t6481 _459_.CLK.t33 a_24452_30344.t0 VPWR.t6480 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4549 a_66988_16839# a_66900_16936# VGND.t1725 VGND.t1724 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4550 a_25643_25273# a_24080_25227# a_25008_25597# VGND.t4263 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4551 a_62564_29032# _229_.I.t10 VPWR.t6875 VPWR.t6874 pfet_06v0 ad=0.1456p pd=1.08u as=0.34437p ps=1.895u w=0.56u l=0.5u
X4552 VPWR.t4404 a_67884_19975# a_67796_20072# VPWR.t4403 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4553 a_52247_31220# a_51791_30644# VPWR.t5456 VPWR.t5455 pfet_06v0 ad=61.19999f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4554 VGND.t4687 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_57276_27208# VGND.t4686 nfet_06v0 ad=0.2132p pd=1.34u as=98.39999f ps=1.06u w=0.82u l=0.6u
X4555 VPWR.t3693 a_3708_15271# a_3620_15368# VPWR.t1970 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4556 _238_.ZN _238_.I VGND.t2131 VGND.t2130 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X4557 VPWR.t6225 a_20956_1159# a_20868_1256# VPWR.t6224 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4558 VPWR.t1818 a_19948_20408# a_19860_20452# VPWR.t1817 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4559 _359_.B.t0 a_45088_29123# VPWR.t4451 VPWR.t4450 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4560 a_40668_20408# a_40580_20452# VGND.t1742 VGND.t1741 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4561 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I VPWR.t1492 VPWR.t1491 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4562 a_8860_1592# a_8772_1636# VGND.t1729 VGND.t1728 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4563 a_58924_12135# a_58836_12232# VGND.t3120 VGND.t3119 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4564 VPWR.t2675 a_21852_21543# a_21764_21640# VPWR.t2674 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4565 a_21292_20408# a_21204_20452# VGND.t1717 VGND.t1716 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4566 a_5052_18840# a_4964_18884# VGND.t2529 VGND.t2528 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4567 VPWR.t6122 a_53884_9432# a_53796_9476# VPWR.t6121 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4568 _460_.Q a_34448_25597# VPWR.t3869 VPWR.t3868 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4569 a_11324_2727# a_11236_2824# VGND.t1731 VGND.t1730 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4570 VPWR.t6096 a_1916_17272# a_1828_17316# VPWR.t2961 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4571 _427_.B1 a_52452_24072# VGND.t5218 VGND.t5217 nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X4572 VPWR.t3046 a_25232_27165# a_25204_26841# VPWR.t3045 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X4573 a_40668_1592# a_40580_1636# VGND.t1052 VGND.t1051 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4574 VPWR.t1485 a_14684_1159# a_14596_1256# VPWR.t1484 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4575 VGND.t4404 _330_.A2 _330_.ZN VGND.t4403 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4576 _474_.CLK.t22 a_48272_25156.t36 VGND.t6282 VGND.t6281 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X4577 a_54604_23263# a_54088_22895# VPWR.t2933 VPWR.t2932 pfet_06v0 ad=43.2f pd=0.6u as=0.1044p ps=0.94u w=0.36u l=0.5u
X4578 VGND.t5804 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t1192 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4579 a_64636_1592# a_64548_1636# VGND.t1054 VGND.t1053 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4580 VPWR.t2045 a_37584_29123# _334_.A1 VPWR.t2044 pfet_06v0 ad=0.854p pd=3.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4581 a_24780_28776# _343_.A2 VGND.t1181 VGND.t1180 nfet_06v0 ad=58.39999f pd=0.685u as=0.23405p ps=1.555u w=0.365u l=0.6u
X4582 VPWR.t3328 a_30364_2727# a_30276_2824# VPWR.t3327 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4583 a_9532_1159# a_9444_1256# VGND.t443 VGND.t442 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4584 VPWR.t1246 a_11548_29816# a_11460_29860# VPWR.t1245 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4585 VPWR.t3334 a_59372_10567# a_59284_10664# VPWR.t3333 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4586 VPWR.t4266 a_65308_8999# a_65220_9096# VPWR.t1342 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4587 a_25660_1159# a_25572_1256# VGND.t5989 VGND.t5988 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4588 VPWR.t5659 a_61052_27815# a_60964_27912# VPWR.t5658 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4589 VPWR.t5171 a_54332_2727# a_54244_2824# VPWR.t5170 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4590 VPWR.t2611 a_1020_5863# a_932_5960# VPWR.t2610 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4591 vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t2395 VPWR.t2394 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4592 a_28908_21976# a_28820_22020# VGND.t2806 VGND.t2805 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4593 a_29020_2727# a_28932_2824# VGND.t596 VGND.t595 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4594 VPWR.t599 a_18828_21976# a_18740_22020# VPWR.t598 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4595 a_41088_17757.t1 _452_.CLK.t48 VGND.t6368 VGND.t6367 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4596 a_38472_30169# _284_.ZN.t31 VPWR.t6520 VPWR.t6519 pfet_06v0 ad=0.2542p pd=1.44u as=0.428p ps=2.02u w=0.82u l=0.5u
X4597 a_28112_27912# _371_.A2 a_27908_27912# VPWR.t3581 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4598 VPWR.t5002 _475_.Q a_49068_20408# VPWR.t5001 pfet_06v0 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X4599 a_31372_21976# a_31284_22020# VGND.t1981 VGND.t1980 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4600 _424_.B1.t2 _324_.C.t23 VPWR.t6803 VPWR.t6802 pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4601 a_20172_25112# a_20084_25156# VGND.t600 VGND.t599 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4602 VPWR.t3514 a_15244_26247# a_15156_26344# VPWR.t2466 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4603 VPWR.t3077 a_1020_2727# a_932_2824# VPWR.t3076 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4604 VPWR.t2587 _379_.Z a_17786_29480# VPWR.t2586 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X4605 a_20250_31048# uio_out[5].t11 _465_.D VPWR.t6899 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4606 VPWR.t3320 a_48060_2727# a_47972_2824# VPWR.t3319 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4607 a_55744_22505# a_55208_22505# VGND.t5894 VGND.t5893 nfet_06v0 ad=43.2f pd=0.6u as=0.2637p ps=1.825u w=0.36u l=0.6u
X4608 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I VPWR.t919 VPWR.t918 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4609 a_46604_16839# a_46516_16936# VGND.t602 VGND.t601 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4610 VPWR.t4098 a_27116_23544# a_27028_23588# VPWR.t4097 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4611 VPWR.t4099 a_28124_1592# a_28036_1636# VPWR.t3136 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4612 a_20172_21976# a_20084_22020# VGND.t2070 VGND.t2069 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4613 VPWR.t3813 a_15244_23111# a_15156_23208# VPWR.t3803 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4614 a_5052_1592# a_4964_1636# VGND.t4924 VGND.t4923 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4615 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I VGND.t1423 VGND.t1422 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4616 VPWR.t443 a_9308_29816# a_9220_29860# VPWR.t442 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4617 VPWR.t6237 a_50076_9432# a_49988_9476# VPWR.t6236 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4618 VPWR.t5081 a_60380_1159# a_60292_1256# VPWR.t821 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4619 a_24468_25641# a_23668_25640.t5 VGND.t6709 VGND.t6708 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4620 _352_.A2.t9 _350_.A1.t8 a_28596_27916.t9 VPWR.t6625 pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X4621 a_61500_9432# a_61412_9476# VGND.t4928 VGND.t4927 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4622 VPWR.t6209 a_54556_12568# a_54468_12612# VPWR.t6208 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4623 a_49936_19325.t0 _474_.CLK.t47 VPWR.t6757 VPWR.t6756 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X4624 VPWR.t3205 a_45820_13703# a_45732_13800# VPWR.t3204 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4625 a_43796_18559# a_42484_18183.t3 a_43452_18191# VPWR.t7046 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X4626 VPWR.t2594 a_61836_25515# _245_.Z VPWR.t2593 pfet_06v0 ad=0.4392p pd=1.94u as=0.3477p ps=1.79u w=1.22u l=0.5u
X4627 VGND.t5871 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I VGND.t5870 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4628 a_59143_31198# a_58687_31220# a_58911_30644# VPWR.t5521 pfet_06v0 ad=61.19999f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X4629 VPWR.t3907 a_61500_26247# a_61412_26344# VPWR.t3906 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4630 a_34716_20937# _319_.ZN a_34548_20937# VGND.t2573 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X4631 a_31820_23544# a_31732_23588# VGND.t693 VGND.t692 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4632 a_64860_26247# a_64772_26344# VGND.t695 VGND.t694 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4633 VPWR.t6185 a_7516_2727# a_7428_2824# VPWR.t6184 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4634 a_42404_17433# _452_.D a_41536_17636# VPWR.t2636 pfet_06v0 ad=54f pd=0.66u as=0.1872p ps=1.4u w=0.36u l=0.5u
X4635 _384_.ZN _473_.Q VGND.t4993 VGND.t4992 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X4636 VGND.t201 _416_.A1.t9 _444_.D VGND.t200 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X4637 a_11996_29816# a_11908_29860# VGND.t696 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4638 _455_.Q.t1 a_22352_25987# VGND.t3851 VGND.t3850 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4639 VPWR.t5638 a_33948_17272# a_33860_17316# VPWR.t651 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4640 a_20620_23544# a_20532_23588# VGND.t698 VGND.t697 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4641 a_42168_25640.t5 _304_.B _284_.ZN.t9 VGND.t4534 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4642 VPWR.t6730 _402_.A1.t18 _411_.A2.t6 VPWR.t6729 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4643 VPWR.t6128 a_53996_24679# a_53908_24776# VPWR.t502 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4644 VPWR.t432 a_6844_1592# a_6756_1636# VPWR.t431 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4645 a_58140_1159# a_58052_1256# VGND.t1164 VGND.t1163 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4646 a_66652_1159# a_66564_1256# VGND.t700 VGND.t699 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4647 a_63516_17272# a_63428_17316# VGND.t702 VGND.t701 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4648 VGND.t1950 a_37584_29123# a_37536_29167# VGND.t1949 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X4649 _238_.I _246_.B2 VPWR.t5211 VPWR.t5210 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X4650 a_40992_17433# a_40040_17675# VPWR.t5251 VPWR.t5250 pfet_06v0 ad=50.4f pd=0.64u as=0.23p ps=1.54u w=0.36u l=0.5u
X4651 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN VPWR.t1388 VPWR.t1387 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4652 VPWR.t7019 _251_.A1.t27 a_59652_25640# VPWR.t7018 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4653 VPWR.t5684 a_62620_15271# a_62532_15368# VPWR.t809 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4654 a_65980_15271# a_65892_15368# VGND.t727 VGND.t726 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4655 a_52316_17272# a_52228_17316# VGND.t729 VGND.t728 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4656 _439_.ZN _260_.A1 VGND.t3772 VGND.t3771 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4657 a_4156_7431# a_4068_7528# VGND.t731 VGND.t730 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4658 a_58140_12568# a_58052_12612# VGND.t733 VGND.t732 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4659 VPWR.t747 a_1916_6296# a_1828_6340# VPWR.t746 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4660 a_33276_2727# a_33188_2824# VGND.t736 VGND.t735 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4661 VPWR.t886 a_38876_19975# a_38788_20072# VPWR.t885 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4662 VPWR.t6928 a_42392_22825.t30 _452_.CLK.t16 VPWR.t6927 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4663 a_9756_29816# a_9668_29860# VGND.t737 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4664 VPWR.t1656 a_1916_3160# a_1828_3204# VPWR.t964 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4665 VPWR.t698 a_1020_28248# a_932_28292# VPWR.t697 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4666 VPWR.t2845 a_40220_15271# a_40132_15368# VPWR.t2844 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4667 VGND.t6611 a_42392_22825.t31 _452_.CLK.t17 VGND.t6610 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X4668 a_43580_15271# a_43492_15368# VGND.t689 VGND.t688 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4669 VPWR.t5461 a_40464_27165# a_40436_26841# VPWR.t5460 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X4670 VPWR.t6132 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I VPWR.t6131 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4671 a_62956_12135# a_62868_12232# VGND.t1531 VGND.t1530 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4672 a_20060_23111# a_19972_23208# VGND.t691 VGND.t690 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4673 VPWR.t4949 a_56348_1592# a_56260_1636# VPWR.t4948 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4674 VPWR.t5344 a_1020_25112# a_932_25156# VPWR.t1013 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4675 VGND.t6471 _359_.B.t10 _461_.D VGND.t38 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X4676 VPWR.t1371 a_29244_21543# a_29156_21640# VPWR.t1370 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4677 a_62560_25112# _251_.A1.t28 VGND.t6702 VGND.t6701 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4678 a_23084_29383# a_22996_29480# VGND.t790 VGND.t491 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4679 VGND.t859 a_54420_21976# a_54040_22366# VGND.t858 nfet_06v0 ad=0.142p pd=1.14u as=0.176p ps=1.68u w=0.4u l=0.6u
X4680 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I VPWR.t1512 VPWR.t1511 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4681 a_55228_27815# a_55140_27912# VGND.t983 VGND.t982 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4682 VPWR.t5154 _473_.Q a_49068_20408# VPWR.t5153 pfet_06v0 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X4683 _424_.B1.t0 _399_.ZN VPWR.t1263 VPWR.t1262 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X4684 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I VPWR.t5338 VPWR.t5337 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4685 vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t2119 VGND.t2118 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4686 VPWR.t4971 a_64748_23544# a_64660_23588# VPWR.t62 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4687 a_20060_1159# a_19972_1256# VGND.t5190 VGND.t5189 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4688 a_44028_27815# a_43940_27912# VGND.t920 VGND.t919 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4689 a_37196_23544# a_37108_23588# VGND.t5192 VGND.t5191 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4690 _352_.A2.t0 _350_.A2.t25 a_28596_27916.t0 VPWR.t6577 pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X4691 _229_.I.t0 a_62532_30736# VPWR.t2530 VPWR.t2529 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X4692 a_61836_16839# a_61748_16936# VGND.t5194 VGND.t5193 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4693 VGND.t314 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN VGND.t313 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4694 a_4940_15271# a_4852_15368# VGND.t5196 VGND.t5195 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4695 a_49492_18840# a_49896_18909# a_49840_19001# VPWR.t5422 pfet_06v0 ad=0.1665p pd=1.285u as=50.4f ps=0.64u w=0.36u l=0.5u
X4696 VPWR.t4748 a_33612_24679# a_33524_24776# VPWR.t4747 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4697 VPWR.t6640 _230_.I.t13 _252_.B VPWR.t6639 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4698 a_4940_12135# a_4852_12232# VGND.t5811 VGND.t5810 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4699 VPWR.t111 _294_.A2.t7 a_34586_27912# VPWR.t110 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X4700 a_1916_15271# a_1828_15368# VGND.t5197 VGND.t4153 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4701 a_31260_16839# a_31172_16936# VGND.t5198 VGND.t4110 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4702 a_35232_24029# a_34939_23705# VGND.t683 VGND.t682 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X4703 VPWR.t4476 a_44364_16839# a_44276_16936# VPWR.t326 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4704 a_51620_19911# a_52024_20083# a_51968_20127# VPWR.t439 pfet_06v0 ad=0.1665p pd=1.285u as=50.4f ps=0.64u w=0.36u l=0.5u
X4705 VPWR.t5910 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN VPWR.t5909 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4706 a_37980_1159# a_37892_1256# VGND.t4664 VGND.t4663 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4707 _302_.Z a_38576_22504# VPWR.t5824 VPWR.t5823 pfet_06v0 ad=0.5368p pd=3.32u as=0.395p ps=2.02u w=1.22u l=0.5u
X4708 a_16672_26841# a_16240_26795# VPWR.t5616 VPWR.t5615 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X4709 a_1916_12135# a_1828_12232# VGND.t5233 VGND.t1708 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4710 a_44961_27912# _400_.ZN _470_.D VPWR.t803 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4711 a_28596_27916.t6 _371_.A2 VPWR.t3580 VPWR.t3579 pfet_06v0 ad=0.48p pd=2u as=0.312p ps=1.72u w=1.2u l=0.5u
X4712 VPWR.t6805 _324_.C.t24 _325_.B VPWR.t6804 pfet_06v0 ad=0.2561p pd=1.505u as=0.44325p ps=2.87u w=0.985u l=0.5u
X4713 a_19696_30345# a_18816_29931# a_19372_30345# VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X4714 VPWR.t3354 a_51084_12135# a_50996_12232# VPWR.t3353 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4715 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I VPWR.t3461 VPWR.t3460 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4716 VPWR.t5197 a_3708_23544# a_3620_23588# VPWR.t5196 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4717 VPWR.t4641 a_65420_10567# a_65332_10664# VPWR.t4640 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4718 VPWR.t4642 a_2364_10567# a_2276_10664# VPWR.t1352 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4719 a_62620_1592# a_62532_1636# VGND.t754 VGND.t753 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4720 VGND.t5899 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I VGND.t5898 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4721 VGND.t645 _386_.A4 _389_.ZN VGND.t644 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4722 a_48732_17272# a_48644_17316# VGND.t756 VGND.t755 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4723 VGND.t5534 a_56964_26724# _241_.Z VGND.t5533 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4724 VPWR.t4644 a_54220_10567# a_54132_10664# VPWR.t4643 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4725 a_28012_23544# a_27924_23588# VGND.t571 VGND.t360 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4726 uo_out[3].t0 a_41160_29083# VPWR.t4182 VPWR.t4181 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4727 VPWR.t4646 a_54444_18407# a_54356_18504# VPWR.t4645 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4728 a_37532_17272# a_37444_17316# VGND.t573 VGND.t572 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4729 a_32380_1592# a_32292_1636# VGND.t574 VGND.t367 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4730 a_45708_17272# a_45620_17316# VGND.t576 VGND.t575 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4731 _336_.A2.t1 a_25936_25597# VGND.t5633 VGND.t5632 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4732 uo_out[0].t1 _296_.ZN VGND.t3514 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4733 VPWR.t4331 a_24988_24679# a_24900_24776# VPWR.t4330 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4734 a_66652_8999# a_66564_9096# VGND.t578 VGND.t577 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4735 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I VGND.t4338 VGND.t4337 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4736 a_48508_12568# a_48420_12612# VGND.t580 VGND.t579 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4737 a_52304_26399# a_51576_25896# VPWR.t2262 VPWR.t2261 pfet_06v0 ad=50.4f pd=0.64u as=0.23p ps=1.54u w=0.36u l=0.5u
X4738 a_37084_21543# a_36996_21640# VGND.t5418 VGND.t5417 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4739 a_32828_23111# a_32740_23208# VGND.t582 VGND.t581 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4740 a_66652_5863# a_66564_5960# VGND.t5773 VGND.t2471 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4741 VGND.t4255 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN VGND.t4254 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4742 a_33540_22505# a_32740_22504.t5 VGND.t95 VGND.t94 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4743 a_59332_29816# _324_.C.t25 a_59948_30352# VGND.t3682 nfet_06v0 ad=0.1672p pd=1.64u as=60.8f ps=0.7u w=0.38u l=0.6u
X4744 VPWR.t5379 a_10876_2727# a_10788_2824# VPWR.t5378 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4745 a_57220_29861# _255_.ZN VPWR.t5269 VPWR.t5268 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4746 VGND.t2272 a_36148_21976# _317_.A2 VGND.t2271 nfet_06v0 ad=0.2424p pd=1.635u as=0.341p ps=2.43u w=0.775u l=0.6u
X4747 a_67741_30600# ena.t0 VPWR.t6818 VPWR.t6817 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4748 VPWR.t3094 a_64300_12135# a_64212_12232# VPWR.t3093 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4749 VPWR.t708 a_11996_29816# a_11908_29860# VPWR.t707 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4750 a_33948_15271# a_33860_15368# VGND.t3449 VGND.t3448 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4751 a_54332_18840# a_54244_18884# VGND.t4543 VGND.t4542 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4752 VPWR.t5010 a_37888_27555# a_37860_27967# VPWR.t5009 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X4753 VPWR.t5222 a_33276_21543# a_33188_21640# VPWR.t5221 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4754 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN VGND.t4456 VGND.t71 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4755 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I VGND.t2378 VGND.t2377 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4756 a_5388_7431# a_5300_7528# VGND.t3451 VGND.t3450 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4757 VPWR.t5695 vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN VPWR.t5694 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4758 VGND.t3754 a_34304_24029# a_34256_24073# VGND.t3753 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X4759 VPWR.t5215 a_15692_26247# a_15604_26344# VPWR.t5214 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4760 VPWR.t4345 a_28572_2727# a_28484_2824# VPWR.t4344 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4761 VPWR.t5217 a_23868_26247# a_23780_26344# VPWR.t5216 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4762 VPWR.t1730 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I VPWR.t1729 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4763 a_17786_29480# _355_.C.t13 _467_.D VPWR.t6674 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4764 clkbuf_1_0__f_clk.I.t24 a_44296_24393.t30 VGND.t281 VGND.t280 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X4765 VPWR.t1160 a_27564_23544# a_27476_23588# VPWR.t1159 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4766 VPWR.t3117 a_64860_4295# a_64772_4392# VPWR.t3116 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4767 VPWR.t5220 a_15692_23111# a_15604_23208# VPWR.t1735 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4768 a_52891_28776# _267_.A1 _267_.ZN VGND.t5600 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4769 a_36948_29860# _287_.A1.t27 uo_out[2].t0 VPWR.t6787 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4770 VPWR.t1634 a_40892_1159# a_40804_1256# VPWR.t1633 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4771 VPWR.t696 a_9756_29816# a_9668_29860# VPWR.t695 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4772 a_51428_20452# _419_.Z a_51240_20452# VPWR.t4462 pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X4773 a_55724_22137# a_55208_22505# VPWR.t6158 VPWR.t6157 pfet_06v0 ad=43.2f pd=0.6u as=0.1044p ps=0.94u w=0.36u l=0.5u
X4774 a_44961_27912# _403_.ZN VPWR.t3730 VPWR.t3729 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4775 VPWR.t974 _435_.A3 a_40468_25157# VPWR.t973 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X4776 VPWR.t2769 _275_.A2 a_51050_29480# VPWR.t2768 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X4777 _324_.B.t17 _304_.ZN.t15 VPWR.t232 VPWR.t231 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4778 a_67741_30600# ena.t1 VGND.t6512 VGND.t45 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4779 VGND.t148 _294_.ZN.t6 uo_out[4].t10 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4780 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[1\].I VGND.t1347 VGND.t1346 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4781 VPWR.t5583 a_55228_20408# a_55140_20452# VPWR.t5582 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4782 _421_.B _474_.Q a_47732_22504# VGND.t4651 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4783 VPWR.t5119 _438_.A2 a_38616_24328# VPWR.t5118 pfet_06v0 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X4784 a_48516_24080# _397_.Z VGND.t870 VGND.t869 nfet_06v0 ad=93.59999f pd=1.02u as=0.3432p ps=2.44u w=0.78u l=0.6u
X4785 VPWR.t262 clkbuf_1_0__f_clk.I.t50 a_48272_25156.t3 VPWR.t261 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X4786 a_32380_1159# a_32292_1256# VGND.t4709 VGND.t4708 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4787 a_40892_1159# a_40804_1256# VGND.t1552 VGND.t1551 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4788 a_4604_29816# a_4516_29860# VGND.t744 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4789 a_62060_13703# a_61972_13800# VGND.t746 VGND.t745 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4790 a_35068_1592# a_34980_1636# VGND.t748 VGND.t747 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4791 a_65644_23544# a_65556_23588# VGND.t750 VGND.t749 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4792 a_49212_26369# _397_.A2.t13 a_48988_26369# VPWR.t6500 pfet_06v0 ad=0.4599p pd=1.935u as=0.33945p ps=1.715u w=1.095u l=0.5u
X4793 VPWR.t3857 a_30364_1592# a_30276_1636# VPWR.t1700 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4794 VPWR.t5467 a_5388_13703# a_5300_13800# VPWR.t5466 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4795 VPWR.t1860 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t1859 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4796 VGND.t2057 _431_.A3 _444_.D VGND.t2056 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X4797 VGND.t4280 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t4279 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4798 VPWR.t2159 a_45416_29885# a_46772_29977# VPWR.t2158 pfet_06v0 ad=0.4554p pd=3.25u as=54f ps=0.66u w=0.36u l=0.5u
X4799 a_59036_1592# a_58948_1636# VGND.t752 VGND.t751 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4800 VGND.t6489 _287_.A1.t28 uo_out[6].t9 VGND.t6488 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4801 VPWR.t3613 a_54332_1592# a_54244_1636# VPWR.t2945 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4802 VPWR.t1166 a_15244_28248# a_15156_28292# VPWR.t1165 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4803 VPWR.t1959 _408_.ZN a_50704_27912# VPWR.t1958 pfet_06v0 ad=0.6588p pd=3.52u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4804 a_54444_23544# a_54356_23588# VGND.t552 VGND.t551 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4805 VPWR.t6021 a_1020_4728# a_932_4772# VPWR.t1757 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4806 a_63964_17272# a_63876_17316# VGND.t554 VGND.t553 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4807 a_4156_25112# a_4068_25156# VGND.t556 VGND.t555 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4808 VGND.t2474 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN VGND.t2473 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4809 a_43819_24372# _447_.Q.t12 _441_.A2 VGND.t6307 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4810 a_2364_19975# a_2276_20072# VGND.t558 VGND.t557 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4811 VGND.t424 a_30160_30301# a_30112_30345# VGND.t137 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X4812 a_13788_2727# a_13700_2824# VGND.t559 VGND.t377 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4813 a_37424_24463# a_35204_24455.t4 a_37179_24831# VGND.t6131 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4814 VPWR.t667 a_15244_25112# a_15156_25156# VPWR.t666 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4815 VPWR.t4878 a_47612_10567# a_47524_10664# VPWR.t1052 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4816 VPWR.t3126 a_1020_1592# a_932_1636# VPWR.t1507 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4817 a_34732_18407# a_34644_18504# VGND.t561 VGND.t560 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4818 a_52764_17272# a_52676_17316# VGND.t563 VGND.t562 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4819 a_4156_21976# a_4068_22020# VGND.t1911 VGND.t1365 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4820 VPWR.t4622 a_62172_18840# a_62084_18884# VPWR.t4621 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4821 VPWR.t3128 a_48060_1592# a_47972_1636# VPWR.t3127 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4822 a_31708_18407# a_31620_18504# VGND.t5650 VGND.t5649 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4823 VPWR.t6930 a_42392_22825.t32 _452_.CLK.t18 VPWR.t6929 pfet_06v0 ad=0.428p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4824 VPWR.t3814 a_62172_15704# a_62084_15748# VPWR.t940 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4825 VGND.t5651 a_14004_31048# uio_oe[2].t0 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4826 VPWR.t3480 _460_.Q _335_.ZN.t10 VPWR.t3479 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4827 VPWR.t1172 a_66428_14136# a_66340_14180# VPWR.t1171 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4828 VGND.t3329 _460_.Q a_34532_27208# VGND.t3328 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4829 _335_.ZN.t7 _334_.A1 a_35914_28776# VGND.t2240 nfet_06v0 ad=0.4161p pd=1.905u as=0.1517p ps=1.19u w=0.82u l=0.6u
X4830 VGND.t109 _294_.A2.t8 _288_.ZN.t2 VGND.t108 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4831 VPWR.t3981 a_45820_12568# a_45732_12612# VPWR.t3980 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4832 a_46848_20893# a_46476_20937# VGND.t1008 VGND.t1007 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X4833 VPWR.t2877 a_29692_21543# a_29604_21640# VPWR.t2876 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4834 VPWR.t473 a_66428_11000# a_66340_11044# VPWR.t472 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4835 VPWR.t996 a_67100_6296# a_67012_6340# VPWR.t995 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4836 a_58924_18840# a_58836_18884# VGND.t2141 VGND.t2140 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4837 _282_.ZN _398_.C VGND.t3154 VGND.t3153 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X4838 VPWR.t4574 a_50412_16839# a_50324_16936# VPWR.t4573 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4839 a_55676_27815# a_55588_27912# VGND.t5396 VGND.t5395 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4840 VPWR.t3378 a_67548_4295# a_67460_4392# VPWR.t3377 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4841 a_1020_13703# a_932_13800# VGND.t2007 VGND.t2006 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4842 a_54108_14136# a_54020_14180# VGND.t4010 VGND.t1371 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4843 VPWR.t5882 a_67100_3160# a_67012_3204# VPWR.t689 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4844 a_47724_18840# a_47636_18884# VGND.t4587 VGND.t4586 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4845 a_50196_22805# _395_.A2 _399_.A1 VGND.t5621 nfet_06v0 ad=0.2119p pd=1.335u as=0.4137p ps=1.9u w=0.815u l=0.6u
X4846 _397_.Z a_46984_23588# VPWR.t850 VPWR.t849 pfet_06v0 ad=0.5368p pd=3.32u as=0.389p ps=2.02u w=1.22u l=0.5u
X4847 a_4604_23544# a_4516_23588# VGND.t2009 VGND.t2008 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4848 a_44476_27815# a_44388_27912# VGND.t5220 VGND.t5219 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4849 a_24304_26795# a_23892_27208.t6 VGND.t6070 VGND.t6069 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4850 VGND.t5466 _328_.A2 _450_.D VGND.t5465 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X4851 a_43750_23544# a_44162_24120# a_44282_24164# VGND.t4836 nfet_06v0 ad=0.369p pd=2.77u as=43.2f ps=0.6u w=0.36u l=0.6u
X4852 VPWR.t89 uio_in[1].t0 a_50436_30689# VPWR.t88 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X4853 VPWR.t2116 a_67548_1159# a_67460_1256# VPWR.t2115 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4854 a_54108_11000# a_54020_11044# VGND.t5718 VGND.t5717 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4855 a_52997_20936# _419_.Z VGND.t4309 VGND.t4308 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4856 a_25744_30345# a_24864_29931# a_25420_30345# VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X4857 VGND.t4083 a_49600_30180# a_49496_30345# VGND.t137 nfet_06v0 ad=0.2637p pd=1.825u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4858 VPWR.t6579 _350_.A2.t26 _340_.A2 VPWR.t6578 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4859 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN VGND.t5409 VGND.t535 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4860 VGND.t4691 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN VGND.t4690 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4861 _324_.B.t13 _302_.Z VPWR.t4989 VPWR.t4988 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4862 a_4156_15704# a_4068_15748# VGND.t2014 VGND.t905 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4863 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t3059 VPWR.t3058 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4864 a_36188_25112# a_36100_25156# VGND.t1472 VGND.t907 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4865 _251_.A1.t3 a_63616_31128# VPWR.t6146 VPWR.t6145 pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X4866 a_2364_3160# a_2276_3204# VGND.t1473 VGND.t371 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4867 a_11100_1592# a_11012_1636# VGND.t1475 VGND.t1474 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4868 a_30812_15704# a_30724_15748# VGND.t1476 VGND.t909 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4869 clkload0.Z a_48384_26724# VPWR.t3002 VPWR.t3001 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4870 a_45456_30301.t0 _474_.CLK.t48 VPWR.t6759 VPWR.t6758 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X4871 a_57692_9432# a_57604_9476# VGND.t1478 VGND.t1477 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4872 a_49856_20936# _474_.Q a_49652_20936# VGND.t4650 nfet_06v0 ad=67.2f pd=0.74u as=88.2f ps=0.84u w=0.42u l=0.6u
X4873 a_44491_20936# _260_.A1 _260_.ZN VGND.t3770 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4874 hold1.Z a_44038_21236# VGND.t5981 VGND.t5980 nfet_06v0 ad=0.3608p pd=2.52u as=0.28262p ps=1.87u w=0.82u l=0.6u
X4875 a_25928_25273# a_24080_25227# a_25643_25273# VPWR.t4421 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X4876 VGND.t15 _397_.A1.t10 _412_.A1 VGND.t14 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X4877 a_14236_29816# a_14148_29860# VGND.t1479 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4878 a_34586_27912# _362_.B.t14 _290_.ZN VPWR.t6537 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4879 VPWR.t5071 a_56236_24679# a_56148_24776# VPWR.t5070 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4880 _402_.A1.t1 a_43736_25896# VPWR.t4112 VPWR.t4111 pfet_06v0 ad=0.3172p pd=1.74u as=0.854p ps=3.84u w=1.22u l=0.5u
X4881 a_43936_27165# a_43564_27209# VPWR.t4570 VPWR.t4569 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X4882 a_7068_29383# a_6980_29480# VGND.t5080 VGND.t5079 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4883 a_24900_27912# _455_.Q.t10 _351_.A2 VPWR.t6854 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4884 a_35616_24776# a_35204_24455.t5 VGND.t6133 VGND.t6132 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4885 a_61164_20408# a_61076_20452# VGND.t5176 VGND.t5175 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4886 VPWR.t3309 _398_.C a_51048_26680# VPWR.t3308 pfet_06v0 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X4887 VGND.t3680 a_43814_21236# a_44290_21236# VGND.t3679 nfet_06v0 ad=0.28262p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X4888 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv1.inv_array_notouch_\[1\].I VGND.t2632 VGND.t2631 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4889 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN VPWR.t4601 VPWR.t4600 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4890 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I VPWR.t2486 VPWR.t2485 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4891 VPWR.t5401 a_3708_30951# a_3620_31048# VPWR.t5400 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4892 a_52891_30644# a_52415_31220# a_52639_30644# VGND.t45 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X4893 VPWR.t4044 a_54444_26680# a_54356_26724# VPWR.t4043 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4894 _383_.ZN _397_.A1.t11 VGND.t17 VGND.t16 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4895 a_52428_13703# a_52340_13800# VGND.t1481 VGND.t1480 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4896 a_46794_25156# _398_.C _282_.ZN VPWR.t3307 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4897 VPWR.t2171 a_21740_29383# a_21652_29480# VPWR.t2170 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4898 a_11324_29383# a_11236_29480# VGND.t1382 VGND.t1381 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4899 a_12892_1592# a_12804_1636# VGND.t1482 VGND.t895 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4900 a_28460_23544# a_28372_23588# VGND.t1484 VGND.t1483 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4901 VPWR.t5421 a_54892_18407# a_54804_18504# VPWR.t5420 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4902 VPWR.t355 a_30476_25112# a_30388_25156# VPWR.t354 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4903 a_37980_17272# a_37892_17316# VGND.t1486 VGND.t1485 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4904 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I VPWR.t1487 VPWR.t1486 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4905 a_51618_22504# _476_.Q a_51414_22504# VGND.t4162 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4906 a_36860_1592# a_36772_1636# VGND.t1488 VGND.t1487 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4907 VPWR.t6976 _459_.Q.t15 _335_.ZN.t18 VPWR.t6975 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4908 a_40004_23233# _303_.ZN _441_.ZN VPWR.t2953 pfet_06v0 ad=0.58035p pd=2.155u as=0.4012p ps=1.85u w=1.095u l=0.5u
X4909 VPWR.t3711 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I VPWR.t3710 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4910 a_32144_26724# _294_.A2.t9 VPWR.t113 VPWR.t112 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4911 a_47388_15704# a_47300_15748# VGND.t1490 VGND.t1489 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4912 VPWR.t4232 _437_.ZN _441_.B VPWR.t4231 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4913 a_48956_12568# a_48868_12612# VGND.t1492 VGND.t1491 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4914 a_53772_26031# _412_.ZN a_52848_25987# VGND.t5091 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X4915 a_49600_30180# a_49112_29885# a_50032_30345# VGND.t137 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X4916 VGND.t6209 _459_.CLK.t34 a_26916_25640.t1 VGND.t6208 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X4917 a_41900_16839# a_41812_16936# VGND.t1494 VGND.t1493 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4918 a_61836_26680# a_61748_26724# VGND.t1778 VGND.t1777 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4919 a_42796_23981# a_43126_24119# a_43246_23610# VPWR.t3360 pfet_06v0 ad=0.3456p pd=2.64u as=61.19999f ps=0.7u w=0.36u l=0.5u
X4920 a_36188_15704# a_36100_15748# VGND.t1496 VGND.t1495 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4921 VGND.t4161 _476_.Q _424_.A1 VGND.t4160 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X4922 VGND.t3421 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I VGND.t3420 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4923 a_1916_28248# a_1828_28292# VGND.t4913 VGND.t1904 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4924 VPWR.t6043 a_19328_28733# a_19320_28409# VPWR.t6042 pfet_06v0 ad=0.2619p pd=1.685u as=50.4f ps=0.64u w=0.36u l=0.5u
X4925 VPWR.t755 a_4604_29816# a_4516_29860# VPWR.t754 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4926 VGND.t1425 _393_.A1 _393_.ZN VGND.t1424 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X4927 VPWR.t5687 a_13340_1159# a_13252_1256# VPWR.t512 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4928 VGND.t4278 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I VGND.t4277 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4929 VGND.t3747 vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN VGND.t3746 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4930 VPWR.t4086 _454_.Q _371_.A2 VPWR.t4085 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4931 a_54780_18840# a_54692_18884# VGND.t1970 VGND.t1969 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4932 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN VGND.t5897 VGND.t5896 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4933 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN VGND.t4455 VGND.t71 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4934 VPWR.t5524 a_4604_26680# a_4516_26724# VPWR.t5523 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4935 VPWR.t644 _386_.A4 a_47924_28292# VPWR.t643 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4936 VPWR.t4854 a_32604_16839# a_32516_16936# VPWR.t4764 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4937 a_17148_1159# a_17060_1256# VGND.t932 VGND.t931 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4938 VPWR.t5789 a_3260_13703# a_3172_13800# VPWR.t3756 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4939 VGND.t5665 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN VGND.t5664 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4940 VPWR.t4202 a_29184_25597# a_29176_25273# VPWR.t4201 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X4941 a_49448_20936# _419_.A4 VGND.t3984 VGND.t3983 nfet_06v0 ad=88.2f pd=0.84u as=0.226p ps=1.515u w=0.42u l=0.6u
X4942 a_44459_18559# a_42896_18504# a_43824_18147# VGND.t5733 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4943 clkbuf_1_0__f_clk.I.t23 a_44296_24393.t31 VGND.t283 VGND.t282 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X4944 VPWR.t5553 a_46848_20893# a_46820_20569# VPWR.t5552 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X4945 VPWR.t4388 a_25884_27815# a_25796_27912# VPWR.t4387 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4946 VGND.t3342 _267_.ZN _275_.A2 VGND.t3341 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X4947 a_11772_2727# a_11684_2824# VGND.t934 VGND.t933 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4948 a_37472_24419# a_37179_24831# VPWR.t1669 VPWR.t1668 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X4949 vgaringosc.workerclkbuff_notouch_.I.t1 _416_.A1.t10 a_51457_29861# VPWR.t203 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4950 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t2399 VPWR.t2398 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4951 VPWR.t6407 _337_.A3.t10 _337_.ZN VPWR.t6406 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4952 a_35740_2727# a_35652_2824# VGND.t2001 VGND.t2000 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4953 VPWR.t1738 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I VPWR.t1737 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4954 VPWR.t192 _424_.A2.t11 a_51988_24776# VPWR.t191 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4955 VPWR.t5181 a_65756_8999# a_65668_9096# VPWR.t989 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4956 VPWR.t453 a_54780_2727# a_54692_2824# VPWR.t452 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4957 a_39548_1592# a_39460_1636# VGND.t2002 VGND.t1085 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4958 a_58687_31220# a_58063_30644# a_58539_30644# VGND.t45 nfet_06v0 ad=0.369p pd=2.77u as=43.2f ps=0.6u w=0.36u l=0.6u
X4959 _379_.A2 uio_out[6].t11 VPWR.t6904 VPWR.t6903 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X4960 a_62503_28293# _250_.A2 _250_.ZN VPWR.t4851 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4961 a_1916_18840# a_1828_18884# VGND.t4157 VGND.t1088 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4962 VGND.t1928 _287_.A2 uo_out[6].t1 VGND.t1927 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4963 a_36076_16839# a_35988_16936# VGND.t2004 VGND.t2003 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4964 a_49034_21640# _324_.B.t32 _416_.A3 VPWR.t6715 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4965 a_54892_23544# a_54804_23588# VGND.t2005 VGND.t1090 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4966 a_42168_25640.t11 _284_.B a_43600_25640# VGND.t5391 nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4967 VPWR.t2621 a_15692_28248# a_15604_28292# VPWR.t2620 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4968 VPWR.t4358 a_65868_13703# a_65780_13800# VPWR.t4357 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4969 VPWR.t2252 a_24540_21543# a_24452_21640# VPWR.t2251 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4970 _260_.A2 _304_.B VGND.t4533 VGND.t4532 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X4971 a_50276_27912# _330_.A1.t18 VPWR.t218 VPWR.t217 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4972 VPWR.t4973 a_4604_17272# a_4516_17316# VPWR.t4972 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4973 a_42168_22504# _302_.Z a_43600_22504# VGND.t4844 nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4974 VPWR.t3692 a_28572_1592# a_28484_1636# VPWR.t3691 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4975 VPWR.t4362 a_54668_13703# a_54580_13800# VPWR.t4361 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4976 VPWR.t4974 a_15692_25112# a_15604_25156# VPWR.t2991 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4977 VPWR.t3695 a_5500_1592# a_5412_1636# VPWR.t3694 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4978 a_53212_1159# a_53124_1256# VGND.t4585 VGND.t4584 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4979 a_51988_24072# _399_.ZN a_51332_24072# VGND.t1186 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4980 VPWR.t6247 a_36636_26680# a_36548_26724# VPWR.t1573 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4981 a_48272_25156.t2 clkbuf_1_0__f_clk.I.t51 VPWR.t264 VPWR.t263 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X4982 VPWR.t4976 a_55228_9432# a_55140_9476# VPWR.t4975 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4983 a_37584_29123# a_37291_29535# VGND.t665 VGND.t664 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X4984 VPWR.t1548 a_14236_29816# a_14148_29860# VPWR.t1547 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4985 VPWR.t5111 a_59708_23111# a_59620_23208# VPWR.t5110 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4986 VGND.t4332 vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I VGND.t4331 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X4987 a_30795_29977# a_29232_29931# a_30160_30301# VGND.t137 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4988 a_57132_10567# a_57044_10664# VGND.t1996 VGND.t1995 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4989 a_18828_23544# a_18740_23588# VGND.t1998 VGND.t1997 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4990 VPWR.t6080 a_35292_1159# a_35204_1256# VPWR.t6079 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4991 a_61276_1592# a_61188_1636# VGND.t1999 VGND.t956 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4992 VPWR.t605 a_66876_14136# a_66788_14180# VPWR.t604 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4993 _434_.ZN _301_.A1 a_38529_22804# VGND.t3201 nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X4994 a_35000_22137# a_33152_22091# a_34715_22137# VPWR.t1469 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X4995 VPWR.t2558 _349_.A4 _371_.A2 VPWR.t2557 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4996 a_18716_30951# a_18628_31048# VGND.t1982 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4997 VPWR.t3989 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I VPWR.t3988 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X4998 VPWR.t1250 a_66876_11000# a_66788_11044# VPWR.t1249 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4999 VPWR.t5502 a_7964_2727# a_7876_2824# VPWR.t5501 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5000 a_43284_18191# a_42484_18183.t4 VGND.t6731 VGND.t6730 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5001 VGND.t6370 _452_.CLK.t49 a_42484_18183.t1 VGND.t6369 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X5002 a_37408_23208# _447_.Q.t13 VPWR.t6588 VPWR.t6587 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5003 VPWR.t5504 a_50860_16839# a_50772_16936# VPWR.t5503 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5004 VPWR.t5314 a_4940_7431# a_4852_7528# VPWR.t5313 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5005 a_54556_14136# a_54468_14180# VGND.t5560 VGND.t960 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5006 VGND.t81 uio_in[1].t1 a_50436_30689# VGND.t80 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5007 VPWR.t3332 a_52092_15271# a_52004_15368# VPWR.t3331 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5008 a_54556_11000# a_54468_11044# VGND.t2326 VGND.t2325 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5009 VPWR.t5167 a_38428_15271# a_38340_15368# VPWR.t5166 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5010 VGND.t166 _336_.A2.t8 a_29028_24072# VGND.t165 nfet_06v0 ad=0.23405p pd=1.555u as=58.39999f ps=0.685u w=0.365u l=0.6u
X5011 VPWR.t5061 a_57244_12568# a_57156_12612# VPWR.t5060 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5012 VPWR.t185 _384_.A3.t16 a_49828_22020# VPWR.t184 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5013 a_35108_28776# _460_.Q a_34084_28776# VGND.t3327 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5014 a_38428_2727# a_38340_2824# VGND.t1984 VGND.t1983 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5015 a_20191_29611# uio_out[5].t12 a_20003_29611# VPWR.t6900 pfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.5u
X5016 VPWR.t2355 _334_.A1 a_35008_27533# VPWR.t2354 pfet_06v0 ad=0.34437p pd=1.895u as=0.1456p ps=1.08u w=0.56u l=0.5u
X5017 VPWR.t2609 _275_.ZN a_51457_29861# VPWR.t2608 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X5018 clkbuf_1_0__f_clk.I.t6 a_44296_24393.t32 VPWR.t286 VPWR.t285 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5019 a_43824_18147# a_43452_18191# VPWR.t57 VPWR.t56 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X5020 VGND.t203 _416_.A1.t11 _475_.D VGND.t202 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X5021 VPWR.t4208 _336_.A1 _337_.ZN VPWR.t4207 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5022 a_33948_18840# a_33860_18884# VGND.t1979 VGND.t1883 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5023 VPWR.t3984 a_53704_23219# a_55060_23263# VPWR.t3983 pfet_06v0 ad=0.4554p pd=3.25u as=54f ps=0.66u w=0.36u l=0.5u
X5024 VPWR.t3063 a_47836_17272# a_47748_17316# VPWR.t3062 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5025 a_1916_30951# a_1828_31048# VGND.t648 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5026 VPWR.t4373 a_57468_2727# a_57380_2824# VPWR.t4372 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5027 VPWR.t3445 a_4156_5863# a_4068_5960# VPWR.t2582 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5028 a_41642_25156# _304_.B _260_.A2 VPWR.t4687 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5029 a_14684_29816# a_14596_29860# VGND.t649 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5030 a_46389_21236# _419_.A4 VGND.t3982 VGND.t3981 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5031 VPWR.t593 a_36636_17272# a_36548_17316# VPWR.t592 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5032 _248_.B1 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I VPWR.t4380 VPWR.t4379 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5033 VPWR.t4294 a_4156_2727# a_4068_2824# VPWR.t4130 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5034 VPWR.t3905 a_56796_1592# a_56708_1636# VPWR.t3904 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5035 a_1468_26247# a_1380_26344# VGND.t651 VGND.t650 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5036 a_1916_7864# a_1828_7908# VGND.t653 VGND.t652 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5037 a_66204_17272# a_66116_17316# VGND.t655 VGND.t654 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5038 a_8188_1592# a_8100_1636# VGND.t657 VGND.t656 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5039 a_29468_1159# a_29380_1256# VGND.t2554 VGND.t2553 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5040 a_39772_20408# a_39684_20452# VGND.t1411 VGND.t1410 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5041 a_18716_24679# a_18628_24776# VGND.t659 VGND.t658 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5042 a_42236_15704# a_42148_15748# VGND.t415 VGND.t414 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5043 a_1468_23111# a_1380_23208# VGND.t417 VGND.t416 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5044 a_29176_25273# a_27328_25227# a_28891_25273# VPWR.t6291 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X5045 a_1916_4728# a_1828_4772# VGND.t5765 VGND.t2142 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5046 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN VPWR.t4599 VPWR.t4598 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5047 a_32380_21543# a_32292_21640# VGND.t3588 VGND.t3587 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5048 a_18716_21543# a_18628_21640# VGND.t3346 VGND.t3345 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5049 VPWR.t5948 a_26668_20408# a_26580_20452# VPWR.t5947 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5050 VPWR.t5516 a_54892_26680# a_54804_26724# VPWR.t5515 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5051 a_37516_27599# _443_.D a_37392_27967# VPWR.t4039 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X5052 a_52876_13703# a_52788_13800# VGND.t419 VGND.t418 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5053 a_35008_22461# a_34715_22137# VPWR.t2241 VPWR.t2240 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X5054 a_35088_20893# a_34716_20937# VGND.t3859 VGND.t3858 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X5055 _345_.A2 _454_.Q VGND.t3938 VGND.t3937 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X5056 VPWR.t382 a_17932_21543# a_17844_21640# VPWR.t381 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5057 a_11772_29383# a_11684_29480# VGND.t4048 VGND.t4047 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5058 a_25548_20408# a_25460_20452# VGND.t1435 VGND.t1434 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5059 a_51956_26183# a_52400_25987.t5 a_52352_26031# VGND.t6098 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X5060 a_51968_26724# _395_.A2 VPWR.t5847 VPWR.t5846 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5061 a_4940_24679# a_4852_24776# VGND.t421 VGND.t420 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5062 a_25124_28776# _454_.Q a_25740_28776# VGND.t3936 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5063 _371_.A2 _337_.A3.t11 a_26954_28776# VGND.t6141 nfet_06v0 ad=0.4161p pd=1.905u as=0.1517p ps=1.19u w=0.82u l=0.6u
X5064 VPWR.t1203 _290_.ZN a_33508_31048# VPWR.t1202 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5065 a_22992_27555# a_22620_27599# VPWR.t4252 VPWR.t4251 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X5066 a_4940_21543# a_4852_21640# VGND.t1748 VGND.t1747 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5067 VPWR.t2843 a_59260_23544# a_59172_23588# VPWR.t2497 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5068 a_1916_24679# a_1828_24776# VGND.t2282 VGND.t2281 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5069 a_16700_29816# a_16612_29860# VGND.t2283 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5070 a_46596_20127# a_45284_19751.t3 a_46252_19759# VPWR.t7031 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X5071 a_21268_27912# _455_.Q.t11 _346_.ZN VPWR.t6855 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X5072 a_5052_9432# a_4964_9476# VGND.t2285 VGND.t2284 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5073 VPWR.t194 _424_.A2.t12 a_52884_18884# VPWR.t193 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5074 a_61164_10567# a_61076_10664# VGND.t2287 VGND.t2286 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5075 a_19328_28733# a_19035_28409# VPWR.t3670 VPWR.t3669 pfet_06v0 ad=0.2457p pd=1.465u as=0.2619p ps=1.685u w=0.945u l=0.5u
X5076 a_1916_21543# a_1828_21640# VGND.t4001 VGND.t1314 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5077 VPWR.t3388 a_56236_23544# a_56148_23588# VPWR.t3387 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5078 a_9532_29383# a_9444_29480# VGND.t3220 VGND.t3219 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5079 a_5052_6296# a_4964_6340# VGND.t5339 VGND.t5338 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5080 a_43804_1592# a_43716_1636# VGND.t2288 VGND.t809 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5081 a_64524_16839# a_64436_16936# VGND.t2290 VGND.t2289 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5082 VPWR.t2926 a_41788_15704# a_41700_15748# VPWR.t2925 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5083 a_1468_16839# a_1380_16936# VGND.t2291 VGND.t1169 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5084 VGND.t3685 _255_.I _255_.ZN VGND.t3684 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X5085 a_24428_21976# a_24340_22020# VGND.t2319 VGND.t2318 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5086 a_37291_29535# a_35316_29159.t3 a_36656_29123# VPWR.t7054 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X5087 VPWR.t559 a_2364_19975# a_2276_20072# VPWR.t316 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5088 a_44571_26841# a_42596_27208.t5 a_43936_27165# VPWR.t141 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X5089 VPWR.t4867 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN VPWR.t4866 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5090 VPWR.t4769 a_58252_16839# a_58164_16936# VPWR.t4768 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5091 a_57020_1159# a_56932_1256# VGND.t4768 VGND.t4767 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5092 a_11548_30951# a_11460_31048# VGND.t2495 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5093 VPWR.t5263 a_5724_29383# a_5636_29480# VPWR.t5262 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5094 VGND.t4969 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN VGND.t4968 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5095 a_37360_19325# a_37067_19001# VGND.t1265 VGND.t1264 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X5096 a_7068_2727# a_6980_2824# VGND.t2497 VGND.t2496 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5097 VPWR.t4519 a_47052_16839# a_46964_16936# VPWR.t4518 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5098 VPWR.t6180 a_60716_13703# a_60628_13800# VPWR.t6179 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5099 VGND.t914 _384_.A1 _398_.C VGND.t913 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5100 VGND.t6339 _350_.A1.t9 _373_.A2 VGND.t102 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X5101 a_23834_28292# _454_.Q _345_.A2 VPWR.t4084 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5102 a_47802_26724# _412_.A1 _419_.A4 VPWR.t3839 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5103 VPWR.t6106 a_51868_17272# a_51780_17316# VPWR.t6105 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5104 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN VPWR.t4722 VPWR.t4721 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5105 _304_.B a_54432_31128# VPWR.t4672 VPWR.t4671 pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X5106 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t4276 VGND.t4275 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5107 a_38652_15704# a_38564_15748# VGND.t2499 VGND.t2498 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5108 _304_.A1.t1 a_35232_24029# VGND.t5473 VGND.t5472 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5109 VPWR.t5324 a_57132_18407# a_57044_18504# VPWR.t5323 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5110 a_52204_18407# a_52116_18504# VGND.t2501 VGND.t2500 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5111 a_35216_27533# _363_.Z.t5 a_35008_27533# VGND.t36 nfet_06v0 ad=57.59999f pd=0.68u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5112 VPWR.t5325 a_65308_18407# a_65220_18504# VPWR.t3056 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5113 VPWR.t659 a_1916_7864# a_1828_7908# VPWR.t2 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5114 VPWR.t5579 a_32604_18840# a_32516_18884# VPWR.t1253 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5115 a_22748_24679# a_22660_24776# VGND.t2293 VGND.t2292 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5116 VPWR.t4257 a_32604_15704# a_32516_15748# VPWR.t3951 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5117 _459_.CLK.t11 a_41048_29816.t15 VGND.t6405 VGND.t6400 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X5118 VPWR.t5053 a_3260_12568# a_3172_12612# VPWR.t2390 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5119 a_16140_26247# a_16052_26344# VGND.t2295 VGND.t2294 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5120 _459_.CLK.t3 a_41048_29816.t16 VPWR.t6691 VPWR.t6690 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5121 a_45696_20072# a_45284_19751.t4 VPWR.t7033 VPWR.t7032 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X5122 a_22748_21543# a_22660_21640# VGND.t1707 VGND.t1706 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5123 a_24316_26247# a_24228_26344# VGND.t2297 VGND.t2296 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5124 VPWR.t4218 a_5388_5863# a_5300_5960# VPWR.t4217 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5125 a_47836_15271# a_47748_15368# VGND.t2299 VGND.t2298 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5126 a_16140_23111# a_16052_23208# VGND.t2301 VGND.t2300 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5127 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN VGND.t5722 VGND.t5721 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5128 a_17932_27815# a_17844_27912# VGND.t3263 VGND.t3262 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5129 a_12444_2727# a_12356_2824# VGND.t2302 VGND.t549 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5130 VPWR.t656 a_14684_29816# a_14596_29860# VPWR.t655 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5131 a_45456_30301.t1 _474_.CLK.t49 VGND.t6459 VGND.t139 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X5132 a_57580_10567# a_57492_10664# VGND.t2304 VGND.t2303 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5133 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN VPWR.t6130 VPWR.t6129 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5134 VPWR.t4533 a_2364_7431# a_2276_7528# VPWR.t791 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5135 VPWR.t4536 a_31484_2727# a_31396_2824# VPWR.t4535 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5136 VGND.t1934 a_39268_18840# a_38644_19368# VGND.t1933 nfet_06v0 ad=0.218p pd=1.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5137 VPWR.t5226 a_11548_1592# a_11460_1636# VPWR.t5225 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5138 VGND.t3437 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t3436 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5139 a_66092_19975# a_66004_20072# VGND.t1018 VGND.t1017 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5140 _327_.A2 a_44752_18147# VPWR.t4172 VPWR.t4171 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5141 VGND.t4498 a_36656_29123# a_36608_29167# VGND.t4497 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X5142 VPWR.t5228 a_35516_1592# a_35428_1636# VPWR.t5227 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5143 VPWR.t3897 a_43400_18909# a_44756_19001# VPWR.t3896 pfet_06v0 ad=0.4554p pd=3.25u as=54f ps=0.66u w=0.36u l=0.5u
X5144 _427_.A2 _324_.C.t26 VPWR.t6807 VPWR.t6806 pfet_06v0 ad=0.44325p pd=2.87u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5145 VPWR.t3478 _460_.Q a_35140_26680# VPWR.t3477 pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X5146 a_49740_16839# a_49652_16936# VGND.t1020 VGND.t1019 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5147 a_36172_24463# _444_.D a_36048_24831# VPWR.t5641 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X5148 a_1020_17272# a_932_17316# VGND.t1021 VGND.t61 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5149 a_63068_19975# a_62980_20072# VGND.t1023 VGND.t1022 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5150 a_59484_1592# a_59396_1636# VGND.t1025 VGND.t1024 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5151 VPWR.t5474 a_54780_1592# a_54692_1636# VPWR.t2936 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5152 VPWR.t5381 a_26556_23111# a_26468_23208# VPWR.t5380 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5153 VPWR.t3151 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN VPWR.t3150 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5154 a_45920_20523# a_45508_20936.t6 VGND.t192 VGND.t191 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X5155 VGND.t5782 a_41188_18840# _327_.Z VGND.t5781 nfet_06v0 ad=0.2424p pd=1.635u as=0.341p ps=2.43u w=0.775u l=0.6u
X5156 VPWR.t2780 a_66204_4295# a_66116_4392# VPWR.t891 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5157 VPWR.t5383 a_38876_15271# a_38788_15368# VPWR.t5382 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5158 a_2364_29383# a_2276_29480# VGND.t1824 VGND.t1823 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5159 VPWR.t2243 a_42236_1159# a_42148_1256# VPWR.t2242 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5160 VPWR.t6110 a_57692_12568# a_57604_12612# VPWR.t6109 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5161 _351_.A2 _455_.Q.t12 a_25108_27508# VGND.t6538 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5162 VPWR.t4846 a_62284_16839# a_62196_16936# VPWR.t4845 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5163 VGND.t6065 _288_.ZN.t8 uo_out[2].t10 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X5164 VPWR.t4553 a_66204_1159# a_66116_1256# VPWR.t4552 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5165 VPWR.t3010 a_32716_20408# a_32628_20452# VPWR.t3009 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5166 a_26556_28776# _349_.A4 VGND.t2431 VGND.t2430 nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5167 clkbuf_1_0__f_clk.I.t5 a_44296_24393.t33 VPWR.t288 VPWR.t287 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5168 a_25184_27209# a_24304_26795# a_24860_27209# VGND.t1099 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X5169 a_21044_27508# _346_.B VGND.t400 VGND.t399 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5170 VPWR.t2404 a_16700_29816# a_16612_29860# VPWR.t2403 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5171 a_34939_23705# a_32964_24072.t7 a_34304_24029# VPWR.t156 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X5172 VPWR.t5924 _293_.A2 a_40644_29480# VPWR.t5923 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5173 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I VPWR.t5908 VPWR.t5907 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5174 VGND.t6211 _459_.CLK.t35 a_35316_29159.t1 VGND.t6210 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X5175 VPWR.t5602 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN VPWR.t5601 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5176 VPWR.t3079 a_47164_12135# a_47076_12232# VPWR.t1335 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5177 a_1020_3160# a_932_3204# VGND.t321 VGND.t320 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5178 VPWR.t1092 a_8636_2727# a_8548_2824# VPWR.t1091 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5179 a_42392_22825.t8 clkbuf_1_0__f_clk.I.t52 VGND.t263 VGND.t262 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X5180 a_57132_23544# a_57044_23588# VGND.t4871 VGND.t4870 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5181 VPWR.t5163 a_68108_13703# a_68020_13800# VPWR.t5162 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5182 a_66652_17272# a_66564_17316# VGND.t4873 VGND.t4872 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5183 VPWR.t5675 a_35232_24029# a_35224_23705# VPWR.t5674 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X5184 _350_.A2.t1 _223_.ZN VPWR.t796 VPWR.t795 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5185 VPWR.t5152 a_61612_23111# a_61524_23208# VPWR.t5151 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5186 _337_.ZN _336_.A1 a_28756_25940# VGND.t4054 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5187 uo_out[0].t0 _296_.ZN VGND.t3513 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X5188 a_61948_26247# a_61860_26344# VGND.t4875 VGND.t4874 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5189 a_42684_15704# a_42596_15748# VGND.t4877 VGND.t4876 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5190 a_64636_2727# a_64548_2824# VGND.t4878 VGND.t1053 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5191 a_36016_20893# a_35723_20569# VGND.t3893 VGND.t3892 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X5192 VPWR.t4489 a_67996_1159# a_67908_1256# VPWR.t4488 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5193 VGND.t1291 a_22560_30288# uio_out[4].t1 VGND.t71 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5194 a_37840_27599# a_36960_27912# a_37516_27599# VGND.t5298 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X5195 a_45820_14136# a_45732_14180# VGND.t3069 VGND.t3068 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5196 VPWR.t3943 a_54824_22045# a_56180_22137# VPWR.t3942 pfet_06v0 ad=0.4554p pd=3.25u as=54f ps=0.66u w=0.36u l=0.5u
X5197 a_67100_7864# a_67012_7908# VGND.t4880 VGND.t4879 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5198 a_66428_12568# a_66340_12612# VGND.t4882 VGND.t4881 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5199 a_33052_17272# a_32964_17316# VGND.t4884 VGND.t4883 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5200 a_44296_24393.t9 clk.t9 VGND.t6531 VGND.t6530 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X5201 a_45820_11000# a_45732_11044# VGND.t3038 VGND.t3037 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5202 VPWR.t3183 a_35140_26680# _363_.Z.t0 VPWR.t3182 pfet_06v0 ad=0.4268p pd=2.175u as=0.5346p ps=3.31u w=1.215u l=0.5u
X5203 VGND.t3529 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN VGND.t3528 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5204 a_67100_4728# a_67012_4772# VGND.t3899 VGND.t3385 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5205 a_14796_20408# a_14708_20452# VGND.t3781 VGND.t1578 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5206 a_33708_22505# _316_.ZN a_33540_22505# VGND.t5286 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X5207 VPWR.t4664 a_53100_16839# a_53012_16936# VPWR.t4663 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5208 VPWR.t6660 _452_.CLK.t50 a_32964_24072.t0 VPWR.t6659 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X5209 VPWR.t3055 a_51196_21543# a_51108_21640# VPWR.t3054 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5210 VPWR.t3442 a_4156_4728# a_4068_4772# VPWR.t1377 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5211 VPWR.t6025 a_65756_27815# a_65668_27912# VPWR.t6024 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5212 _274_.A3 _268_.A1.t7 a_52640_29860# VPWR.t6738 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X5213 a_40668_15271# a_40580_15368# VGND.t4888 VGND.t4887 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5214 VPWR.t5430 a_48060_30951# a_47972_31048# VPWR.t5429 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5215 a_36188_1159# a_36100_1256# VGND.t616 VGND.t615 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5216 VPWR.t5801 a_56684_23544# a_56596_23588# VPWR.t5800 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5217 a_9980_29383# a_9892_29480# VGND.t6021 VGND.t6020 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5218 VPWR.t5802 a_4156_1592# a_4068_1636# VPWR.t4249 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5219 _340_.ZN _349_.A4 VGND.t2429 VGND.t2428 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X5220 VPWR.t2604 vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN VPWR.t1710 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5221 VPWR.t1341 a_64188_1159# a_64100_1256# VPWR.t1009 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5222 VGND.t134 _417_.A2.t10 a_51240_23340# VGND.t133 nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X5223 a_65308_9432# a_65220_9476# VGND.t1277 VGND.t1276 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5224 a_64972_16839# a_64884_16936# VGND.t1279 VGND.t1278 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5225 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN VPWR.t4061 VPWR.t4060 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5226 a_56236_22505# _427_.ZN a_55312_22340# VGND.t3639 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X5227 a_26148_28776# _454_.Q a_25124_28776# VGND.t3935 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5228 a_24876_21976# a_24788_22020# VGND.t3360 VGND.t3359 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5229 VPWR.t2384 a_14796_21976# a_14708_22020# VPWR.t1657 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5230 a_33500_15704# a_33412_15748# VGND.t1280 VGND.t404 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5231 VPWR.t6263 a_39264_18147# a_39256_18559# VPWR.t6262 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X5232 a_65308_6296# a_65220_6340# VGND.t2948 VGND.t2947 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5233 VPWR.t6703 vgaringosc.workerclkbuff_notouch_.I.t8 a_41048_29816.t1 VPWR.t6702 pfet_06v0 ad=0.3608p pd=2.52u as=0.2952p ps=1.54u w=0.82u l=0.5u
X5234 VPWR.t4936 a_30588_23111# a_30500_23208# VPWR.t4935 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5235 VPWR.t3159 a_45904_30180# a_45800_30345# VPWR.t3158 pfet_06v0 ad=0.1044p pd=0.94u as=0.1791p ps=1.355u w=0.36u l=0.5u
X5236 VPWR.t5781 a_23084_23544# a_22996_23588# VPWR.t5780 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5237 a_59036_9432# a_58948_9476# VGND.t1282 VGND.t1281 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5238 a_42572_16839# a_42484_16936# VGND.t1284 VGND.t1283 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5239 VPWR.t3528 a_17932_20408# a_17844_20452# VPWR.t3527 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5240 a_48708_29816# a_49112_29885# a_49056_29977# VPWR.t2337 pfet_06v0 ad=0.1665p pd=1.285u as=50.4f ps=0.64u w=0.36u l=0.5u
X5241 a_26720_30301# a_26427_29977# VGND.t5061 VGND.t2052 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X5242 VGND.t2995 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I VGND.t2994 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5243 VPWR.t2332 _316_.A3 a_35268_21640# VPWR.t2331 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5244 a_40416_27209# a_39536_26795# a_40092_27209# VGND.t3118 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X5245 VPWR.t4412 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN VPWR.t4411 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5246 _350_.A2.t19 _335_.ZN.t26 VPWR.t7003 VPWR.t7002 pfet_06v0 ad=0.2561p pd=1.505u as=0.3766p ps=1.815u w=0.985u l=0.5u
X5247 _416_.A1.t1 _324_.C.t27 VPWR.t6809 VPWR.t6808 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5248 _448_.D _325_.A2.t8 VGND.t6124 VGND.t6123 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5249 VGND.t3861 a_35088_20893# a_35040_20937# VGND.t3860 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X5250 a_66316_13703# a_66228_13800# VGND.t1199 VGND.t1198 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5251 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN VGND.t3990 VGND.t3989 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5252 VPWR.t730 _427_.A2 a_53108_21640# VPWR.t729 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5253 VGND.t6284 a_48272_25156.t37 _474_.CLK.t23 VGND.t6283 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5254 _409_.ZN _330_.A1.t19 a_50068_27508# VGND.t218 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5255 a_22059_26399# a_20084_26023.t6 a_21424_25987# VPWR.t7005 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X5256 a_55116_13703# a_55028_13800# VGND.t1201 VGND.t1200 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5257 VPWR.t3121 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN VPWR.t3120 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5258 a_44906_23588# a_44786_24120# a_44162_24120# VPWR.t1787 pfet_06v0 ad=61.19999f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X5259 a_52652_18407# a_52564_18504# VGND.t1203 VGND.t1202 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5260 VPWR.t4927 a_57580_18407# a_57492_18504# VPWR.t4926 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5261 a_23627_27967# a_21652_27591.t7 a_22992_27555# VPWR.t105 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X5262 a_63740_1592# a_63652_1636# VGND.t1205 VGND.t1204 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5263 a_40416_18885# _452_.Q.t15 VPWR.t6961 VPWR.t6960 pfet_06v0 ad=0.44955p pd=1.955u as=0.5346p ps=3.31u w=1.215u l=0.5u
X5264 a_14236_1592# a_14148_1636# VGND.t1207 VGND.t1206 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5265 VPWR.t2336 a_49112_29885# a_50468_29977# VPWR.t2335 pfet_06v0 ad=0.4554p pd=3.25u as=54f ps=0.66u w=0.36u l=0.5u
X5266 a_28596_27916.t8 _350_.A1.t10 _352_.A2.t8 VPWR.t6626 pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X5267 VPWR.t5078 a_64412_8999# a_64324_9096# VPWR.t5077 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5268 a_16700_1159# a_16612_1256# VGND.t3466 VGND.t3465 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5269 VPWR.t4930 a_62508_10567# a_62420_10664# VPWR.t4929 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5270 a_38204_1592# a_38116_1636# VGND.t634 VGND.t633 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5271 VPWR.t5192 a_36300_23544# a_36212_23588# VPWR.t5191 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5272 a_26427_29977# a_24864_29931# a_25792_30301# VGND.t137 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X5273 a_46198_27060# _424_.A2.t13 VGND.t188 VGND.t187 nfet_06v0 ad=0.3608p pd=2.52u as=0.2911p ps=1.53u w=0.82u l=0.6u
X5274 _459_.CLK.t10 a_41048_29816.t17 VGND.t6406 VGND.t6400 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X5275 _313_.ZN _330_.A1.t20 VGND.t220 VGND.t219 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5276 _459_.CLK.t2 a_41048_29816.t18 VPWR.t6693 VPWR.t6692 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5277 VPWR.t4303 a_35180_18407# a_35092_18504# VPWR.t4302 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5278 _474_.Q a_48888_19243# VPWR.t2893 VPWR.t2892 pfet_06v0 ad=0.3172p pd=1.74u as=0.854p ps=3.84u w=1.22u l=0.5u
X5279 VPWR.t2703 _319_.A3 a_35716_20072# VPWR.t2702 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5280 VGND.t3836 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I VGND.t3835 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5281 VPWR.t5310 a_44924_15271# a_44836_15368# VPWR.t3640 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5282 _448_.Q.t1 a_37360_19325# VGND.t5501 VGND.t5500 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5283 a_1468_26680# a_1380_26724# VGND.t5932 VGND.t5798 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5284 VPWR.t3816 a_63740_12568# a_63652_12612# VPWR.t3815 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5285 VPWR.t5415 a_21404_23111# a_21316_23208# VPWR.t5414 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5286 a_4604_28248# a_4516_28292# VGND.t1238 VGND.t1237 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5287 VPWR.t5035 a_67100_7864# a_67012_7908# VPWR.t5034 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5288 VPWR.t5407 a_55228_15704# a_55140_15748# VPWR.t5406 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5289 a_63616_31128# ui_in[0].t2 VGND.t6736 VGND.t80 nfet_06v0 ad=0.51425p pd=2.91u as=0.2662p ps=2.09u w=0.605u l=0.6u
X5290 _411_.A2.t3 _397_.A2.t14 a_48580_27508# VGND.t6226 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5291 VPWR.t4444 a_32156_18407# a_32068_18504# VPWR.t4443 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5292 VPWR.t3818 a_52540_12568# a_52452_12612# VPWR.t3817 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5293 VPWR.t507 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I VPWR.t506 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5294 VPWR.t4356 a_44028_15704# a_43940_15748# VPWR.t3703 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5295 a_62396_27815# a_62308_27912# VGND.t1737 VGND.t1736 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5296 VGND.t6150 _451_.Q.t7 a_38548_21327# VGND.t6149 nfet_06v0 ad=0.23405p pd=1.555u as=58.39999f ps=0.685u w=0.365u l=0.6u
X5297 _267_.ZN _267_.A1 VPWR.t5818 VPWR.t5817 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X5298 VPWR.t4624 a_59932_2727# a_59844_2824# VPWR.t4623 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5299 a_2812_18407# a_2724_18504# VGND.t355 VGND.t354 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5300 _334_.A1 a_37584_29123# VGND.t1948 VGND.t1947 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5301 a_43253_25940# _451_.Q.t8 VGND.t6152 VGND.t6151 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5302 _352_.A2.t6 _371_.A2 VGND.t3431 VGND.t3430 nfet_06v0 ad=0.1326p pd=1.03u as=0.1326p ps=1.03u w=0.51u l=0.6u
X5303 VPWR.t3794 a_61948_9432# a_61860_9476# VPWR.t3793 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5304 a_4940_4295# a_4852_4392# VGND.t2060 VGND.t2059 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5305 VPWR.t3796 a_57132_17272# a_57044_17316# VPWR.t3795 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5306 VPWR.t4733 a_6620_2727# a_6532_2824# VPWR.t4732 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5307 VPWR.t4122 a_65308_17272# a_65220_17316# VPWR.t4121 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5308 VPWR.t368 a_22748_1159# a_22660_1256# VPWR.t367 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5309 VGND.t3597 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN VGND.t3596 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5310 a_61500_17272# a_61412_17316# VGND.t359 VGND.t358 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5311 VPWR.t2069 a_46716_1159# a_46628_1256# VPWR.t2068 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5312 VPWR.t4078 a_55676_9432# a_55588_9476# VPWR.t4077 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5313 a_28012_24679# a_27924_24776# VGND.t361 VGND.t360 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5314 a_3260_7431# a_3172_7528# VGND.t363 VGND.t362 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5315 a_7740_29816# a_7652_29860# VGND.t364 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5316 a_66428_1592# a_66340_1636# VGND.t366 VGND.t365 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5317 VPWR.t4275 a_37868_16839# a_37780_16936# VPWR.t4274 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5318 a_32380_2727# a_32292_2824# VGND.t368 VGND.t367 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5319 a_40644_31048# _284_.ZN.t32 uo_out[0].t7 VPWR.t6521 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X5320 VPWR.t4001 a_2364_9432# a_2276_9476# VPWR.t4000 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5321 VPWR.t4784 a_61724_1592# a_61636_1636# VPWR.t4783 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5322 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I VGND.t3435 VGND.t3434 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5323 VPWR.t1221 a_8627_30644# uio_oe[6].t0 VPWR.t1220 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5324 a_20844_20408# a_20756_20452# VGND.t2750 VGND.t2749 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5325 a_40196_29480# _293_.A2 VPWR.t5922 VPWR.t5921 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X5326 VGND.t1421 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN VGND.t1420 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5327 a_4604_18840# a_4516_18884# VGND.t2226 VGND.t2225 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5328 VPWR.t4453 a_56124_2727# a_56036_2824# VPWR.t4452 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5329 a_57580_23544# a_57492_23588# VGND.t1152 VGND.t1151 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5330 VPWR.t2379 _226_.ZN a_41488_24072# VPWR.t2378 pfet_06v0 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X5331 a_48508_13703# a_48420_13800# VGND.t1153 VGND.t579 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5332 a_39256_18559# a_37408_18504# a_38971_18559# VPWR.t1846 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X5333 a_53212_27815# a_53124_27912# VGND.t3609 VGND.t3608 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5334 VPWR.t2794 a_18380_25112# a_18292_25156# VPWR.t2793 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5335 a_45820_10567# a_45732_10664# VGND.t1155 VGND.t1154 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5336 VPWR.t4459 a_58924_10567# a_58836_10664# VPWR.t4458 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5337 VPWR.t2902 a_60604_27815# a_60516_27912# VPWR.t2901 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5338 VPWR.t6811 _324_.C.t28 _424_.A2.t2 VPWR.t6810 pfet_06v0 ad=0.2938p pd=1.65u as=0.2938p ps=1.65u w=1.13u l=0.5u
X5339 _346_.ZN _455_.Q.t13 a_21044_27508# VGND.t6539 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5340 a_38759_24072# _437_.ZN a_38575_24072# VGND.t4073 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5341 vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN VGND.t2688 VGND.t2687 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5342 VPWR.t1883 a_28124_26680# a_28036_26724# VPWR.t1882 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5343 a_66876_12568# a_66788_12612# VGND.t1157 VGND.t1156 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5344 a_30924_21976# a_30836_22020# VGND.t2775 VGND.t2774 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5345 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I VPWR.t3709 VPWR.t3708 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5346 VPWR.t18 _397_.A1.t12 _412_.A1 VPWR.t17 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5347 a_29164_25940# _336_.A1 _337_.ZN VGND.t4053 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5348 a_59620_27208# _244_.Z _247_.B VGND.t1776 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5349 a_53412_29480# _274_.A1 _274_.ZN VPWR.t2654 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X5350 a_9532_2727# a_9444_2824# VGND.t1159 VGND.t1158 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5351 a_57244_14136# a_57156_14180# VGND.t2039 VGND.t2038 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5352 VPWR.t5341 a_47164_14136# a_47076_14180# VPWR.t975 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5353 a_57244_11000# a_57156_11044# VGND.t5839 VGND.t5838 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5354 VPWR.t4051 a_47164_11000# a_47076_11044# VPWR.t3381 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5355 a_16240_26795# a_15828_27208.t6 VGND.t6114 VGND.t6113 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X5356 _231_.I vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN VPWR.t540 VPWR.t539 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5357 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I VGND.t4385 VGND.t4384 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5358 VGND.t6533 clk.t10 a_44296_24393.t10 VGND.t6532 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X5359 VPWR.t1438 a_60909_30600# a_61029_31220# VPWR.t1437 pfet_06v0 ad=0.1116p pd=0.98u as=61.19999f ps=0.7u w=0.36u l=0.5u
X5360 a_42168_25640.t2 _284_.A2.t6 _284_.ZN.t2 VGND.t28 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5361 VPWR.t6019 a_3708_6296# a_3620_6340# VPWR.t1188 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5362 VPWR.t585 a_42392_19243# _325_.A1.t0 VPWR.t584 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5363 VGND.t5663 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I VGND.t5662 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5364 VGND.t2239 _334_.A1 _293_.A2 VGND.t102 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X5365 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN VGND.t2085 VGND.t2084 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5366 VGND.t2117 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN VGND.t2116 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5367 VPWR.t4268 a_39324_17272# a_39236_17316# VPWR.t4267 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5368 VPWR.t1168 a_48529_22460# _279_.Z VPWR.t1167 pfet_06v0 ad=0.38705p pd=2.08u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5369 _330_.A1.t3 a_46198_27060# VGND.t1539 VGND.t1538 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5370 a_59036_2727# a_58948_2824# VGND.t1362 VGND.t751 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5371 VPWR.t5094 a_3708_3160# a_3620_3204# VPWR.t3110 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5372 a_54444_24679# a_54356_24776# VGND.t1363 VGND.t551 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5373 VPWR.t5318 a_23084_30951# a_22996_31048# VPWR.t5317 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5374 a_4156_26247# a_4068_26344# VGND.t1364 VGND.t555 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5375 VGND.t4730 _340_.A2 _340_.ZN VGND.t4729 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X5376 VPWR.t2683 a_9084_1159# a_8996_1256# VPWR.t2682 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5377 VPWR.t2353 _334_.A1 _335_.ZN.t2 VPWR.t2352 pfet_06v0 ad=0.4056p pd=1.805u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5378 a_4156_23111# a_4068_23208# VGND.t1366 VGND.t1365 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5379 VPWR.t736 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I VPWR.t735 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5380 a_66764_13703# a_66676_13800# VGND.t1368 VGND.t1367 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5381 _384_.A3.t0 _281_.A1 VPWR.t3296 VPWR.t3295 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5382 VPWR.t1748 a_53660_21543# a_53572_21640# VPWR.t1747 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5383 VPWR.t1058 a_66092_19975# a_66004_20072# VPWR.t1057 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5384 VGND.t6613 a_42392_22825.t33 _452_.CLK.t19 VGND.t6612 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5385 VPWR.t3889 vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN VPWR.t3888 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5386 VPWR.t567 a_29356_20408# a_29268_20452# VPWR.t566 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5387 a_55564_13703# a_55476_13800# VGND.t1370 VGND.t1369 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5388 a_25232_27165# a_24860_27209# VGND.t5185 VGND.t5184 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X5389 VGND.t1361 a_60909_30600# a_61029_30644# VGND.t45 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X5390 VPWR.t1064 a_63068_19975# a_62980_20072# VPWR.t1063 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5391 a_22636_29383# a_22548_29480# VGND.t5095 VGND.t2617 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5392 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I VPWR.t1742 VPWR.t1741 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5393 a_34716_20937# _319_.ZN a_34592_20569# VPWR.t2708 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X5394 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I VPWR.t5888 VPWR.t5887 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5395 a_48292_26369# _381_.A2.t5 VPWR.t6983 VPWR.t6982 pfet_06v0 ad=0.4599p pd=1.935u as=0.3918p ps=1.815u w=1.095u l=0.5u
X5396 VGND.t2156 a_51576_25896# _397_.A1.t1 VGND.t2155 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5397 a_17036_20408# a_16948_20452# VGND.t2026 VGND.t2025 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5398 a_26970_29480# _355_.C.t14 _373_.ZN VPWR.t6675 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5399 a_46100_26399# _402_.ZN a_45232_25987# VPWR.t3630 pfet_06v0 ad=54f pd=0.66u as=0.1872p ps=1.4u w=0.36u l=0.5u
X5400 VPWR.t392 a_62956_10567# a_62868_10664# VPWR.t391 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5401 a_57132_12135# a_57044_12232# VGND.t3392 VGND.t3391 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5402 VPWR.t5732 a_20060_21543# a_19972_21640# VPWR.t5731 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5403 a_54108_15271# a_54020_15368# VGND.t1372 VGND.t1371 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5404 a_36748_23544# a_36660_23588# VGND.t1374 VGND.t1373 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5405 VPWR.t888 a_28054_30196# _355_.C.t0 VPWR.t887 pfet_06v0 ad=0.4941p pd=2.03u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5406 VPWR.t682 a_50188_13703# a_50100_13800# VPWR.t681 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5407 VPWR.t878 a_54420_21976# a_54040_22366# VPWR.t877 pfet_06v0 ad=0.23p pd=1.54u as=0.352p ps=2.48u w=0.8u l=0.5u
X5408 _474_.CLK.t24 a_48272_25156.t38 VPWR.t6565 VPWR.t6564 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5409 _336_.Z a_28820_24072# VGND.t3699 VGND.t3698 nfet_06v0 ad=0.3586p pd=2.51u as=0.23405p ps=1.555u w=0.815u l=0.6u
X5410 VGND.t285 a_44296_24393.t34 clkbuf_1_0__f_clk.I.t22 VGND.t284 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5411 VPWR.t6200 a_25100_30951# a_25012_31048# VPWR.t6199 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5412 a_31168_24419# a_30796_24463# VPWR.t3131 VPWR.t3130 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X5413 a_58588_26247# a_58500_26344# VGND.t902 VGND.t901 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5414 a_64972_26680# a_64884_26724# VGND.t2306 VGND.t2305 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5415 VPWR.t4670 a_54432_31128# _304_.B VPWR.t4669 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5416 VPWR.t3997 a_21852_23111# a_21764_23208# VPWR.t3996 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5417 VGND.t3248 _327_.A2 _433_.ZN VGND.t3247 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5418 VPWR.t376 a_7740_29816# a_7652_29860# VPWR.t375 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5419 _304_.ZN.t0 _303_.ZN a_42252_20936# VGND.t2812 nfet_06v0 ad=0.30965p pd=1.685u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5420 VPWR.t925 a_44700_1159# a_44612_1256# VPWR.t924 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5421 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN VGND.t536 VGND.t535 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5422 a_29163_24394# _336_.Z _355_.ZN VGND.t4412 nfet_06v0 ad=85.2f pd=0.95u as=0.21175p ps=1.41u w=0.71u l=0.6u
X5423 a_3260_20408# a_3172_20452# VGND.t5443 VGND.t3668 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5424 _349_.A4 a_26720_30301# VGND.t4242 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5425 VGND.t2991 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN VGND.t2990 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5426 VPWR.t6135 a_44476_15704# a_44388_15748# VPWR.t1894 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5427 VPWR.t2952 _303_.ZN a_43380_20452# VPWR.t2951 pfet_06v0 ad=0.3918p pd=1.815u as=0.4599p ps=1.935u w=1.095u l=0.5u
X5428 VPWR.t6001 a_62396_14136# a_62308_14180# VPWR.t6000 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5429 a_4156_16839# a_4068_16936# VGND.t906 VGND.t905 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5430 vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN VGND.t5992 VGND.t5991 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5431 a_27116_21976# a_27028_22020# VGND.t5448 VGND.t5447 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5432 a_36188_26247# a_36100_26344# VGND.t908 VGND.t907 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5433 a_2364_4295# a_2276_4392# VGND.t372 VGND.t371 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5434 a_30812_16839# a_30724_16936# VGND.t910 VGND.t909 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5435 VPWR.t2490 a_17036_21976# a_16948_22020# VPWR.t2489 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5436 VPWR.t4577 a_43916_16839# a_43828_16936# VPWR.t4576 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5437 VPWR.t5484 a_56348_15271# a_56260_15368# VPWR.t5483 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5438 _250_.C _230_.I.t14 a_61940_29076# VGND.t6349 nfet_06v0 ad=0.4161p pd=1.905u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5439 a_24392_28248# _454_.Q a_24780_28776# VGND.t3934 nfet_06v0 ad=0.1606p pd=1.61u as=58.39999f ps=0.685u w=0.365u l=0.6u
X5440 VGND.t2313 a_48104_30219# _397_.A2.t2 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5441 VPWR.t1926 a_62396_11000# a_62308_11044# VPWR.t1925 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5442 VPWR.t4239 a_51196_14136# a_51108_14180# VPWR.t4238 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5443 VGND.t4336 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN VGND.t4335 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5444 VPWR.t4585 a_1020_7431# a_932_7528# VPWR.t482 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5445 uo_out[1].t7 _284_.ZN.t33 a_39300_29480# VPWR.t6522 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5446 VPWR.t3518 a_10204_1592# a_10116_1636# VPWR.t3517 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5447 VPWR.t1184 a_51196_11000# a_51108_11044# VPWR.t1183 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5448 VPWR.t4786 a_4940_10567# a_4852_10664# VPWR.t4785 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5449 a_31932_1159# a_31844_1256# VGND.t3791 VGND.t3790 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5450 VPWR.t3390 a_57580_17272# a_57492_17316# VPWR.t3389 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5451 VPWR.t3392 a_65756_17272# a_65668_17316# VPWR.t3391 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5452 VPWR.t2524 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I VPWR.t2523 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5453 a_34172_1592# a_34084_1636# VGND.t893 VGND.t892 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5454 VPWR.t6054 a_50636_12135# a_50548_12232# VPWR.t6053 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5455 VPWR.t4368 a_63404_13703# a_63316_13800# VPWR.t4367 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5456 VPWR.t4030 a_3260_21976# a_3172_22020# VPWR.t3819 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5457 VPWR.t4787 a_1916_10567# a_1828_10664# VPWR.t1800 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5458 a_58140_1592# a_58052_1636# VGND.t894 VGND.t848 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5459 VPWR.t6539 _362_.B.t15 _335_.ZN.t12 VPWR.t6538 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5460 VPWR.t4789 a_42908_2727# a_42820_2824# VPWR.t4788 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5461 VPWR.t4790 a_45820_18407# a_45732_18504# VPWR.t2515 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5462 _384_.A3.t8 _475_.Q VPWR.t5000 VPWR.t4999 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5463 VGND.t4649 _474_.Q a_52434_22504# VGND.t4648 nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X5464 uio_out[7].t5 a_18096_27165# VGND.t390 VGND.t389 nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X5465 VPWR.t5774 a_14796_27815# a_14708_27912# VPWR.t4177 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5466 a_12892_2727# a_12804_2824# VGND.t896 VGND.t895 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5467 a_56368_26344# vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I VPWR.t4436 VPWR.t4435 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5468 VGND.t113 _411_.A2.t11 a_51016_25940# VGND.t112 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5469 a_46800_20937# a_45920_20523# a_46476_20937# VGND.t1976 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X5470 VGND.t1304 a_66787_30600# _256_.A2.t1 VGND.t34 nfet_06v0 ad=0.28262p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5471 a_49672_19668# _474_.Q _417_.Z VGND.t4647 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5472 VPWR.t1357 a_19744_30301# a_19716_29977# VPWR.t1356 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X5473 VPWR.t4897 a_36636_2727# a_36548_2824# VPWR.t4896 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5474 VPWR.t2906 a_32156_17272# a_32068_17316# VPWR.t2905 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5475 VPWR.t6306 a_43296_28733# a_43288_28409# VPWR.t6305 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X5476 a_3260_14136# a_3172_14180# VGND.t3618 VGND.t854 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5477 VPWR.t1382 a_11091_30644# uio_oe[4].t0 VPWR.t1381 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5478 VPWR.t4745 a_11996_1592# a_11908_1636# VPWR.t4744 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5479 a_36636_21543# a_36548_21640# VGND.t2095 VGND.t2094 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5480 a_25436_24679# a_25348_24776# VGND.t1307 VGND.t1306 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5481 a_56720_26344# a_55956_25940# a_56516_26344# VPWR.t2499 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5482 a_3260_11000# a_3172_11044# VGND.t3221 VGND.t2707 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5483 VPWR.t4751 a_35964_1592# a_35876_1636# VPWR.t4750 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5484 VPWR.t3929 a_53212_14136# a_53124_14180# VPWR.t3928 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5485 VGND.t4029 a_41160_29083# uo_out[3].t5 VGND.t4028 nfet_06v0 ad=0.23432p pd=1.94u as=0.1183p ps=0.975u w=0.455u l=0.6u
X5486 a_40464_27165# a_40092_27209# VGND.t528 VGND.t527 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X5487 a_25436_21543# a_25348_21640# VGND.t1790 VGND.t1789 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5488 VPWR.t4593 a_19164_24679# a_19076_24776# VPWR.t4592 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5489 a_53660_27815# a_53572_27912# VGND.t4320 VGND.t4319 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5490 VPWR.t4475 a_59932_1592# a_59844_1636# VPWR.t2551 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5491 vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN VGND.t3595 VGND.t3594 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5492 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN VGND.t826 VGND.t825 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5493 VPWR.t3713 a_53212_11000# a_53124_11044# VPWR.t3712 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5494 VGND.t4840 a_43750_23544# a_43890_24164# VGND.t4839 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X5495 VPWR.t5764 a_32828_21543# a_32740_21640# VPWR.t5763 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5496 a_27004_23111# a_26916_23208# VGND.t1309 VGND.t1308 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5497 a_29575_28293# _369_.ZN _370_.ZN VPWR.t3101 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5498 VPWR.t3858 a_66652_4295# a_66564_4392# VPWR.t3436 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5499 a_32268_20408# a_32180_20452# VGND.t2848 VGND.t2847 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5500 a_49840_19001# a_48888_19243# VPWR.t2891 VPWR.t2890 pfet_06v0 ad=50.4f pd=0.64u as=0.23p ps=1.54u w=0.36u l=0.5u
X5501 _265_.ZN _324_.C.t29 VPWR.t6813 VPWR.t6812 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X5502 a_39324_15271# a_39236_15368# VGND.t1229 VGND.t1228 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5503 a_5388_10567# a_5300_10664# VGND.t1231 VGND.t1230 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5504 VGND.t4241 a_26720_30301# a_26672_30345# VGND.t137 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X5505 VPWR.t712 a_66652_1159# a_66564_1256# VPWR.t711 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5506 _424_.B2 _424_.A1 a_51912_20452# VPWR.t302 pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5507 a_61164_12135# a_61076_12232# VGND.t4089 VGND.t4088 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5508 VPWR.t953 a_17148_1159# a_17060_1256# VPWR.t952 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5509 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[1\].I VPWR.t1425 VPWR.t1424 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5510 a_40880_23588# _260_.A1 a_40656_23588# VPWR.t3913 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5511 VPWR.t5040 _274_.A3 a_53616_29480# VPWR.t5039 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X5512 a_36836_20072# _325_.A2.t9 a_36612_20072# VPWR.t6395 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5513 VPWR.t969 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I VPWR.t968 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5514 VPWR.t621 a_2364_24679# a_2276_24776# VPWR.t620 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5515 a_57020_2727# a_56932_2824# VGND.t1233 VGND.t1232 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5516 a_46268_18407# a_46180_18504# VGND.t1235 VGND.t1234 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5517 VGND.t5228 _245_.I1 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t5227 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5518 VGND.t3731 a_34448_25597# a_34400_25641# VGND.t3730 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X5519 a_57692_14136# a_57604_14180# VGND.t3863 VGND.t3862 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5520 VPWR.t4528 a_29244_23111# a_29156_23208# VPWR.t4527 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5521 a_36404_19001# a_35092_19368.t5 a_36060_19369# VPWR.t90 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X5522 VGND.t987 a_55312_22340# a_55208_22505# VGND.t986 nfet_06v0 ad=0.2637p pd=1.825u as=93.59999f ps=0.88u w=0.36u l=0.6u
X5523 VPWR.t3781 a_32268_21976# a_32180_22020# VPWR.t3780 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5524 a_21292_30951# a_21204_31048# VGND.t1236 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5525 a_60940_28248# a_60852_28292# VGND.t3169 VGND.t3168 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5526 vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN VPWR.t5612 VPWR.t5611 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5527 VGND.t6490 _287_.A1.t29 uo_out[4].t4 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X5528 a_61297_30300# _229_.I.t11 a_61689_29860# VPWR.t6876 pfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.5u
X5529 a_48321_23208# _399_.A1 _399_.ZN VPWR.t4236 pfet_06v0 ad=0.32805p pd=1.755u as=0.37665p ps=1.835u w=1.215u l=0.5u
X5530 a_57692_11000# a_57604_11044# VGND.t2886 VGND.t2885 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5531 a_60013_26344# _252_.B a_59397_26344# VPWR.t790 pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X5532 VPWR.t4200 a_21068_21976# a_20980_22020# VPWR.t4199 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5533 a_10092_30951# a_10004_31048# VGND.t1080 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5534 VPWR.t4770 a_59820_13703# a_59732_13800# VPWR.t3787 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5535 a_61612_13703# a_61524_13800# VGND.t1082 VGND.t1081 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5536 _304_.ZN.t8 _452_.Q.t16 a_42252_20936# VGND.t6641 nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5537 a_4940_19975# a_4852_20072# VGND.t1084 VGND.t1083 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5538 VPWR.t3845 a_24204_20408# a_24116_20452# VPWR.t3844 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5539 a_39548_2727# a_39460_2824# VGND.t1086 VGND.t1085 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5540 a_62796_25640# a_62560_25112# a_61836_25515# VGND.t2464 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5541 a_3708_25112# a_3620_25156# VGND.t1087 VGND.t63 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5542 a_1916_19975# a_1828_20072# VGND.t1089 VGND.t1088 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5543 VGND.t4531 _304_.B a_52081_21236# VGND.t4530 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5544 a_54892_24679# a_54804_24776# VGND.t1091 VGND.t1090 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5545 VPWR.t626 a_58588_2727# a_58500_2824# VPWR.t625 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5546 a_16700_1592# a_16612_1636# VGND.t1092 VGND.t67 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5547 VPWR.t3589 a_58028_12135# a_57940_12232# VPWR.t3588 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5548 _461_.D _362_.ZN VGND.t5564 VGND.t38 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X5549 a_3708_21976# a_3620_22020# VGND.t2936 VGND.t2935 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5550 VPWR.t4844 a_64300_23111# a_64212_23208# VPWR.t4409 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5551 VPWR.t6483 _459_.CLK.t36 a_28820_30344.t0 VPWR.t6482 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X5552 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I VPWR.t1588 VPWR.t1587 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5553 _412_.ZN _412_.A1 a_51332_24372# VGND.t1186 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5554 VPWR.t5296 a_5276_2727# a_5188_2824# VPWR.t5295 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5555 a_45372_15704# a_45284_15748# VGND.t1094 VGND.t1093 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5556 a_18760_29032# _379_.A2 a_19140_29612# VPWR.t2734 pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X5557 _432_.ZN _441_.A3 VGND.t1680 VGND.t1679 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5558 a_44752_18147# a_44459_18559# VPWR.t3207 VPWR.t3206 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X5559 VPWR.t4350 a_9308_1592# a_9220_1636# VPWR.t4349 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5560 a_35740_1159# a_35652_1256# VGND.t4631 VGND.t4630 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5561 VPWR.t1086 a_2364_15271# a_2276_15368# VPWR.t1085 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5562 VPWR.t5150 a_50524_15704# a_50436_15748# VPWR.t5149 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5563 a_26112_27209# a_23892_27208.t7 a_25867_26841# VGND.t6071 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X5564 a_61276_2727# a_61188_2824# VGND.t957 VGND.t956 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5565 VPWR.t6841 clk.t11 a_44296_24393.t11 VPWR.t6840 pfet_06v0 ad=0.3608p pd=2.52u as=0.2542p ps=1.44u w=0.82u l=0.5u
X5566 VPWR.t4709 a_34396_24679# a_34308_24776# VPWR.t4708 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5567 a_45396_22020# _304_.B _324_.B.t4 VPWR.t4686 pfet_06v0 ad=0.4599p pd=1.935u as=0.2847p ps=1.615u w=1.095u l=0.5u
X5568 a_65756_9432# a_65668_9476# VGND.t959 VGND.t958 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5569 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN VGND.t5661 VGND.t5660 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5570 a_48272_25156.t9 clkbuf_1_0__f_clk.I.t53 VGND.t265 VGND.t264 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X5571 VGND.t6643 _452_.Q.t17 _439_.ZN VGND.t6642 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X5572 VPWR.t4715 a_23196_24679# a_23108_24776# VPWR.t4714 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5573 a_65756_6296# a_65668_6340# VGND.t4035 VGND.t4034 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5574 a_17484_20408# a_17396_20452# VGND.t3541 VGND.t3540 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5575 a_57580_12135# a_57492_12232# VGND.t3551 VGND.t3550 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5576 a_54556_15271# a_54468_15368# VGND.t961 VGND.t960 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5577 a_4156_3160# a_4068_3204# VGND.t2541 VGND.t2540 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5578 a_52036_22504# _281_.A1 _384_.A3.t2 VGND.t3144 nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5579 a_31036_23111# a_30948_23208# VGND.t963 VGND.t962 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5580 a_59484_9432# a_59396_9476# VGND.t5065 VGND.t5064 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5581 a_43288_28409# a_41440_28363# a_43003_28409# VPWR.t1519 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X5582 VPWR.t3806 a_5388_27815# a_5300_27912# VPWR.t3805 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5583 VPWR.t4511 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN VPWR.t4510 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5584 VPWR.t309 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN VPWR.t308 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5585 _350_.A1.t1 a_29856_29123# VGND.t3057 VGND.t3056 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5586 a_52081_21236# _476_.Q a_51877_21236# VGND.t4159 nfet_06v0 ad=0.1312p pd=1.14u as=0.1722p ps=1.24u w=0.82u l=0.6u
X5587 VGND.t6143 _337_.A3.t12 _351_.A2 VGND.t6142 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X5588 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I VPWR.t6176 VPWR.t2525 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5589 a_43892_20072# _325_.A1.t17 _325_.B VPWR.t4699 pfet_06v0 ad=0.3172p pd=1.74u as=0.4016p ps=1.94u w=1.22u l=0.5u
X5590 VPWR.t3810 a_57244_27815# a_57156_27912# VPWR.t3809 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5591 a_3708_15704# a_3620_15748# VGND.t1878 VGND.t1877 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5592 a_14796_23544# a_14708_23588# VGND.t1880 VGND.t1879 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5593 a_32156_15271# a_32068_15368# VGND.t1882 VGND.t1881 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5594 a_33948_19975# a_33860_20072# VGND.t1884 VGND.t1883 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5595 VPWR.t4685 _304_.B _304_.ZN.t2 VPWR.t4684 pfet_06v0 ad=0.5292p pd=3.14u as=0.2808p ps=1.6u w=1.08u l=0.5u
X5596 a_27564_21976# a_27476_22020# VGND.t3095 VGND.t3094 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5597 VPWR.t1697 a_17484_21976# a_17396_22020# VPWR.t1696 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5598 VPWR.t4613 a_18940_1159# a_18852_1256# VPWR.t4612 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5599 VPWR.t2381 a_25792_30301# a_25764_29977# VPWR.t2380 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X5600 VPWR.t4666 a_56796_15271# a_56708_15368# VPWR.t4665 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5601 VPWR.t4668 a_33276_23111# a_33188_23208# VPWR.t4667 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5602 VGND.t4529 _304_.B a_49764_26724# VGND.t4528 nfet_06v0 ad=0.224p pd=1.52u as=0.14p ps=1.1u w=0.4u l=0.6u
X5603 VPWR.t6502 _397_.A2.t15 _411_.A2.t0 VPWR.t6501 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5604 VPWR.t4811 a_34620_2727# a_34532_2824# VPWR.t4810 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5605 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN VPWR.t3149 VPWR.t3148 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5606 a_45260_16839# a_45172_16936# VGND.t1886 VGND.t1885 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5607 a_14684_1592# a_14596_1636# VGND.t1888 VGND.t1887 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5608 a_35156_29860# _287_.A1.t30 uo_out[4].t6 VPWR.t6788 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X5609 VPWR.t5920 _293_.A2 a_39748_29480# VPWR.t5919 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5610 a_1916_8999# a_1828_9096# VGND.t1889 VGND.t652 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5611 VPWR.t4754 a_64860_8999# a_64772_9096# VPWR.t3967 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5612 a_39300_31048# _296_.ZN VPWR.t3661 VPWR.t3660 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X5613 a_38652_1592# a_38564_1636# VGND.t1891 VGND.t1890 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5614 a_19500_20408# a_19412_20452# VGND.t2346 VGND.t2345 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5615 VPWR.t4848 a_63852_13703# a_63764_13800# VPWR.t4847 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5616 uo_out[1].t9 _293_.A2 VGND.t5701 VGND.t5700 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X5617 a_38523_27967# a_36960_27912# a_37888_27555# VGND.t5297 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X5618 a_1916_5863# a_1828_5960# VGND.t2143 VGND.t2142 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5619 VPWR.t6163 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I VPWR.t6162 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5620 VPWR.t3764 a_55228_28248# a_55140_28292# VPWR.t1149 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5621 VPWR.t5812 a_60604_9432# a_60516_9476# VPWR.t5811 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5622 VPWR.t5478 a_21404_1159# a_21316_1256# VPWR.t5477 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5623 VGND.t3611 _267_.A2 a_52891_28776# VGND.t3610 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5624 a_66540_18407# a_66452_18504# VGND.t1893 VGND.t1892 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5625 a_3260_10567# a_3172_10664# VGND.t1894 VGND.t646 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5626 a_28891_25273# a_27328_25227# a_28256_25597# VGND.t6028 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X5627 vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN VGND.t2018 VGND.t2017 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5628 a_35504_18955# a_35092_19368.t6 VPWR.t92 VPWR.t91 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X5629 VPWR.t6992 _352_.A2.t26 a_25524_26344# VPWR.t6991 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5630 a_39475_21236# _451_.Q.t9 VGND.t6154 VGND.t6153 nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5631 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I VGND.t2022 VGND.t2021 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5632 VPWR.t5787 a_54332_9432# a_54244_9476# VPWR.t5786 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5633 a_63516_18407# a_63428_18504# VGND.t1895 VGND.t701 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5634 VPWR.t3421 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN VPWR.t3068 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5635 VPWR.t3230 a_40264_30320# _294_.A2.t0 VPWR.t3229 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5636 a_41116_1592# a_41028_1636# VGND.t1897 VGND.t1896 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5637 VPWR.t3842 a_15132_1159# a_15044_1256# VPWR.t2606 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5638 VPWR.t4942 a_46940_15704# a_46852_15748# VPWR.t4305 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5639 VPWR.t4420 a_5388_18407# a_5300_18504# VPWR.t4419 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5640 a_46804_28292# _389_.ZN a_46580_28292# VPWR.t5305 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5641 a_25888_25641# a_23668_25640.t6 a_25643_25273# VGND.t6710 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X5642 a_31803_24831# a_29828_24455.t6 a_31168_24419# VPWR.t6387 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X5643 a_25884_24679# a_25796_24776# VGND.t1899 VGND.t1898 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5644 VPWR.t628 a_39100_1159# a_39012_1256# VPWR.t627 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5645 VPWR.t2931 a_54192_22851# a_54088_22895# VPWR.t2930 pfet_06v0 ad=0.1044p pd=0.94u as=0.1791p ps=1.355u w=0.36u l=0.5u
X5646 a_62172_17272# a_62084_17316# VGND.t965 VGND.t964 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5647 VPWR.t5788 a_1020_9432# a_932_9476# VPWR.t4883 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5648 a_63740_14136# a_63652_14180# VGND.t2391 VGND.t2390 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5649 vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN VPWR.t4650 VPWR.t4649 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5650 a_40644_17272# a_41048_17341# a_40992_17433# VPWR.t5011 pfet_06v0 ad=0.1665p pd=1.285u as=50.4f ps=0.64u w=0.36u l=0.5u
X5651 a_60380_1592# a_60292_1636# VGND.t806 VGND.t805 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5652 VPWR.t1845 a_53660_14136# a_53572_14180# VPWR.t1844 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5653 VPWR.t5069 a_35740_15704# a_35652_15748# VPWR.t5068 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5654 _241_.Z a_56964_26724# VGND.t5532 VGND.t5531 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5655 a_36828_28776# _362_.B.t16 a_34084_28776# VGND.t6256 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5656 a_25884_21543# a_25796_21640# VGND.t2113 VGND.t2112 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5657 VPWR.t2460 a_48060_9432# a_47972_9476# VPWR.t2459 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5658 VGND.t4862 a_37888_27555# a_37840_27599# VGND.t4861 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X5659 a_63740_11000# a_63652_11044# VGND.t496 VGND.t495 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5660 a_52540_14136# a_52452_14180# VGND.t498 VGND.t497 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5661 a_4156_26680# a_4068_26724# VGND.t3109 VGND.t1574 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5662 VPWR.t534 a_53660_11000# a_53572_11044# VPWR.t533 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5663 a_27452_23111# a_27364_23208# VGND.t808 VGND.t807 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5664 VPWR.t1238 a_16588_24679# a_16500_24776# VPWR.t1237 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5665 a_52540_11000# a_52452_11044# VGND.t2350 VGND.t2349 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5666 a_43804_2727# a_43716_2824# VGND.t810 VGND.t809 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5667 VPWR.t4925 a_36412_15271# a_36324_15368# VPWR.t4924 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5668 VPWR.t4660 a_2812_13703# a_2724_13800# VPWR.t3908 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5669 a_39772_15271# a_39684_15368# VGND.t812 VGND.t811 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5670 a_29351_28293# _359_.B.t11 VPWR.t6775 VPWR.t6774 pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X5671 VPWR.t775 _282_.ZN _284_.B VPWR.t774 pfet_06v0 ad=0.3918p pd=1.815u as=0.2808p ps=1.6u w=1.08u l=0.5u
X5672 VPWR.t2668 a_62844_2727# a_62756_2824# VPWR.t2667 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5673 VPWR.t5309 a_42908_1592# a_42820_1636# VPWR.t5308 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5674 a_53996_25112# a_53908_25156# VGND.t5505 VGND.t5504 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5675 a_65868_10567# a_65780_10664# VGND.t814 VGND.t813 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5676 a_37532_2727# a_37444_2824# VGND.t816 VGND.t815 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5677 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I VGND.t2783 VGND.t2782 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5678 a_65308_18840# a_65220_18884# VGND.t2904 VGND.t2903 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5679 _495_.I a_41056_30669# VPWR.t6228 VPWR.t6227 pfet_06v0 ad=0.31207p pd=1.665u as=0.34437p ps=1.895u w=1.095u l=0.5u
X5680 a_66876_1592# a_66788_1636# VGND.t818 VGND.t817 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5681 VPWR.t1937 a_14796_26680# a_14708_26724# VPWR.t1936 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5682 VGND.t6444 _268_.A1.t8 _275_.A2 VGND.t6443 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X5683 a_54668_10567# a_54580_10664# VGND.t792 VGND.t791 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5684 VPWR.t4304 a_67548_8999# a_67460_9096# VPWR.t4010 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5685 a_62620_15704# a_62532_15748# VGND.t794 VGND.t793 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5686 VPWR.t1240 a_56572_2727# a_56484_2824# VPWR.t1239 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5687 VPWR.t4442 a_29692_23111# a_29604_23208# VPWR.t4441 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5688 VGND.t1458 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN _249_.A2 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5689 a_28596_27916.t5 _371_.A2 VPWR.t3578 VPWR.t3577 pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X5690 a_37348_27599# a_36548_27591.t4 VGND.t6325 VGND.t6324 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5691 VPWR.t6816 a_3260_5863# a_3172_5960# VPWR.t2754 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5692 a_51420_15704# a_51332_15748# VGND.t796 VGND.t795 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5693 a_59605_25962# _231_.ZN VGND.t4199 VGND.t4198 nfet_06v0 ad=85.2f pd=0.95u as=0.3124p ps=2.3u w=0.71u l=0.6u
X5694 VPWR.t6523 _284_.ZN.t34 a_38472_30169# VPWR.t6517 pfet_06v0 ad=0.3608p pd=2.52u as=0.2542p ps=1.44u w=0.82u l=0.5u
X5695 _371_.ZN _371_.A1.t17 a_28112_27912# VPWR.t6512 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5696 VPWR.t1244 a_3260_2727# a_3172_2824# VPWR.t1243 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5697 a_35040_20937# a_34160_20523# a_34716_20937# VGND.t2764 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X5698 a_27900_21543# a_27812_21640# VGND.t2062 VGND.t2061 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5699 a_37179_24831# a_35204_24455.t6 a_36544_24419# VPWR.t6398 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X5700 a_27716_25641# a_26916_25640.t6 VGND.t6474 VGND.t6473 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5701 VPWR.t2326 a_17036_27815# a_16948_27912# VPWR.t2325 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5702 VPWR.t5399 a_43356_1159# a_43268_1256# VPWR.t2072 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5703 a_37860_27967# a_36548_27591.t5 a_37516_27599# VPWR.t6615 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X5704 a_7292_1592# a_7204_1636# VGND.t798 VGND.t797 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5705 VGND.t722 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I VGND.t721 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5706 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN VGND.t6015 VGND.t6014 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5707 VPWR.t1893 a_24652_20408# a_24564_20452# VPWR.t1892 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5708 a_35628_16839# a_35540_16936# VGND.t800 VGND.t799 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5709 a_68108_20408# a_68020_20452# VGND.t994 VGND.t993 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5710 VPWR.t2512 a_58028_20408# a_57940_20452# VPWR.t2511 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5711 a_63740_9432# a_63652_9476# VGND.t4851 VGND.t4850 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5712 VPWR.t2601 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN VPWR.t2600 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5713 a_40644_17272# a_41088_17757.t7 a_41040_17801# VGND.t162 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X5714 a_36188_26680# a_36100_26724# VGND.t2197 VGND.t2196 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5715 VPWR.t5194 a_51084_28248# a_50996_28292# VPWR.t5193 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5716 VPWR.t853 a_37084_1159# a_36996_1256# VPWR.t852 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5717 VPWR.t1422 a_58476_12135# a_58388_12232# VPWR.t1421 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5718 a_63068_1592# a_62980_1636# VGND.t839 VGND.t838 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5719 a_51968_20127# a_51240_19624# VPWR.t4566 VPWR.t4565 pfet_06v0 ad=50.4f pd=0.64u as=0.23p ps=1.54u w=0.36u l=0.5u
X5720 a_24860_27209# _351_.ZN a_24692_27209# VGND.t2191 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X5721 VGND.t6023 _260_.A2 a_44491_20936# VGND.t6022 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X5722 a_19320_28409# a_17472_28363# a_19035_28409# VPWR.t2637 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X5723 VPWR.t2886 a_3260_27815# a_3172_27912# VPWR.t2885 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5724 VGND.t1378 a_40644_17272# a_40040_17675# VGND.t1377 nfet_06v0 ad=0.142p pd=1.14u as=0.176p ps=1.68u w=0.4u l=0.6u
X5725 a_36560_22512# _311_.A2.t9 VGND.t6109 VGND.t6108 nfet_06v0 ad=79.8f pd=0.8u as=0.2424p ps=1.635u w=0.38u l=0.6u
X5726 a_9980_2727# a_9892_2824# VGND.t841 VGND.t840 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5727 a_39780_22805# _441_.A2 _441_.ZN VGND.t4146 nfet_06v0 ad=0.2119p pd=1.335u as=0.4137p ps=1.9u w=0.815u l=0.6u
X5728 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I VPWR.t3119 VPWR.t3118 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5729 _432_.ZN _260_.A1 VGND.t3769 VGND.t3768 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X5730 VPWR.t4910 a_2364_23544# a_2276_23588# VPWR.t3965 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5731 a_56964_26724# _251_.A1.t29 a_56816_26724# VPWR.t7020 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X5732 _284_.ZN.t8 _304_.B a_42168_25640.t4 VGND.t4527 nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5733 a_5276_30951# a_5188_31048# VGND.t842 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5734 _268_.A2.t0 a_50436_30689# VPWR.t2114 VPWR.t2113 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X5735 a_41788_2727# a_41700_2824# VGND.t844 VGND.t843 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5736 VPWR.t4913 a_52092_1592# a_52004_1636# VPWR.t4912 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5737 VGND.t6111 _311_.A2.t10 a_35188_22895# VGND.t6110 nfet_06v0 ad=0.23405p pd=1.555u as=58.39999f ps=0.685u w=0.365u l=0.6u
X5738 VPWR.t4917 a_50972_15704# a_50884_15748# VPWR.t4916 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5739 a_66787_30600# a_67117_30600# a_67237_30644# VGND.t45 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X5740 a_65756_2727# a_65668_2824# VGND.t846 VGND.t845 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5741 VPWR.t1648 a_23532_21976# a_23444_22020# VPWR.t1647 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5742 a_52415_31220# a_51791_30644# a_52247_31220# VPWR.t5454 pfet_06v0 ad=0.3852p pd=2.86u as=61.19999f ps=0.7u w=0.36u l=0.5u
X5743 a_44364_17272# a_44276_17316# VGND.t679 VGND.t678 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5744 a_28596_26725# _336_.A2.t9 _355_.B VPWR.t172 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X5745 VGND.t6519 _325_.A1.t18 _439_.ZN VGND.t3247 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X5746 a_32848_29123# a_32476_29167# VGND.t4849 VGND.t4848 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X5747 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].I VPWR.t5201 VPWR.t1430 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5748 VPWR.t4457 a_51644_15271# a_51556_15368# VPWR.t4456 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5749 _452_.CLK.t20 a_42392_22825.t34 VPWR.t6932 VPWR.t6931 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5750 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I _258_.ZN VPWR.t2151 VPWR.t2150 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5751 a_59484_2727# a_59396_2824# VGND.t5634 VGND.t1024 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5752 a_47164_12568# a_47076_12612# VGND.t1733 VGND.t1732 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5753 a_31484_23111# a_31396_23208# VGND.t5636 VGND.t5635 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5754 VPWR.t3737 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN VPWR.t3736 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5755 uio_out[5].t7 a_20672_30301# VGND.t4868 VGND.t71 nfet_06v0 ad=0.2119p pd=1.335u as=0.2608p ps=1.455u w=0.815u l=0.6u
X5756 _452_.CLK.t21 a_42392_22825.t35 VGND.t6615 VGND.t6614 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5757 _399_.A1 _395_.A1 a_50196_22805# VGND.t887 nfet_06v0 ad=0.4137p pd=1.9u as=0.2119p ps=1.335u w=0.815u l=0.6u
X5758 _288_.ZN.t1 _460_.Q VGND.t3326 VGND.t108 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X5759 a_6172_2727# a_6084_2824# VGND.t5638 VGND.t5637 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5760 _417_.Z _474_.Q a_49448_20072# VPWR.t4795 pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5761 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I VPWR.t505 VPWR.t504 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5762 VPWR.t457 a_58588_1592# a_58500_1636# VPWR.t456 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5763 a_3708_7864# a_3620_7908# VGND.t5640 VGND.t5639 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5764 a_45080_29535# a_43232_29480# a_44795_29535# VPWR.t804 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X5765 VPWR.t4829 a_56348_30951# a_56260_31048# VPWR.t4828 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5766 a_35008_22461# a_34715_22137# VGND.t2137 VGND.t2136 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X5767 a_35660_27508# _363_.Z.t6 _365_.ZN VGND.t37 nfet_06v0 ad=0.3608p pd=2.52u as=0.4161p ps=1.905u w=0.82u l=0.6u
X5768 a_3708_4728# a_3620_4772# VGND.t5946 VGND.t1130 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5769 a_50972_1159# a_50884_1256# VGND.t5642 VGND.t5641 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5770 VPWR.t1814 a_3260_18407# a_3172_18504# VPWR.t1813 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5771 VGND.t1907 a_37384_19624# _325_.A2.t1 VGND.t1906 nfet_06v0 ad=0.23405p pd=1.555u as=0.3586p ps=2.51u w=0.815u l=0.6u
X5772 a_36656_29123# a_36284_29167# VPWR.t4938 VPWR.t4937 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X5773 VGND.t2170 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN VGND.t2169 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5774 VPWR.t4284 a_45148_30951# a_45060_31048# VPWR.t4283 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5775 a_34960_22505# a_32740_22504.t6 a_34715_22137# VGND.t96 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X5776 clkbuf_1_0__f_clk.I.t21 a_44296_24393.t35 VGND.t287 VGND.t286 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5777 a_1020_4295# a_932_4392# VGND.t1675 VGND.t320 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5778 a_45408_30345# a_44632_30206# VGND.t819 VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=0.142p ps=1.14u w=0.36u l=0.6u
X5779 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv1.inv_array_notouch_\[1\].I VPWR.t2773 VPWR.t2772 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5780 VPWR.t1816 a_66988_16839# a_66900_16936# VPWR.t1815 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5781 a_31932_21543# a_31844_21640# VGND.t6035 VGND.t6034 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5782 VPWR.t1080 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I VPWR.t1079 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5783 a_33188_25940# _460_.Q _360_.ZN VGND.t3325 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5784 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I VGND.t1859 VGND.t1858 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5785 VPWR.t2522 a_55676_28248# a_55588_28292# VPWR.t2521 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5786 _402_.ZN _402_.A1.t19 a_46352_22021# VPWR.t6731 pfet_06v0 ad=0.3159p pd=1.735u as=0.44955p ps=1.955u w=1.215u l=0.5u
X5787 a_54108_21543# a_54020_21640# VGND.t1759 VGND.t1758 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5788 a_24636_25641# _457_.D a_24468_25641# VGND.t2817 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X5789 VPWR.t6070 a_1468_21543# a_1380_21640# VPWR.t4760 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5790 VGND.t6617 a_42392_22825.t36 _452_.CLK.t22 VGND.t6616 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5791 VPWR.t6072 a_9084_29383# a_8996_29480# VPWR.t6071 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5792 VPWR.t6485 _459_.CLK.t37 a_23892_27208.t0 VPWR.t6484 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X5793 a_42796_23981# a_43126_24119# a_43246_24163# VGND.t3216 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X5794 a_67100_8999# a_67012_9096# VGND.t4943 VGND.t4879 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5795 a_22300_23111# a_22212_23208# VGND.t4945 VGND.t4944 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5796 a_3260_29816# a_3172_29860# VGND.t4946 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5797 VPWR.t5520 a_58687_31220# a_59143_31198# VPWR.t5519 pfet_06v0 ad=0.379p pd=2.37u as=61.19999f ps=0.7u w=0.36u l=0.5u
X5798 a_21628_1592# a_21540_1636# VGND.t4948 VGND.t4947 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5799 a_45820_12135# a_45732_12232# VGND.t5535 VGND.t3037 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5800 a_34620_15271# a_34532_15368# VGND.t4950 VGND.t4949 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5801 a_63964_18407# a_63876_18504# VGND.t4951 VGND.t553 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5802 a_67100_5863# a_67012_5960# VGND.t3386 VGND.t3385 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5803 _231_.ZN _231_.I VPWR.t6167 VPWR.t6166 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5804 VPWR.t6662 _452_.CLK.t51 a_42484_18183.t0 VPWR.t6661 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X5805 VPWR.t1822 a_11324_2727# a_11236_2824# VPWR.t1821 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5806 VPWR.t2092 a_35740_26247# a_35652_26344# VPWR.t2091 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5807 VPWR.t3629 a_20844_26680# a_20756_26724# VPWR.t3628 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5808 a_60716_10567# a_60628_10664# VGND.t4953 VGND.t4952 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5809 VPWR.t4323 _476_.Q _424_.A1 VPWR.t4322 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5810 VPWR.t6233 a_13340_29383# a_13252_29480# VPWR.t5572 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5811 a_36516_24831# a_35204_24455.t7 a_36172_24463# VPWR.t6399 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X5812 VPWR.t4292 a_10652_1592# a_10564_1636# VPWR.t4291 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5813 VPWR.t1136 a_4940_19975# a_4852_20072# VPWR.t1135 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5814 vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN VGND.t2746 VGND.t1849 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5815 VGND.t4886 _274_.A3 a_52756_29076# VGND.t4885 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5816 VPWR.t4392 a_24540_23111# a_24452_23208# VPWR.t4391 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5817 VPWR.t4295 a_34620_1592# a_34532_1636# VPWR.t2314 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5818 a_45904_30180# a_45456_30301.t3 a_46316_29977# VPWR.t7058 pfet_06v0 ad=0.1872p pd=1.4u as=43.2f ps=0.6u w=0.36u l=0.5u
X5819 a_17036_23544# a_16948_23588# VGND.t403 VGND.t402 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5820 a_50308_26476# _411_.A2.t12 a_50120_26476# VPWR.t118 pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X5821 VPWR.t597 a_29020_2727# a_28932_2824# VPWR.t596 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5822 VPWR.t4394 a_36860_15271# a_36772_15368# VPWR.t4393 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5823 VPWR.t1142 a_1916_19975# a_1828_20072# VPWR.t1141 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5824 _324_.B.t16 _304_.ZN.t16 VPWR.t234 VPWR.t233 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5825 a_62396_12568# a_62308_12612# VGND.t1535 VGND.t1534 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5826 uio_out[0].t0 a_28124_30600# VGND.t5211 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5827 VPWR.t5679 a_65084_14136# a_64996_14180# VPWR.t5678 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5828 a_33500_16839# a_33412_16936# VGND.t405 VGND.t404 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5829 VPWR.t420 a_41340_1159# a_41252_1256# VPWR.t419 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5830 VPWR.t603 a_46604_16839# a_46516_16936# VPWR.t602 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5831 VPWR.t290 a_44296_24393.t36 clkbuf_1_0__f_clk.I.t4 VPWR.t289 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5832 a_51196_12568# a_51108_12612# VGND.t3526 VGND.t3525 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5833 VPWR.t2061 a_65084_11000# a_64996_11044# VPWR.t2060 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5834 a_57580_18840# a_57492_18884# VGND.t5819 VGND.t5818 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5835 _424_.B2 a_51240_20452# VGND.t461 VGND.t460 nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X5836 vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I VGND.t2692 VGND.t2691 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5837 a_65756_18840# a_65668_18884# VGND.t5823 VGND.t5822 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5838 VGND.t926 a_26160_27165# a_26112_27209# VGND.t925 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X5839 a_34155_25273# a_32180_25640.t6 a_33520_25597# VPWR.t40 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X5840 a_3260_23544# a_3172_23588# VGND.t409 VGND.t408 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5841 VPWR.t5278 a_1468_12135# a_1380_12232# VPWR.t1857 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5842 VPWR.t818 a_41392_27165# a_41384_26841# VPWR.t817 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X5843 VGND.t5720 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN VGND.t5719 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X5844 a_52400_25987.t1 _474_.CLK.t50 VGND.t6461 VGND.t6460 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X5845 VGND.t4454 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].I VGND.t71 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5846 VPWR.t5356 a_39884_27815# a_39796_27912# VPWR.t5355 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5847 VPWR.t5865 a_3708_7864# a_3620_7908# VPWR.t4244 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5848 VPWR.t1655 a_53324_12135# a_53236_12232# VPWR.t1654 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5849 a_49888_19369# a_48888_19243# VGND.t2762 VGND.t2761 nfet_06v0 ad=43.2f pd=0.6u as=0.142p ps=1.14u w=0.36u l=0.6u
X5850 _304_.A1.t0 a_35232_24029# VPWR.t5673 VPWR.t5672 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5851 VGND.t6372 _452_.CLK.t52 a_35092_19368.t1 VGND.t6371 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X5852 _305_.A2 a_41488_24072# VGND.t5428 VGND.t5427 nfet_06v0 ad=0.3586p pd=2.51u as=0.226p ps=1.515u w=0.815u l=0.6u
X5853 a_50464_24908# _281_.ZN.t8 VPWR.t124 VPWR.t123 pfet_06v0 ad=0.224p pd=1.36u as=0.389p ps=2.02u w=0.56u l=0.5u
X5854 a_20508_2727# a_20420_2824# VGND.t2831 VGND.t2830 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5855 VPWR.t2973 a_23868_1159# a_23780_1256# VPWR.t2972 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5856 a_43824_18147# a_43452_18191# VGND.t48 VGND.t47 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X5857 a_32156_18840# a_32068_18884# VGND.t5181 VGND.t5180 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5858 VPWR.t4581 a_19164_30951# a_19076_31048# VPWR.t4580 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5859 VPWR.t5545 a_17484_27815# a_17396_27912# VPWR.t5544 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5860 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN VGND.t6013 VGND.t6012 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5861 VPWR.t3306 _398_.C a_49316_23588# VPWR.t3305 pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X5862 a_48560_26369# _397_.A2.t16 a_48292_26369# VPWR.t6503 pfet_06v0 ad=0.33945p pd=1.715u as=0.4599p ps=1.935u w=1.095u l=0.5u
X5863 a_63740_2727# a_63652_2824# VGND.t2834 VGND.t1204 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5864 VPWR.t4631 a_16588_23544# a_16500_23588# VPWR.t1643 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5865 VPWR.t3522 a_56796_9432# a_56708_9476# VPWR.t3521 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5866 VPWR.t1965 a_58476_20408# a_58388_20452# VPWR.t1964 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5867 a_14236_2727# a_14148_2824# VGND.t2835 VGND.t1206 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5868 VPWR.t2978 a_17596_1159# a_17508_1256# VPWR.t2624 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5869 VPWR.t3078 a_2812_12568# a_2724_12612# VPWR.t3047 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5870 _438_.A2 a_37472_24419# VPWR.t2022 VPWR.t2021 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5871 a_26152_26841# a_24304_26795# a_25867_26841# VPWR.t1155 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X5872 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN VPWR.t1709 VPWR.t1708 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5873 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN VGND.t2728 VGND.t2727 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5874 uo_out[4].t9 _294_.ZN.t7 VGND.t149 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X5875 VPWR.t743 a_4156_7431# a_4068_7528# VPWR.t742 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5876 a_53212_12568# a_53124_12612# VGND.t1387 VGND.t1386 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5877 VPWR.t3399 _327_.A2 _303_.ZN VPWR.t3398 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X5878 VPWR.t749 a_33276_2727# a_33188_2824# VPWR.t748 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5879 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t734 VPWR.t733 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5880 a_42392_22825.t2 clkbuf_1_0__f_clk.I.t54 VPWR.t266 VPWR.t265 pfet_06v0 ad=0.2542p pd=1.44u as=0.428p ps=2.02u w=0.82u l=0.5u
X5881 a_54780_1159# a_54692_1256# VGND.t2804 VGND.t2803 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5882 _330_.A2 _327_.Z a_38644_19368# VGND.t5365 nfet_06v0 ad=0.4161p pd=1.905u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5883 VPWR.t1977 a_33948_19975# a_33860_20072# VPWR.t1976 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5884 _336_.A2.t0 a_25936_25597# VPWR.t5856 VPWR.t5855 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5885 a_1468_27815# a_1380_27912# VGND.t5799 VGND.t5798 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5886 VPWR.t5048 a_42778_21812# a_43214_21812# VPWR.t5047 pfet_06v0 ad=0.1656p pd=1.28u as=61.19999f ps=0.7u w=0.36u l=0.5u
X5887 VPWR.t4775 a_37308_1592# a_37220_1636# VPWR.t4774 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5888 vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN VGND.t1058 VGND.t1057 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5889 VPWR.t4893 a_2364_30951# a_2276_31048# VPWR.t4892 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5890 a_17472_28363# a_17060_28776.t6 VGND.t6595 VGND.t6594 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X5891 VPWR.t4396 a_49292_13703# a_49204_13800# VPWR.t4395 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5892 a_51084_13703# a_50996_13800# VGND.t3395 VGND.t3394 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5893 VGND.t1286 a_19744_30301# a_19696_30345# VGND.t137 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X5894 VPWR.t5898 a_3260_4728# a_3172_4772# VPWR.t4167 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5895 VPWR.t2983 a_16140_21543# a_16052_21640# VPWR.t2982 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5896 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I VGND.t4685 VGND.t4684 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5897 VPWR.t4903 a_17932_26247# a_17844_26344# VPWR.t4902 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5898 _324_.B.t12 _302_.Z VPWR.t4987 VPWR.t4986 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X5899 VPWR.t394 a_46268_13703# a_46180_13800# VPWR.t393 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5900 a_59260_21976# a_59172_22020# VGND.t4932 VGND.t823 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5901 VPWR.t2724 a_23980_21976# a_23892_22020# VPWR.t2723 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5902 a_50176_26724# _402_.A1.t20 a_49952_26724# VPWR.t6732 pfet_06v0 ad=0.224p pd=1.36u as=0.1736p ps=1.18u w=0.56u l=0.5u
X5903 _371_.A2 _337_.A3.t13 VPWR.t6409 VPWR.t6408 pfet_06v0 ad=0.2197p pd=1.365u as=0.4056p ps=1.805u w=0.845u l=0.5u
X5904 VPWR.t4885 a_3260_1592# a_3172_1636# VPWR.t2279 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5905 VPWR.t5884 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I VPWR.t5883 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5906 _427_.A2 _384_.A3.t17 a_51540_23588# VPWR.t186 pfet_06v0 ad=0.4016p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5907 a_30812_1159# a_30724_1256# VGND.t3766 VGND.t3765 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5908 a_54444_19975# a_54356_20072# VGND.t3397 VGND.t3396 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5909 a_68108_10567# a_68020_10664# VGND.t3399 VGND.t3398 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5910 a_22300_1159# a_22212_1256# VGND.t3401 VGND.t3400 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5911 VPWR.t4889 a_29804_23544# a_29716_23588# VPWR.t4888 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5912 VPWR.t2224 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN VPWR.t2223 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5913 VPWR.t3450 a_19500_27815# a_19412_27912# VPWR.t3449 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5914 VPWR.t4591 a_17932_23111# a_17844_23208# VPWR.t2491 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5915 a_39996_2727# a_39908_2824# VGND.t3403 VGND.t3402 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5916 VPWR.t4772 a_63292_1159# a_63204_1256# VPWR.t4771 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5917 a_64412_9432# a_64324_9476# VGND.t5450 VGND.t5449 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5918 a_32268_23544# a_32180_23588# VGND.t708 VGND.t707 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5919 VPWR.t4683 _304_.B _438_.ZN VPWR.t4682 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5920 a_43356_30951# a_43268_31048# VGND.t709 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5921 _371_.A1.t6 _362_.B.t17 VPWR.t6541 VPWR.t6540 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5922 VPWR.t836 a_44632_30206# _388_.B VPWR.t835 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5923 a_1916_29383# a_1828_29480# VGND.t1905 VGND.t1904 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5924 a_64412_6296# a_64324_6340# VGND.t5855 VGND.t3471 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5925 a_21068_23544# a_20980_23588# VGND.t711 VGND.t710 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5926 uio_out[5].t6 a_20672_30301# VGND.t4867 VGND.t71 nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X5927 _325_.ZN _325_.A1.t19 a_43664_17317# VPWR.t6828 pfet_06v0 ad=0.3159p pd=1.735u as=0.44955p ps=1.955u w=1.215u l=0.5u
X5928 VGND.t6491 _287_.A1.t31 uo_out[2].t5 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X5929 VPWR.t5368 a_61836_16839# a_61748_16936# VPWR.t5367 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5930 VPWR.t5101 a_3260_29816# a_3172_29860# VPWR.t3742 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5931 a_35914_28776# _362_.B.t18 a_35710_28776# VGND.t6257 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X5932 a_58140_9432# a_58052_9476# VGND.t4715 VGND.t4714 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5933 a_47483_20569# a_45920_20523# a_46848_20893# VGND.t1975 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X5934 VGND.t802 a_41392_27165# a_41344_27209# VGND.t801 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X5935 VPWR.t5273 a_49740_12135# a_49652_12232# VPWR.t5272 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5936 VPWR.t4405 a_63068_15271# a_62980_15368# VPWR.t2676 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5937 a_64300_13703# a_64212_13800# VGND.t713 VGND.t712 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5938 VPWR.t4549 a_3260_26680# a_3172_26724# VPWR.t2185 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5939 a_50792_26344# _411_.A2.t13 _412_.B2 VPWR.t119 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5940 VGND.t3152 _398_.C _399_.A2 VGND.t3151 nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X5941 VPWR.t4923 a_9756_1592# a_9668_1636# VPWR.t4922 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5942 VPWR.t767 a_31260_16839# a_31172_16936# VPWR.t766 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5943 _399_.A1 _395_.A3 a_50196_22805# VGND.t5299 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X5944 _438_.A2 a_37472_24419# VGND.t1920 VGND.t1919 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5945 VPWR.t1380 a_66787_30600# _256_.A2.t0 VPWR.t1379 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5946 VPWR.t6326 a_46716_12135# a_46628_12232# VPWR.t2527 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5947 VPWR.t623 a_45596_30951# a_45508_31048# VPWR.t622 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5948 a_36188_2727# a_36100_2824# VGND.t715 VGND.t714 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5949 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t1035 VGND.t1034 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5950 a_45800_30345# a_45456_30301.t4 a_45012_29816# VPWR.t7059 pfet_06v0 ad=0.1791p pd=1.355u as=0.1665p ps=1.285u w=0.36u l=0.5u
X5951 a_9980_1159# a_9892_1256# VGND.t4579 VGND.t4578 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5952 VPWR.t3051 a_64412_18840# a_64324_18884# VPWR.t1721 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5953 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I VGND.t741 VGND.t740 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5954 VPWR.t6144 a_63616_31128# _251_.A1.t2 VPWR.t6143 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X5955 a_13340_1592# a_13252_1636# VGND.t514 VGND.t513 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5956 VPWR.t4337 a_50076_17272# a_49988_17316# VPWR.t4336 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5957 _272_.B1 _251_.A1.t30 a_57120_31048# VPWR.t7021 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X5958 VPWR.t4378 a_64412_15704# a_64324_15748# VPWR.t1871 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5959 a_41384_26841# a_39536_26795# a_41099_26841# VPWR.t3264 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X5960 a_54556_21543# a_54468_21640# VGND.t1852 VGND.t1851 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5961 VGND.t6619 a_42392_22825.t37 _452_.CLK.t23 VGND.t6618 nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X5962 a_32604_17272# a_32516_17316# VGND.t4984 VGND.t4983 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5963 a_51883_27508# _411_.A2.t14 _408_.ZN VGND.t114 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5964 VPWR.t4839 a_53212_15704# a_53124_15748# VPWR.t4838 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5965 a_56124_23111# a_56036_23208# VGND.t516 VGND.t515 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5966 VPWR.t4083 _454_.Q _371_.A2 VPWR.t4082 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5967 VPWR.t6411 _337_.A3.t14 _371_.A2 VPWR.t6410 pfet_06v0 ad=0.4056p pd=1.805u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5968 _399_.A2 _474_.Q a_48516_24080# VGND.t4646 nfet_06v0 ad=0.2028p pd=1.3u as=93.59999f ps=1.02u w=0.78u l=0.6u
X5969 VPWR.t4515 a_32848_29123# a_32820_29535# VPWR.t4514 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X5970 a_17168_27165# a_16796_27209# VGND.t930 VGND.t929 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X5971 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN VGND.t4724 VGND.t71 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X5972 a_5388_15271# a_5300_15368# VGND.t518 VGND.t517 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5973 VPWR.t196 _424_.A2.t14 a_50644_21640# VPWR.t195 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5974 a_34448_25597# a_34155_25273# VGND.t5693 VGND.t5692 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X5975 VPWR.t3410 a_62564_29032# _250_.C VPWR.t3409 pfet_06v0 ad=0.34437p pd=1.895u as=0.31207p ps=1.665u w=1.095u l=0.5u
X5976 a_62396_9432# a_62308_9476# VGND.t1108 VGND.t1107 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5977 a_62864_25156# _251_.A1.t31 a_61836_25515# VPWR.t7022 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X5978 VPWR.t5298 a_47612_30951# a_47524_31048# VPWR.t5297 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5979 a_5388_12135# a_5300_12232# VGND.t1543 VGND.t1542 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5980 a_60212_25156# a_59652_25640# a_60084_25640# VGND.t725 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X5981 a_19836_1592# a_19748_1636# VGND.t520 VGND.t519 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5982 VPWR.t4348 a_3260_17272# a_3172_17316# VPWR.t2179 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5983 VPWR.t6891 _448_.Q.t11 _438_.ZN VPWR.t6890 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X5984 _371_.A1.t0 _334_.A1 VPWR.t2351 VPWR.t2350 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5985 a_46044_15271# a_45956_15368# VGND.t522 VGND.t521 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5986 a_46308_20937# a_45508_20936.t7 VGND.t194 VGND.t193 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X5987 a_16140_27815# a_16052_27912# VGND.t5695 VGND.t5694 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5988 VPWR.t5304 a_15460_31048# a_15460_31048# VPWR.t5303 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5989 VPWR.t3836 _255_.I _255_.ZN VPWR.t3835 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5990 a_17484_23544# a_17396_23588# VGND.t524 VGND.t523 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X5991 VPWR.t6316 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN VPWR.t6315 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X5992 VPWR.t174 _336_.A2.t10 _337_.ZN VPWR.t173 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X5993 VPWR.t3604 a_5388_7431# a_5300_7528# VPWR.t3603 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5994 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I VPWR.t5126 VPWR.t5125 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5995 VPWR.t5686 a_21852_1159# a_21764_1256# VPWR.t5685 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5996 VPWR.t4982 a_43750_23544# a_43850_23588# VPWR.t4981 pfet_06v0 ad=0.1656p pd=1.28u as=61.19999f ps=0.7u w=0.36u l=0.5u
X5997 _397_.A2.t0 a_48104_30219# VPWR.t2438 VPWR.t2437 pfet_06v0 ad=0.3172p pd=1.74u as=0.854p ps=3.84u w=1.22u l=0.5u
X5998 a_47476_28292# _397_.A2.t17 _389_.ZN VPWR.t6504 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X5999 a_27328_25227# a_26916_25640.t7 VGND.t6476 VGND.t6475 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X6000 VPWR.t5332 a_22636_23544# a_22548_23588# VPWR.t5331 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6001 a_17372_30951# a_17284_31048# VGND.t1804 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6002 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN VGND.t2168 VGND.t2084 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6003 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I VPWR.t967 VPWR.t966 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6004 VPWR.t2298 a_1468_20408# a_1380_20452# VPWR.t2297 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6005 VPWR.t5375 a_54780_9432# a_54692_9476# VPWR.t5374 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6006 VGND.t6374 _452_.CLK.t53 a_42596_27208.t1 VGND.t6373 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X6007 _393_.ZN _389_.ZN VGND.t5132 VGND.t5131 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6008 VPWR.t5852 a_64972_12135# a_64884_12232# VPWR.t5851 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6009 a_63404_20408# a_63316_20452# VGND.t2214 VGND.t2213 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6010 a_41564_1592# a_41476_1636# VGND.t4853 VGND.t4852 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6011 VPWR.t4939 a_15580_1159# a_15492_1256# VPWR.t1629 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6012 VPWR.t4731 a_48284_15271# a_48196_15368# VPWR.t1631 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6013 a_33708_22505# _316_.ZN a_33584_22137# VPWR.t5470 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X6014 a_31484_26680# a_31396_26724# VGND.t3496 VGND.t3495 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6015 a_65532_1592# a_65444_1636# VGND.t1110 VGND.t1109 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6016 VPWR.t3726 a_53772_12135# a_53684_12232# VPWR.t3725 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6017 a_16028_1592# a_15940_1636# VGND.t830 VGND.t829 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6018 _274_.A2 _258_.I a_56596_29861# VPWR.t322 pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X6019 a_39548_1159# a_39460_1256# VGND.t4388 VGND.t4387 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6020 VPWR.t4877 a_35740_25112# a_35652_25156# VPWR.t4876 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6021 VPWR.t884 a_66204_8999# a_66116_9096# VPWR.t883 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6022 a_34620_1159# a_34532_1256# VGND.t2207 VGND.t2206 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6023 a_43666_21812# a_42982_21730# VPWR.t5439 VPWR.t5438 pfet_06v0 ad=61.19999f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X6024 a_52660_24072# _424_.A2.t15 a_52452_24072# VGND.t189 nfet_06v0 ad=58.39999f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X6025 a_44704_18191# a_42484_18183.t5 a_44459_18559# VGND.t6732 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6026 VPWR.t5428 a_46492_17272# a_46404_17316# VPWR.t5427 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6027 VPWR.t3019 _305_.A2 a_45396_22020# VPWR.t3018 pfet_06v0 ad=0.4818p pd=3.07u as=0.4599p ps=1.935u w=1.095u l=0.5u
X6028 a_45800_30345# a_45416_29885# a_45012_29816# VGND.t137 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6029 VPWR.t5434 a_21516_25112# a_21428_25156# VPWR.t5433 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6030 VPWR.t4572 a_35292_17272# a_35204_17316# VPWR.t4571 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6031 _441_.A2 _447_.Q.t14 VPWR.t6590 VPWR.t6589 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X6032 VPWR.t2556 _349_.A4 _371_.A2 VPWR.t2555 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X6033 VPWR.t4756 a_29020_1592# a_28932_1636# VPWR.t4262 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6034 a_49628_15704# a_49540_15748# VGND.t941 VGND.t940 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6035 VPWR.t561 a_13788_2727# a_13700_2824# VPWR.t560 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6036 VPWR.t563 a_34732_18407# a_34644_18504# VPWR.t562 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6037 a_48068_21236# _419_.A4 VGND.t3980 VGND.t3979 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6038 a_37980_2727# a_37892_2824# VGND.t2663 VGND.t2662 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6039 a_53660_12568# a_53572_12612# VGND.t3869 VGND.t3868 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6040 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I VGND.t5758 VGND.t5757 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6041 VGND.t1244 vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t1243 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6042 a_42392_22825.t1 clkbuf_1_0__f_clk.I.t55 VPWR.t268 VPWR.t267 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X6043 VGND.t2665 a_47297_25596# _381_.A2.t1 VGND.t2664 nfet_06v0 ad=0.2288p pd=1.58u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6044 VPWR.t2217 a_1468_14136# a_1380_14180# VPWR.t2216 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6045 VPWR.t5871 a_31708_18407# a_31620_18504# VPWR.t3511 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6046 a_38808_27967# a_36960_27912# a_38523_27967# VPWR.t5487 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X6047 VPWR.t2003 a_1468_11000# a_1380_11044# VPWR.t1897 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6048 a_61948_27815# a_61860_27912# VGND.t1836 VGND.t1835 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6049 VGND.t2053 a_45012_29816# a_44632_30206# VGND.t2052 nfet_06v0 ad=0.142p pd=1.14u as=0.176p ps=1.68u w=0.4u l=0.6u
X6050 a_45820_18840# a_45732_18884# VGND.t2389 VGND.t2388 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6051 VGND.t6156 _451_.Q.t10 _260_.A2 VGND.t6155 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X6052 VPWR.t2807 a_48508_1159# a_48420_1256# VPWR.t2194 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6053 a_14796_28248# a_14708_28292# VGND.t4023 VGND.t4022 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6054 a_40444_2727# a_40356_2824# VGND.t2669 VGND.t2668 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6055 _359_.ZN _460_.Q a_34516_25940# VGND.t3324 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6056 a_61276_15271# a_61188_15368# VGND.t2671 VGND.t2670 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6057 VPWR.t4503 a_7740_1592# a_7652_1636# VPWR.t4502 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6058 a_67100_1159# a_67012_1256# VGND.t2673 VGND.t2672 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6059 a_54892_19975# a_54804_20072# VGND.t2675 VGND.t2674 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6060 VPWR.t1233 a_29804_30951# a_29716_31048# VPWR.t1232 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6061 VPWR.t1235 a_62396_26247# a_62308_26344# VPWR.t1234 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6062 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I VPWR.t4509 VPWR.t4508 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6063 VPWR.t2187 a_2812_6296# a_2724_6340# VPWR.t780 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6064 a_34172_2727# a_34084_2824# VGND.t2676 VGND.t892 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6065 VGND.t4967 a_60401_30300# _255_.I VGND.t71 nfet_06v0 ad=0.2288p pd=1.58u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6066 VPWR.t5076 a_4156_9432# a_4068_9476# VPWR.t3188 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6067 VGND.t2686 vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I VGND.t2685 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6068 vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN VGND.t4007 VGND.t4006 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6069 a_40668_19975# a_40580_20072# VGND.t2678 VGND.t2677 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6070 a_58140_2727# a_58052_2824# VGND.t849 VGND.t848 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6071 VGND.t6100 a_52400_25987.t6 a_53772_26031# VGND.t6099 nfet_06v0 ad=0.1584p pd=1.6u as=43.2f ps=0.6u w=0.36u l=0.6u
X6072 VPWR.t4659 a_2812_3160# a_2724_3204# VPWR.t1296 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6073 a_23084_25112# a_22996_25156# VGND.t5317 VGND.t5316 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6074 VPWR.t5723 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t5722 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6075 a_42896_18504# a_42484_18183.t6 VGND.t6734 VGND.t6733 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X6076 VPWR.t4301 a_33276_1592# a_33188_1636# VPWR.t4300 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6077 a_63180_16839# a_63092_16936# VGND.t851 VGND.t850 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6078 uo_out[1].t8 _293_.A2 VGND.t5699 VGND.t5698 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X6079 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN VPWR.t4869 VPWR.t4868 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6080 a_41048_29816.t0 vgaringosc.workerclkbuff_notouch_.I.t9 VPWR.t6705 VPWR.t6704 pfet_06v0 ad=0.2952p pd=1.54u as=0.367p ps=1.92u w=0.82u l=0.5u
X6081 VPWR.t4440 a_57244_1592# a_57156_1636# VPWR.t4439 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6082 a_23084_21976# a_22996_22020# VGND.t2680 VGND.t2679 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6083 VPWR.t4398 a_26720_30301# a_26712_29977# VPWR.t4397 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X6084 a_52640_29860# _474_.CLK.t51 VPWR.t6761 VPWR.t6760 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6085 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I _241_.I0 VPWR.t3879 VPWR.t3878 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6086 a_17168_27165# a_16796_27209# VPWR.t951 VPWR.t950 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X6087 a_38316_16839# a_38228_16936# VGND.t853 VGND.t852 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6088 a_3260_15271# a_3172_15368# VGND.t855 VGND.t854 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6089 a_35060_20569# a_33748_20936.t4 a_34716_20937# VPWR.t49 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X6090 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].I VGND.t5047 VGND.t5046 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6091 a_26220_20408# a_26132_20452# VGND.t3601 VGND.t3600 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6092 VGND.t4866 a_20672_30301# uio_out[5].t5 VGND.t71 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X6093 VPWR.t2309 a_16140_20408# a_16052_20452# VPWR.t2308 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6094 a_3260_12135# a_3172_12232# VGND.t2708 VGND.t2707 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6095 VPWR.t2128 a_17932_25112# a_17844_25156# VPWR.t2127 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6096 VPWR.t4575 a_46268_12568# a_46180_12612# VPWR.t3385 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6097 VPWR.t6161 a_64860_18840# a_64772_18884# VPWR.t2247 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6098 VGND.t4383 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN VGND.t4382 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6099 VPWR.t6142 a_63616_31128# _251_.A1.t1 VPWR.t6141 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6100 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I VGND.t3192 VGND.t3191 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6101 _452_.Q.t3 a_40040_17675# VGND.t5088 VGND.t5087 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6102 VPWR.t4626 a_64860_15704# a_64772_15748# VPWR.t4625 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6103 VPWR.t4628 a_5052_23544# a_4964_23588# VPWR.t4627 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6104 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I VGND.t3131 VGND.t3130 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6105 VPWR.t1906 a_47776_20893# a_47768_20569# VPWR.t1905 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X6106 a_23532_23544# a_23444_23588# VGND.t334 VGND.t333 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6107 VGND.t2083 vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I VGND.t2082 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6108 a_59820_14136# a_59732_14180# VGND.t3641 VGND.t3640 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6109 VPWR.t4736 a_53660_15704# a_53572_15748# VPWR.t387 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6110 a_36432_19325# a_36060_19369# VPWR.t1695 VPWR.t1694 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X6111 VPWR.t2026 a_26220_21976# a_26132_22020# VPWR.t2025 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6112 a_56572_23111# a_56484_23208# VGND.t857 VGND.t856 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6113 a_64748_23111# a_64660_23208# VGND.t56 VGND.t55 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6114 VGND.t6296 _350_.A2.t27 a_30128_27508# VGND.t6295 nfet_06v0 ad=0.2132p pd=1.34u as=98.39999f ps=1.06u w=0.82u l=0.6u
X6115 VPWR.t5689 a_65532_15271# a_65444_15368# VPWR.t5688 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6116 VPWR.t5744 a_31260_18840# a_31172_18884# VPWR.t2963 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6117 VGND.t2611 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I VGND.t2610 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6118 VPWR.t4390 a_18760_29032# a_18264_29480# VPWR.t4389 pfet_06v0 ad=0.4005p pd=2.12u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6119 VGND.t5245 a_49492_18840# a_48888_19243# VGND.t5244 nfet_06v0 ad=0.142p pd=1.14u as=0.176p ps=1.68u w=0.4u l=0.6u
X6120 a_42161_24776# _260_.ZN hold2.I VPWR.t3623 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X6121 a_62396_2727# a_62308_2824# VGND.t58 VGND.t57 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6122 VPWR.t1837 a_46716_14136# a_46628_14180# VPWR.t348 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6123 VPWR.t1564 a_41900_16839# a_41812_16936# VPWR.t1563 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6124 VGND.t5806 vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t5227 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6125 a_33060_31048# _290_.ZN VPWR.t1201 VPWR.t1200 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X6126 VPWR.t4271 a_31260_15704# a_31172_15748# VPWR.t1569 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6127 _264_.B _260_.A1 a_40676_25640# VGND.t3767 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6128 VPWR.t1418 a_60380_11000# a_60292_11044# VPWR.t1417 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6129 a_41600_19376# _325_.A2.t10 VGND.t6126 VGND.t6125 nfet_06v0 ad=79.8f pd=0.8u as=0.2424p ps=1.635u w=0.38u l=0.6u
X6130 a_50196_21640# _417_.Z VPWR.t5392 VPWR.t5391 pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X6131 VPWR.t1420 a_46716_11000# a_46628_11044# VPWR.t1419 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6132 a_35723_20569# a_34160_20523# a_35088_20893# VGND.t2763 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6133 VGND.t1179 _343_.A2 _345_.A2 VGND.t1178 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X6134 VPWR.t451 a_43132_15271# a_43044_15368# VPWR.t450 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6135 a_46492_15271# a_46404_15368# VGND.t60 VGND.t59 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6136 a_31124_25156# _355_.C.t15 _459_.D VPWR.t6676 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6137 a_52744_26031# a_52360_26355# a_51956_26183# VGND.t3135 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6138 a_65868_12135# a_65780_12232# VGND.t2756 VGND.t2755 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6139 VGND.t6704 _251_.A1.t32 a_59652_25640# VGND.t6703 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6140 a_54668_12135# a_54580_12232# VGND.t5960 VGND.t5959 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6141 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN VGND.t5573 VGND.t5572 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6142 VPWR.t544 a_14460_30951# a_14372_31048# VPWR.t543 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6143 VPWR.t546 a_22636_30951# a_22548_31048# VPWR.t545 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6144 a_1020_18407# a_932_18504# VGND.t62 VGND.t61 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6145 a_3708_26247# a_3620_26344# VGND.t64 VGND.t63 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6146 a_13788_1159# a_13700_1256# VGND.t2854 VGND.t2853 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6147 VPWR.t6190 a_22188_29383# a_22100_29480# VPWR.t6189 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6148 VPWR.t3155 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I VPWR.t3154 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6149 _421_.B _416_.A3 a_47524_22021# VPWR.t4465 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X6150 a_50188_10567# a_50100_10664# VGND.t66 VGND.t65 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6151 a_16700_2727# a_16612_2824# VGND.t68 VGND.t67 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6152 VPWR.t955 a_11772_2727# a_11684_2824# VPWR.t954 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6153 a_43452_18191# _450_.D a_43284_18191# VGND.t3711 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X6154 a_34160_20523# a_33748_20936.t5 VPWR.t51 VPWR.t50 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X6155 a_3708_23111# a_3620_23208# VGND.t6764 VGND.t2935 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6156 a_41040_17801# a_40040_17675# VGND.t5086 VGND.t5085 nfet_06v0 ad=43.2f pd=0.6u as=0.142p ps=1.14u w=0.36u l=0.6u
X6157 _241_.Z a_56964_26724# VPWR.t5741 VPWR.t5740 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X6158 VPWR.t2102 a_35740_2727# a_35652_2824# VPWR.t2101 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6159 VPWR.t2254 a_50748_20408# a_50660_20452# VPWR.t2253 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6160 a_53548_16839# a_53460_16936# VGND.t6766 VGND.t6765 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6161 VPWR.t6300 a_28908_20408# a_28820_20452# VPWR.t6299 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6162 _460_.Q a_34448_25597# VGND.t3729 VGND.t3728 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6163 VPWR.t3549 a_54444_19975# a_54356_20072# VPWR.t3548 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6164 _435_.A3 _304_.B a_43253_25940# VGND.t4526 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6165 _371_.ZN _371_.A3 VGND.t955 VGND.t954 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X6166 VPWR.t2328 a_31372_20408# a_31284_20452# VPWR.t2327 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6167 a_60416_25156# a_59652_25640# a_60212_25156# VPWR.t737 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6168 a_43888_19204# a_43440_19325.t5 a_44300_19001# VPWR.t6462 pfet_06v0 ad=0.1872p pd=1.4u as=43.2f ps=0.6u w=0.36u l=0.5u
X6169 VPWR.t6152 a_4156_21543# a_4068_21640# VPWR.t2007 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6170 VPWR.t684 a_58364_25112# a_58276_25156# VPWR.t683 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6171 VPWR.t2106 a_36076_16839# a_35988_16936# VPWR.t2105 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6172 VPWR.t5499 a_21964_25112# a_21876_25156# VPWR.t5498 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6173 a_39587_24372# _430_.ZN VGND.t4672 VGND.t4671 nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6174 _379_.Z _379_.A2 a_18264_29480# VPWR.t2733 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6175 a_63404_10567# a_63316_10664# VGND.t6768 VGND.t6767 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6176 a_34548_20937# a_33748_20936.t6 VGND.t43 VGND.t42 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X6177 a_4156_4295# a_4068_4392# VGND.t5860 VGND.t2540 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6178 VPWR.t5727 a_16252_1159# a_16164_1256# VPWR.t5726 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6179 a_24304_29480# _340_.ZN a_24100_29480# VPWR.t1158 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6180 VPWR.t2096 a_57132_10567# a_57044_10664# VPWR.t2095 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6181 uio_out[6].t0 a_19328_28733# VPWR.t6041 VPWR.t6040 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6182 a_37772_19759# _319_.A3 VGND.t2570 VGND.t2569 nfet_06v0 ad=58.39999f pd=0.685u as=0.23405p ps=1.555u w=0.365u l=0.6u
X6183 a_2812_20408# a_2724_20452# VGND.t4097 VGND.t2208 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6184 a_40452_22504# _448_.Q.t12 a_39796_22504# VGND.t6578 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6185 VPWR.t2010 a_61948_14136# a_61860_14180# VPWR.t2009 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6186 a_3708_16839# a_3620_16936# VGND.t6769 VGND.t1877 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6187 a_28928_29123# a_28556_29167# VGND.t1533 VGND.t1532 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X6188 a_41340_1159# a_41252_1256# VGND.t407 VGND.t406 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6189 a_33052_18407# a_32964_18504# VGND.t6770 VGND.t4883 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6190 VPWR.t5845 a_58028_18840# a_57940_18884# VPWR.t5844 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6191 a_14796_24679# a_14708_24776# VGND.t6771 VGND.t1879 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6192 VPWR.t4364 a_49180_9432# a_49092_9476# VPWR.t4363 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6193 a_37536_29167# a_35316_29159.t4 a_37291_29535# VGND.t6739 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6194 a_20956_2727# a_20868_2824# VGND.t6773 VGND.t6772 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6195 VPWR.t2094 a_31260_1592# a_31172_1636# VPWR.t2093 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6196 a_65084_12568# a_64996_12612# VGND.t4611 VGND.t4610 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6197 VPWR.t2193 a_61948_11000# a_61860_11044# VPWR.t2192 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6198 VPWR.t3187 a_50748_14136# a_50660_14180# VPWR.t3186 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6199 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN VPWR.t3572 VPWR.t3571 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6200 a_14796_21543# a_14708_21640# VGND.t1579 VGND.t1578 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6201 VPWR.t4096 a_58588_21543# a_58500_21640# VPWR.t4095 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6202 a_51252_19001# _474_.D a_50384_19204# VPWR.t2673 pfet_06v0 ad=54f pd=0.66u as=0.1872p ps=1.4u w=0.36u l=0.5u
X6203 a_47768_20569# a_45920_20523# a_47483_20569# VPWR.t2076 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X6204 VPWR.t1640 vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I VPWR.t1639 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6205 VPWR.t3444 a_50748_11000# a_50660_11044# VPWR.t3443 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6206 a_43440_26841# a_43008_26795# VPWR.t6007 VPWR.t6006 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X6207 a_36160_29535# a_35728_29480# VPWR.t669 VPWR.t668 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X6208 a_14684_2727# a_14596_2824# VGND.t6774 VGND.t1887 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6209 VPWR.t2133 a_67212_12135# a_67124_12232# VPWR.t2132 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6210 VPWR.t6212 a_4156_12135# a_4068_12232# VPWR.t2233 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6211 _437_.A1.t0 a_38816_27555# VPWR.t5806 VPWR.t5805 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6212 VPWR.t1299 a_2812_21976# a_2724_22020# VPWR.t1298 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6213 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN VGND.t5424 VGND.t5423 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6214 VGND.t5598 _301_.Z a_39172_22504# VGND.t5597 nfet_06v0 ad=0.226p pd=1.515u as=88.2f ps=0.84u w=0.42u l=0.6u
X6215 _284_.ZN.t14 _304_.B a_44948_25156# VPWR.t4681 pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X6216 VPWR.t2084 a_38428_2727# a_38340_2824# VPWR.t2083 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6217 VPWR.t6089 a_56012_12135# a_55924_12232# VPWR.t6088 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6218 a_29348_25940# _336_.A2.t11 a_29164_25940# VGND.t167 nfet_06v0 ad=0.1148p pd=1.1u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6219 VPWR.t390 a_13788_1592# a_13700_1636# VPWR.t389 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6220 uio_out[7].t4 a_18096_27165# VGND.t388 VGND.t387 nfet_06v0 ad=0.2119p pd=1.335u as=0.2608p ps=1.455u w=0.815u l=0.6u
X6221 VPWR.t396 a_37756_1592# a_37668_1636# VPWR.t395 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6222 a_65308_7431# a_65220_7528# VGND.t6795 VGND.t2947 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6223 VPWR.t5426 a_49492_18840# a_48888_19243# VPWR.t5425 pfet_06v0 ad=0.23p pd=1.54u as=0.352p ps=2.48u w=0.8u l=0.5u
X6224 VPWR.t3994 a_31708_17272# a_31620_17316# VPWR.t1934 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6225 a_2812_14136# a_2724_14180# VGND.t3762 VGND.t2461 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6226 _324_.B.t8 _304_.B a_42168_22504# VGND.t4525 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6227 VPWR.t4944 a_19276_23544# a_19188_23588# VPWR.t4943 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6228 a_38764_16839# a_38676_16936# VGND.t6797 VGND.t6796 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6229 a_2812_11000# a_2724_11044# VGND.t3808 VGND.t2896 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6230 a_40220_26247# a_40132_26344# VGND.t6799 VGND.t6798 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6231 VPWR.t665 a_18716_24679# a_18628_24776# VPWR.t664 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6232 uo_out[2].t11 _288_.ZN.t9 VGND.t6066 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X6233 a_60380_2727# a_60292_2824# VGND.t6800 VGND.t805 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6234 a_64860_9432# a_64772_9476# VGND.t1389 VGND.t1388 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6235 VPWR.t6027 _390_.ZN _392_.A2 VPWR.t6026 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X6236 VPWR.t706 a_64860_26247# a_64772_26344# VPWR.t705 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6237 a_49056_29977# a_48104_30219# VPWR.t2436 VPWR.t2435 pfet_06v0 ad=50.4f pd=0.64u as=0.23p ps=1.54u w=0.36u l=0.5u
X6238 a_52540_15271# a_52452_15368# VGND.t6801 VGND.t497 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6239 VGND.t222 _330_.A1.t21 _319_.ZN VGND.t221 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X6240 a_4156_27815# a_4068_27912# VGND.t1575 VGND.t1574 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6241 a_59820_10567# a_59732_10664# VGND.t6803 VGND.t6802 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6242 a_64188_1592# a_64100_1636# VGND.t981 VGND.t980 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6243 a_64860_6296# a_64772_6340# VGND.t2700 VGND.t2699 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6244 a_35728_29480# a_35316_29159.t5 VGND.t6741 VGND.t6740 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X6245 a_17596_1159# a_17508_1256# VGND.t2837 VGND.t2836 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6246 a_23980_23544# a_23892_23588# VGND.t4340 VGND.t4339 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6247 a_60716_12135# a_60628_12232# VGND.t5347 VGND.t5346 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6248 a_3260_3160# a_3172_3204# VGND.t3295 VGND.t3294 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6249 VPWR.t6592 _447_.Q.t15 a_35816_21192# VPWR.t6591 pfet_06v0 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X6250 VPWR.t430 a_4940_24679# a_4852_24776# VPWR.t429 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6251 a_67237_31198# a_67117_30600# VPWR.t3326 VPWR.t3325 pfet_06v0 ad=61.19999f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X6252 VGND.t6785 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN VGND.t6784 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6253 _241_.I0 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I VGND.t3356 VGND.t3355 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6254 VPWR.t4951 a_27004_21543# a_26916_21640# VPWR.t4950 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6255 a_34032_22505# a_33152_22091# a_33708_22505# VGND.t1395 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X6256 a_29371_30644# _350_.A1.t11 _340_.A2 VGND.t34 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6257 VPWR.t739 a_65980_15271# a_65892_15368# VPWR.t738 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6258 a_42610_21812# a_42154_21236# VPWR.t2506 VPWR.t2505 pfet_06v0 ad=61.19999f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X6259 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN VGND.t4960 VGND.t4959 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6260 VGND.t6046 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN VGND.t6045 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6261 VPWR.t2402 a_1916_24679# a_1828_24776# VPWR.t1397 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6262 VPWR.t2278 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN VPWR.t2277 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6263 a_65308_19975# a_65220_20072# VGND.t6804 VGND.t2903 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6264 _336_.Z a_28820_24072# VPWR.t3849 VPWR.t3848 pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X6265 a_42460_17801# _452_.D a_41536_17636# VGND.t2502 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X6266 a_44160_29123# a_43788_29167# VGND.t4931 VGND.t4930 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X6267 VPWR.t2408 a_61164_10567# a_61076_10664# VPWR.t2407 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6268 a_46044_30951# a_45956_31048# VGND.t6805 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6269 VPWR.t4298 a_59932_12568# a_59844_12612# VPWR.t4297 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6270 _375_.Z a_20003_29611# VGND.t5809 VGND.t5808 nfet_06v0 ad=0.3608p pd=2.52u as=0.2288p ps=1.58u w=0.82u l=0.6u
X6271 a_46620_22504# _402_.A1.t21 _402_.ZN VGND.t6440 nfet_06v0 ad=0.1312p pd=1.14u as=0.2569p ps=1.56u w=0.82u l=0.6u
X6272 a_63180_26680# a_63092_26724# VGND.t4820 VGND.t4819 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6273 VPWR.t700 a_43580_15271# a_43492_15368# VPWR.t699 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6274 a_33140_29860# _362_.ZN a_32916_29860# VPWR.t5777 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6275 a_61052_9432# a_60964_9476# VGND.t2216 VGND.t2215 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6276 VPWR.t2412 a_64524_16839# a_64436_16936# VPWR.t2411 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6277 VGND.t1684 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN VGND.t1683 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6278 VPWR.t702 a_20060_23111# a_19972_23208# VPWR.t701 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6279 a_3260_28248# a_3172_28292# VGND.t2768 VGND.t2767 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6280 _424_.B1.t5 _324_.C.t30 a_50532_24072# VGND.t6511 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6281 VPWR.t2414 a_1468_16839# a_1380_16936# VPWR.t2413 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6282 _304_.ZN.t5 _304_.A1.t11 a_42252_20936# VGND.t6319 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6283 _247_.B _252_.B a_59620_27208# VGND.t768 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6284 a_17803_26841# a_15828_27208.t7 a_17168_27165# VPWR.t6385 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X6285 vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN VGND.t2957 VGND.t2956 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6286 a_5388_4295# a_5300_4392# VGND.t3687 VGND.t3686 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6287 _447_.Q.t1 a_36016_20893# VGND.t1674 VGND.t1673 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6288 VPWR.t2631 a_7068_2727# a_6980_2824# VPWR.t2630 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6289 a_47259_20127# a_45696_20072# a_46624_19715# VGND.t2470 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6290 VPWR.t3252 a_54040_22366# _281_.A1 VPWR.t3251 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6291 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I VGND.t2609 VGND.t2608 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6292 a_58588_1159# a_58500_1256# VGND.t5043 VGND.t5042 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6293 a_33808_23705# a_33376_23659# VPWR.t1912 VPWR.t1911 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X6294 VPWR.t4402 a_6396_1592# a_6308_1636# VPWR.t4401 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6295 a_53660_1159# a_53572_1256# VGND.t5943 VGND.t5942 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6296 a_44924_15704# a_44836_15748# VGND.t4351 VGND.t4350 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6297 a_5388_24679# a_5300_24776# VGND.t6807 VGND.t6806 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6298 a_67548_9432# a_67460_9476# VGND.t3857 VGND.t3856 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6299 VPWR.t5370 a_4940_15271# a_4852_15368# VPWR.t5369 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6300 VPWR.t1675 a_67100_18840# a_67012_18884# VPWR.t1674 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6301 a_28208_25641# a_27328_25227# a_27884_25641# VGND.t6027 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X6302 a_48529_22460# _475_.Q a_48921_22020# VPWR.t4998 pfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.5u
X6303 VPWR.t4548 a_1468_6296# a_1380_6340# VPWR.t3744 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6304 a_40220_1592# a_40132_1636# VGND.t2845 VGND.t2844 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6305 a_53996_16839# a_53908_16936# VGND.t6809 VGND.t6808 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6306 a_52660_21640# _427_.B2 VPWR.t3933 VPWR.t3932 pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X6307 a_5388_21543# a_5300_21640# VGND.t1457 VGND.t1456 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6308 a_67548_6296# a_67460_6340# VGND.t4058 VGND.t1321 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6309 a_17148_29816# a_17060_29860# VGND.t6810 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6310 VPWR.t5371 a_1916_15271# a_1828_15368# VPWR.t2039 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6311 VPWR.t619 a_67100_15704# a_67012_15748# VPWR.t618 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6312 a_37067_19001# a_35092_19368.t7 a_36432_19325# VPWR.t93 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X6313 VGND.t6812 a_31088_30301# a_31040_30345# VGND.t137 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X6314 VPWR.t2815 a_54892_19975# a_54804_20072# VPWR.t2814 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6315 VPWR.t2635 a_52204_18407# a_52116_18504# VPWR.t2634 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6316 a_44948_22020# _305_.A2 VPWR.t3017 VPWR.t3016 pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X6317 VPWR.t3178 a_1468_3160# a_1380_3204# VPWR.t529 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6318 a_26108_1159# a_26020_1256# VGND.t6814 VGND.t6813 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6319 a_38784_22504# _447_.Q.t16 a_38576_22504# VGND.t6308 nfet_06v0 ad=67.2f pd=0.74u as=0.1848p ps=1.72u w=0.42u l=0.6u
X6320 VPWR.t2416 a_22748_24679# a_22660_24776# VPWR.t2415 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6321 VGND.t4645 _474_.Q a_47297_25596# VGND.t4644 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6322 a_39268_18840# _327_.Z a_39648_19435# VGND.t5364 nfet_06v0 ad=0.1584p pd=1.6u as=57.59999f ps=0.68u w=0.36u l=0.6u
X6323 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN VPWR.t4607 VPWR.t4606 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6324 VGND.t2895 a_25232_27165# a_25184_27209# VGND.t2894 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X6325 VPWR.t6815 _324_.C.t31 _416_.A1.t0 VPWR.t6814 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6326 VPWR.t4538 a_55788_25112# a_55700_25156# VPWR.t4537 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6327 a_28756_25940# _336_.A2.t12 a_28552_25940# VGND.t168 nfet_06v0 ad=0.1312p pd=1.14u as=0.1722p ps=1.24u w=0.82u l=0.6u
X6328 a_43440_19325.t1 _452_.CLK.t54 VGND.t6376 VGND.t6375 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X6329 a_3260_18840# a_3172_18884# VGND.t5214 VGND.t5213 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6330 VPWR.t2818 a_40668_19975# a_40580_20072# VPWR.t1831 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6331 _474_.CLK.t25 a_48272_25156.t39 VGND.t6286 VGND.t6285 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X6332 a_63852_10567# a_63764_10664# VGND.t6816 VGND.t6815 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6333 a_46624_19715# a_46252_19759# VPWR.t1919 VPWR.t1918 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X6334 VPWR.t4377 a_59932_9432# a_59844_9476# VPWR.t4376 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6335 a_47164_13703# a_47076_13800# VGND.t1822 VGND.t1732 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6336 a_54088_22895# a_53744_22851.t6 a_53300_23047# VPWR.t27 pfet_06v0 ad=0.1791p pd=1.355u as=0.1665p ps=1.285u w=0.36u l=0.5u
X6337 VGND.t136 _417_.A2.t11 a_49672_19668# VGND.t135 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6338 a_25936_25597# a_25643_25273# VGND.t3924 VGND.t3923 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X6339 VPWR.t2424 a_12444_2727# a_12356_2824# VPWR.t2423 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6340 a_42460_20452# _303_.ZN VPWR.t2950 VPWR.t2949 pfet_06v0 ad=0.4599p pd=1.935u as=0.4818p ps=3.07u w=1.095u l=0.5u
X6341 a_14236_29383# a_14148_29480# VGND.t5543 VGND.t5542 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6342 VPWR.t2426 a_57580_10567# a_57492_10664# VPWR.t2425 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6343 a_44276_20072# _325_.A1.t20 _328_.A2 VPWR.t6829 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X6344 a_31708_15271# a_31620_15368# VGND.t6818 VGND.t6817 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6345 a_68108_12135# a_68020_12232# VGND.t3173 VGND.t3172 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6346 VPWR.t1002 a_31036_21543# a_30948_21640# VPWR.t1001 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6347 a_65980_1592# a_65892_1636# VGND.t4801 VGND.t4800 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6348 vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN VGND.t2724 VGND.t2723 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6349 a_41392_27165# a_41099_26841# VGND.t5280 VGND.t5279 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X6350 a_27004_27815# a_26916_27912# VGND.t1564 VGND.t1563 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6351 a_3708_8999# a_3620_9096# VGND.t6073 VGND.t5639 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6352 _460_.D _360_.ZN VPWR.t6214 VPWR.t6213 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6353 VPWR.t579 a_66652_8999# a_66564_9096# VPWR.t578 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6354 VPWR.t1628 a_58476_18840# a_58388_18884# VPWR.t1627 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6355 VGND.t2016 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN VGND.t2015 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6356 VGND.t2020 vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I VGND.t2019 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6357 a_39324_19975# a_39236_20072# VGND.t6075 VGND.t6074 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6358 VPWR.t1154 a_10428_29383# a_10340_29480# VPWR.t1153 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6359 a_3708_5863# a_3620_5960# VGND.t1131 VGND.t1130 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6360 VPWR.t583 a_32828_23111# a_32740_23208# VPWR.t582 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6361 VPWR.t6567 a_48272_25156.t40 _474_.CLK.t26 VPWR.t6566 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6362 VGND.t1504 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t1503 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6363 a_26746_26344# _355_.C.t16 _457_.D VPWR.t6677 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6364 a_44812_16839# a_44724_16936# VGND.t6077 VGND.t6076 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6365 VPWR.t1060 a_49740_16839# a_49652_16936# VPWR.t1059 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6366 VPWR.t5300 a_25324_23544# a_25236_23588# VPWR.t5299 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6367 VGND.t5516 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t2169 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6368 VPWR.t3802 a_67212_20408# a_67124_20452# VPWR.t3801 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6369 a_34708_29860# _294_.ZN.t8 VPWR.t150 VPWR.t149 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X6370 VPWR.t3212 a_4156_20408# a_4068_20452# VPWR.t2338 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6371 _395_.A2 a_49764_26724# VPWR.t1022 VPWR.t1021 pfet_06v0 ad=0.5368p pd=3.32u as=0.389p ps=2.02u w=1.22u l=0.5u
X6372 a_24988_23111# a_24900_23208# VGND.t6079 VGND.t6078 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6373 a_48988_27508# _397_.A2.t18 _411_.A2.t2 VGND.t6227 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6374 VPWR.t4190 a_67660_12135# a_67572_12232# VPWR.t4189 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6375 VPWR.t3602 a_33948_15271# a_33860_15368# VPWR.t2011 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6376 a_47297_25596# _474_.Q a_47689_25156# VPWR.t4794 pfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.5u
X6377 a_49013_22805# _399_.A2 VGND.t1403 VGND.t1402 nfet_06v0 ad=92.99999f pd=1.015u as=0.23975p ps=1.475u w=0.775u l=0.6u
X6378 VPWR.t6963 _452_.Q.t18 a_41488_24072# VPWR.t6962 pfet_06v0 ad=0.395p pd=2.02u as=0.156p ps=1.12u w=0.6u l=0.5u
X6379 VPWR.t1094 a_56124_9432# a_56036_9476# VPWR.t1093 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6380 a_38852_18884# _327_.Z VPWR.t5566 VPWR.t5565 pfet_06v0 ad=0.55297p pd=2.105u as=0.4818p ps=3.07u w=1.095u l=0.5u
X6381 _274_.A3 _474_.CLK.t52 VGND.t6462 VGND.t108 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X6382 VPWR.t1162 _373_.A2 a_26970_29480# VPWR.t1161 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X6383 VPWR.t4009 a_56460_12135# a_56372_12232# VPWR.t4008 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6384 a_47028_18884# _416_.A1.t12 _416_.ZN VPWR.t204 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6385 VGND.t205 _416_.A1.t13 _442_.ZN VGND.t204 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X6386 _384_.A3.t6 _474_.Q VPWR.t4793 VPWR.t4792 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X6387 a_41099_26841# a_39536_26795# a_40464_27165# VGND.t3117 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6388 a_2812_10567# a_2724_10664# VGND.t6080 VGND.t2586 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6389 VGND.t1946 a_37584_29123# _334_.A1 VGND.t1945 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6390 a_62172_1592# a_62084_1636# VGND.t3506 VGND.t3505 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6391 VPWR.t3453 a_1916_4295# a_1828_4392# VPWR.t1362 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6392 a_63404_23544# a_63316_23588# VGND.t5035 VGND.t5034 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6393 VPWR.t5334 a_49180_17272# a_49092_17316# VPWR.t5333 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6394 VGND.t3429 _371_.A2 _352_.A2.t5 VGND.t3428 nfet_06v0 ad=0.2405p pd=1.52u as=0.1326p ps=1.03u w=0.51u l=0.6u
X6395 a_63105_28293# _248_.B1 VPWR.t1215 VPWR.t1214 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X6396 a_31116_26020# _336_.Z a_30932_26020# VGND.t4411 nfet_06v0 ad=79.8f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X6397 a_3260_30951# a_3172_31048# VGND.t336 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6398 a_20928_26399# a_20496_26344# VPWR.t4817 VPWR.t4816 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X6399 a_32800_29167# a_31920_29480# a_32476_29167# VGND.t3139 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X6400 VPWR.t4730 a_1916_1159# a_1828_1256# VPWR.t1300 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6401 a_40892_2727# a_40804_2824# VGND.t6082 VGND.t6081 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6402 VPWR.t3312 a_48956_1159# a_48868_1256# VPWR.t3085 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6403 a_31068_28292# _371_.A1.t18 _350_.A2.t14 VPWR.t6513 pfet_06v0 ad=0.3942p pd=1.815u as=0.2847p ps=1.615u w=1.095u l=0.5u
X6404 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t1606 VGND.t1605 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6405 _431_.A3 _438_.A2 a_38752_26344# VPWR.t5117 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X6406 a_50524_17272# a_50436_17316# VGND.t3819 VGND.t3818 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6407 VGND.t4934 a_25008_25597# a_24960_25641# VGND.t4933 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X6408 a_3708_26680# a_3620_26724# VGND.t3457 VGND.t3009 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6409 VPWR.t5033 a_64636_2727# a_64548_2824# VPWR.t5032 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6410 a_60656_29612# _252_.ZN VPWR.t6271 VPWR.t6270 pfet_06v0 ad=0.224p pd=1.36u as=0.389p ps=2.02u w=0.56u l=0.5u
X6411 a_1468_12568# a_1380_12612# VGND.t1765 VGND.t1764 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6412 a_59744_30352# _255_.I VGND.t3683 VGND.t3682 nfet_06v0 ad=79.8f pd=0.8u as=0.2424p ps=1.635u w=0.38u l=0.6u
X6413 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I VGND.t1850 VGND.t1849 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6414 VPWR.t3053 a_4156_14136# a_4068_14180# VPWR.t3052 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6415 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN VPWR.t5783 VPWR.t5782 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6416 VPWR.t6934 a_42392_22825.t38 _452_.CLK.t24 VPWR.t6933 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6417 a_32240_31048# _363_.Z.t7 _370_.B VPWR.t45 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X6418 _417_.Z a_48776_20204# VGND.t3456 VGND.t3455 nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X6419 VGND.t5278 a_40464_27165# a_40416_27209# VGND.t5277 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X6420 a_59332_29816# _255_.I VPWR.t3834 VPWR.t3833 pfet_06v0 ad=0.1391p pd=1.055u as=0.4268p ps=2.175u w=0.535u l=0.5u
X6421 VPWR.t1778 a_28928_29123# a_28900_29535# VPWR.t1777 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X6422 VGND.t5216 _417_.Z a_49988_21236# VGND.t5215 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6423 a_17036_24679# a_16948_24776# VGND.t6083 VGND.t402 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6424 VPWR.t4161 a_4156_11000# a_4068_11044# VPWR.t2943 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6425 VPWR.t7024 _251_.A1.t33 a_56404_27208# VPWR.t7023 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6426 VPWR.t1338 a_17803_26841# a_18096_27165# VPWR.t1337 pfet_06v0 ad=0.38575p pd=1.92u as=0.2457p ps=1.465u w=0.945u l=0.5u
X6427 a_36008_20569# a_34160_20523# a_35723_20569# VPWR.t2900 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X6428 VPWR.t6082 a_61297_30300# _246_.B2 VPWR.t6081 pfet_06v0 ad=0.38705p pd=2.08u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6429 VPWR.t3044 a_27452_21543# a_27364_21640# VPWR.t3043 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6430 VGND.t6634 a_49152_30301.t6 a_50524_30345# VGND.t137 nfet_06v0 ad=0.1584p pd=1.6u as=43.2f ps=0.6u w=0.36u l=0.6u
X6431 uo_out[3].t4 a_41160_29083# VGND.t4027 VGND.t4026 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X6432 a_17036_21543# a_16948_21640# VGND.t2882 VGND.t2025 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6433 _346_.ZN _346_.B VPWR.t412 VPWR.t411 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X6434 VPWR.t4619 a_57692_1592# a_57604_1636# VPWR.t4618 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6435 a_2812_7864# a_2724_7908# VGND.t6084 VGND.t4074 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6436 _296_.ZN _350_.A1.t12 VGND.t6340 VGND.t102 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X6437 a_40452_18180# _451_.Q.t11 a_40244_18180# VGND.t6157 nfet_06v0 ad=60.8f pd=0.7u as=0.1672p ps=1.64u w=0.38u l=0.6u
X6438 a_42236_27815# a_42148_27912# VGND.t3272 VGND.t3271 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6439 VPWR.t6356 a_45148_1159# a_45060_1256# VPWR.t4931 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6440 _438_.ZN _304_.B a_39873_21236# VGND.t4524 nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X6441 a_38428_1159# a_38340_1256# VGND.t3180 VGND.t3179 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6442 a_3260_24679# a_3172_24776# VGND.t6087 VGND.t408 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6443 VPWR.t7133 a_17148_29816# a_17060_29860# VPWR.t3074 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6444 VPWR.t5873 a_14004_31048# a_14004_31048# VPWR.t5872 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6445 a_2812_4728# a_2724_4772# VGND.t2889 VGND.t762 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6446 a_60793_29860# _246_.B2 VPWR.t5209 VPWR.t5208 pfet_06v0 ad=0.1469p pd=1.085u as=0.38705p ps=2.08u w=0.565u l=0.5u
X6447 a_3260_21543# a_3172_21640# VGND.t3669 VGND.t3668 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6448 VPWR.t1345 a_64972_16839# a_64884_16936# VPWR.t1344 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6449 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I VPWR.t6314 VPWR.t6313 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6450 VGND.t5412 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN VGND.t5411 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6451 a_40656_23588# _300_.ZN a_40452_23588# VPWR.t5713 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6452 a_45904_30180# a_45416_29885# a_46336_30345# VGND.t137 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X6453 a_35292_30951# a_35204_31048# VGND.t1358 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6454 _393_.A1 _386_.ZN a_47525_29480# VPWR.t1881 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X6455 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN VPWR.t4865 VPWR.t4864 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6456 a_38548_21327# _301_.A1 a_38340_21327# VGND.t3200 nfet_06v0 ad=58.39999f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X6457 a_50384_19204# a_49936_19325.t4 a_50796_19001# VPWR.t120 pfet_06v0 ad=0.1872p pd=1.4u as=43.2f ps=0.6u w=0.36u l=0.5u
X6458 a_3260_1159# a_3172_1256# VGND.t2174 VGND.t2173 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6459 a_32156_19975# a_32068_20072# VGND.t6088 VGND.t5180 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6460 _412_.B2 a_50120_26476# VGND.t2354 VGND.t2353 nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X6461 VPWR.t5360 a_58588_11000# a_58500_11044# VPWR.t5359 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6462 VPWR.t1351 a_42572_16839# a_42484_16936# VPWR.t1350 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6463 a_20379_29977# a_18404_30344.t7 a_19744_30301# VPWR.t140 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X6464 a_52064_19715.t0 _474_.CLK.t53 VPWR.t6763 VPWR.t6762 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X6465 _407_.A1 _397_.A2.t19 VPWR.t6506 VPWR.t6505 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6466 a_46268_14136# a_46180_14180# VGND.t2336 VGND.t2335 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6467 VPWR.t152 _294_.ZN.t9 a_34260_29860# VPWR.t151 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6468 a_41440_28363# a_41028_28776.t6 VGND.t6779 VGND.t6778 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X6469 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN _248_.B1 VPWR.t1213 VPWR.t1212 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6470 VPWR.t2540 hold2.I _284_.ZN.t5 VPWR.t2539 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6471 VPWR.t2823 a_2812_27815# a_2724_27912# VPWR.t2822 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6472 a_46268_11000# a_46180_11044# VGND.t2340 VGND.t2339 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6473 a_67548_2727# a_67460_2824# VGND.t6090 VGND.t6089 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6474 a_20732_1592# a_20644_1636# VGND.t6007 VGND.t6006 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6475 VPWR.t757 a_62060_13703# a_61972_13800# VPWR.t756 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6476 a_42252_20936# _304_.A1.t12 _304_.ZN.t6 VGND.t6320 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6477 VPWR.t2670 a_1916_23544# a_1828_23588# VPWR.t2669 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6478 _284_.ZN.t3 _284_.A2.t7 a_42168_25640.t3 VGND.t29 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6479 a_4828_30951# a_4740_31048# VGND.t3527 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6480 a_44700_1592# a_44612_1636# VGND.t3264 VGND.t923 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6481 a_46940_17272# a_46852_17316# VGND.t5846 VGND.t5845 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6482 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I VGND.t1682 VGND.t1681 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6483 a_17596_29816# a_17508_29860# VGND.t6091 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6484 VPWR.t2913 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I VPWR.t2273 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6485 a_67548_15704# a_67460_15748# VGND.t5678 VGND.t5677 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6486 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN VGND.t5744 VGND.t5743 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6487 a_26220_23544# a_26132_23588# VGND.t2955 VGND.t2954 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6488 VPWR.t1281 a_52652_18407# a_52564_18504# VPWR.t1280 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6489 VPWR.t2848 a_1468_18840# a_1380_18884# VPWR.t1393 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6490 a_46772_29977# _393_.ZN a_45904_30180# VPWR.t3157 pfet_06v0 ad=54f pd=0.66u as=0.1872p ps=1.4u w=0.36u l=0.5u
X6491 a_35740_17272# a_35652_17316# VGND.t1417 VGND.t1416 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6492 a_28679_24776# _355_.C.t17 VPWR.t6679 VPWR.t6678 pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X6493 _324_.B.t11 _304_.B a_44028_22020# VPWR.t4680 pfet_06v0 ad=0.2847p pd=1.615u as=0.4599p ps=1.935u w=1.095u l=0.5u
X6494 VPWR.t1242 a_1468_15704# a_1380_15748# VPWR.t1241 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6495 a_59260_23111# a_59172_23208# VGND.t824 VGND.t823 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6496 a_34308_26344# _460_.Q _359_.ZN VPWR.t3476 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X6497 a_60380_12568# a_60292_12612# VGND.t2403 VGND.t2402 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6498 a_28820_24072# _336_.A1 VPWR.t4206 VPWR.t4205 pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X6499 a_46716_12568# a_46628_12612# VGND.t5471 VGND.t341 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6500 a_24092_24679# a_24004_24776# VGND.t6093 VGND.t6092 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6501 VPWR.t6160 a_49404_14136# a_49316_14180# VPWR.t6159 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6502 VPWR.t6275 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN VPWR.t6274 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X6503 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I VPWR.t4434 VPWR.t4433 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6504 VPWR.t2324 a_31168_24419# a_31140_24831# VPWR.t2323 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X6505 _474_.CLK.t27 a_48272_25156.t41 VGND.t6288 VGND.t6287 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X6506 a_60380_1159# a_60292_1256# VGND.t4926 VGND.t4925 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6507 a_40316_23233# _441_.A2 a_40004_23233# VPWR.t4309 pfet_06v0 ad=0.2847p pd=1.615u as=0.58035p ps=2.155u w=1.095u l=0.5u
X6508 VPWR.t3475 _460_.Q _335_.ZN.t9 VPWR.t3474 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X6509 a_35660_27508# a_35008_27533# VGND.t1986 VGND.t1985 nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X6510 a_24092_21543# a_24004_21640# VGND.t4268 VGND.t4267 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6511 VPWR.t1410 a_49404_11000# a_49316_11044# VPWR.t1409 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6512 a_25867_26841# a_24304_26795# a_25232_27165# VGND nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6513 a_58539_30644# a_58063_30644# VGND.t3084 VGND.t45 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6514 a_14684_29383# a_14596_29480# VGND.t4270 VGND.t4269 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6515 _331_.ZN _452_.Q.t19 VGND.t6645 VGND.t6644 nfet_06v0 ad=0.2569p pd=1.56u as=0.2244p ps=1.9u w=0.51u l=0.6u
X6516 _407_.ZN _397_.A4 VPWR.t1325 VPWR.t1324 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X6517 _330_.A2 _451_.Q.t12 a_38852_18884# VPWR.t5565 pfet_06v0 ad=0.31207p pd=1.665u as=0.55297p ps=2.105u w=1.095u l=0.5u
X6518 a_49180_15271# a_49092_15368# VGND.t1209 VGND.t1208 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6519 a_52228_19368# _424_.B1.t13 VGND.t6337 VGND.t6336 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6520 VPWR.t4074 a_31484_21543# a_31396_21640# VPWR.t4073 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6521 a_43776_18191# a_42896_18504# a_43452_18191# VGND.t5732 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X6522 VPWR.t2110 a_1020_13703# a_932_13800# VPWR.t2109 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6523 a_47172_23588# _397_.A1.t13 a_46984_23588# VPWR.t19 pfet_06v0 ad=0.196p pd=1.26u as=0.2464p ps=2u w=0.56u l=0.5u
X6524 VPWR.t366 a_2812_18407# a_2724_18504# VPWR.t365 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6525 a_39772_19975# a_39684_20072# VGND.t6165 VGND.t6164 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6526 VGND.t4152 _388_.B _393_.A1 VGND.t4151 nfet_06v0 ad=0.1209p pd=0.985u as=0.21175p ps=1.41u w=0.465u l=0.6u
X6527 VPWR.t2838 _407_.ZN _408_.ZN VPWR.t2837 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X6528 VPWR.t3999 a_10876_29383# a_10788_29480# VPWR.t3998 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6529 VPWR.t6355 a_2812_7864# a_2724_7908# VPWR.t5345 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6530 VPWR.t3337 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t3336 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6531 VPWR.t6569 a_48272_25156.t42 _474_.CLK.t28 VPWR.t6568 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6532 clkbuf_1_0__f_clk.I.t20 a_44296_24393.t37 VGND.t289 VGND.t288 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X6533 VPWR.t449 a_25772_23544# a_25684_23588# VPWR.t448 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6534 VPWR.t6664 _452_.CLK.t55 a_35204_24455.t0 VPWR.t6663 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X6535 VGND.t6246 _284_.ZN.t35 uo_out[0].t9 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X6536 a_35492_20072# _330_.A1.t22 _319_.ZN VPWR.t219 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6537 _433_.ZN _226_.ZN VGND.t2261 VGND.t2260 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6538 a_32628_26725# _460_.Q _362_.ZN VPWR.t3473 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X6539 VPWR.t5177 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN VPWR.t5176 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6540 VGND.t116 _411_.A2.t15 _419_.A4 VGND.t115 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X6541 _480_.Q a_43296_28733# VPWR.t6304 VPWR.t6303 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6542 VGND.t2745 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN VGND.t1847 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6543 a_53996_26680# a_53908_26724# VGND.t3930 VGND.t3929 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6544 a_33520_25597# a_33148_25641# VPWR.t6154 VPWR.t6153 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X6545 a_67436_16839# a_67348_16936# VGND.t6167 VGND.t6166 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6546 VPWR.t3284 a_52360_26355# a_53716_26399# VPWR.t3283 pfet_06v0 ad=0.4554p pd=3.25u as=54f ps=0.66u w=0.36u l=0.5u
X6547 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I VPWR.t5721 VPWR.t5720 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6548 a_13340_2727# a_13252_2824# VGND.t6168 VGND.t513 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6549 VPWR.t2292 a_6723_30644# uio_oe[7].t0 VPWR.t2291 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6550 VPWR.t2800 a_8636_29383# a_8548_29480# VPWR.t2799 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6551 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN VPWR.t5113 VPWR.t5112 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6552 VPWR.t372 a_28012_24679# a_27924_24776# VPWR.t371 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6553 a_16700_29383# a_16612_29480# VGND.t2736 VGND.t2735 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6554 VPWR.t374 a_3260_7431# a_3172_7528# VPWR.t373 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6555 VPWR.t7126 a_65308_19975# a_65220_20072# VPWR.t7125 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6556 a_2812_29816# a_2724_29860# VGND.t6169 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6557 VGND.t5779 _390_.ZN a_48859_29076# VGND.t5778 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6558 VPWR.t380 a_32380_2727# a_32292_2824# VPWR.t379 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6559 a_17148_1592# a_17060_1636# VGND.t5375 VGND.t1136 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6560 a_63852_23544# a_63764_23588# VGND.t3270 VGND.t3269 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6561 VPWR.t844 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN VPWR.t843 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6562 VPWR.t550 a_12444_1592# a_12356_1636# VPWR.t549 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6563 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I VPWR.t3585 VPWR.t3584 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6564 VPWR.t4447 a_64188_12568# a_64100_12612# VPWR.t4446 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6565 VGND.t2690 vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I VGND.t2689 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6566 a_20396_26680# a_20308_26724# VGND.t2655 VGND.t2654 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6567 a_51050_29480# _416_.A1.t14 _275_.ZN VPWR.t205 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6568 VPWR.t1812 a_36412_1592# a_36324_1636# VPWR.t1811 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6569 VPWR.t1699 a_21628_28248# a_21540_28292# VPWR.t1698 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6570 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I VGND.t1502 VGND.t1501 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6571 VPWR.t3211 a_22300_21543# a_22212_21640# VPWR.t3210 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6572 a_2364_25112# a_2276_25156# VGND.t5476 VGND.t5330 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6573 a_44270_21790# a_43814_21236# a_44038_21236# VPWR.t3829 pfet_06v0 ad=61.19999f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X6574 a_52848_25987# a_52360_26355# a_53280_26031# VGND.t3134 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X6575 VGND.t4516 a_54432_31128# _304_.B VGND.t4514 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X6576 VPWR.t1227 a_45820_10567# a_45732_10664# VPWR.t1226 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6577 VPWR.t1550 a_52428_13703# a_52340_13800# VPWR.t1549 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6578 a_50972_17272# a_50884_17316# VGND.t1437 VGND.t1436 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6579 a_2364_21976# a_2276_22020# VGND.t4954 VGND.t2977 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6580 VPWR.t6136 a_67100_4295# a_67012_4392# VPWR.t4054 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6581 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN VGND.t4920 VGND.t4919 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6582 VPWR.t7049 ui_in[4].t1 a_58063_30644# VPWR.t7048 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X6583 a_20379_29977# a_18816_29931# a_19744_30301# VGND.t137 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6584 VPWR.t5671 _375_.Z _378_.I VPWR.t5670 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6585 a_52434_22504# _475_.Q a_52240_22504# VGND.t4855 nfet_06v0 ad=0.1517p pd=1.19u as=0.1517p ps=1.19u w=0.82u l=0.6u
X6586 a_28256_25597# a_27884_25641# VGND.t2828 VGND.t2827 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X6587 VPWR.t6936 a_42392_22825.t39 _452_.CLK.t25 VPWR.t6935 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6588 VPWR.t2813 a_67100_1159# a_67012_1256# VPWR.t2812 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6589 a_61948_12568# a_61860_12612# VGND.t3745 VGND.t3744 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6590 VPWR.t5769 a_64636_14136# a_64548_14180# VPWR.t5768 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6591 a_42168_22504# _304_.B _324_.B.t7 VGND.t4523 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6592 a_17484_24679# a_17396_24776# VGND.t6170 VGND.t523 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6593 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I VPWR.t2868 VPWR.t2867 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6594 _369_.ZN _371_.A3 VGND.t953 VGND.t952 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X6595 VPWR.t6843 clk.t12 a_44296_24393.t12 VPWR.t6842 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X6596 a_50748_12568# a_50660_12612# VGND.t5957 VGND.t5956 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6597 VPWR.t2450 a_64636_11000# a_64548_11044# VPWR.t2449 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6598 a_17484_21543# a_17396_21640# VGND.t5840 VGND.t3540 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6599 a_65756_7431# a_65668_7528# VGND.t6171 VGND.t4034 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6600 a_27228_26247# a_27140_26344# VGND.t681 VGND.t680 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6601 VPWR.t3322 a_67741_30600# a_67861_31220# VPWR.t3321 pfet_06v0 ad=0.1116p pd=0.98u as=61.19999f ps=0.7u w=0.36u l=0.5u
X6602 VGND.t2726 vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I VGND.t2725 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6603 VPWR.t1435 a_9532_2727# a_9444_2824# VPWR.t1434 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6604 a_2812_23544# a_2724_23588# VGND.t3408 VGND.t1398 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6605 VPWR.t6666 _452_.CLK.t56 a_32740_22504.t0 VPWR.t6665 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X6606 a_42684_27815# a_42596_27912# VGND.t5866 VGND.t5865 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6607 a_31080_29977# a_29232_29931# a_30795_29977# VPWR.t1030 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X6608 VPWR.t3513 a_65308_5863# a_65220_5960# VPWR.t3102 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6609 a_8188_29816# a_8100_29860# VGND.t6172 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6610 VPWR.t6362 a_17596_29816# a_17508_29860# VPWR.t6361 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6611 a_67996_21976# a_67908_22020# VGND.t5263 VGND.t5262 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6612 VPWR.t1820 a_8860_1592# a_8772_1636# VPWR.t1819 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6613 VPWR.t4455 a_55004_12568# a_54916_12612# VPWR.t4454 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6614 VGND.t1056 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I VGND.t1055 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6615 VPWR.t6668 _452_.CLK.t57 a_45508_20936.t0 VPWR.t6667 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X6616 VPWR.t2088 a_58588_9432# a_58500_9476# VPWR.t2087 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6617 VPWR.t538 vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN VPWR.t537 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6618 a_44752_18147# a_44459_18559# VGND.t3047 VGND.t3046 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X6619 _351_.ZN _351_.A2 VGND.t3105 VGND.t3104 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6620 VPWR.t4928 a_19388_1159# a_19300_1256# VPWR.t2042 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6621 a_49292_10567# a_49204_10664# VGND.t6174 VGND.t6173 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6622 VPWR.t1096 a_40668_1592# a_40580_1636# VPWR.t1095 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6623 VGND.t4683 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t4682 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6624 VPWR.t2082 a_18716_30951# a_18628_31048# VPWR.t2081 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6625 a_23644_29816# a_23556_29860# VGND.t6175 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6626 a_31708_18840# a_31620_18884# VGND.t3361 VGND.t77 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6627 a_2364_15704# a_2276_15748# VGND.t4082 VGND.t3511 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6628 a_35292_2727# a_35204_2824# VGND.t6177 VGND.t6176 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6629 VPWR.t1098 a_64636_1592# a_64548_1636# VPWR.t1097 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6630 a_50188_12135# a_50100_12232# VGND.t3012 VGND.t3011 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6631 a_46268_10567# a_46180_10664# VGND.t6178 VGND.t3897 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6632 a_12444_29816# a_12356_29860# VGND.t6179 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6633 VGND.t6672 _352_.A2.t27 a_29163_24394# VGND.t6671 nfet_06v0 ad=0.3124p pd=2.3u as=85.2f ps=0.95u w=0.71u l=0.6u
X6634 VPWR.t1440 a_59036_2727# a_58948_2824# VPWR.t1439 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6635 VGND.t3786 _427_.B2 a_52452_21236# VGND.t3785 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6636 VPWR.t1442 a_54444_24679# a_54356_24776# VPWR.t1441 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6637 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN VPWR.t3153 VPWR.t3152 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6638 VGND.t3175 a_67741_30600# a_67861_30644# VGND.t45 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X6639 a_5276_29383# a_5188_29480# VGND.t5907 VGND.t5906 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6640 VPWR.t5551 a_5052_4728# a_4964_4772# VPWR.t5550 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6641 a_46580_23588# _402_.A1.t22 _402_.B VPWR.t267 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X6642 a_30140_21543# a_30052_21640# VGND.t5950 VGND.t5949 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6643 a_45148_1159# a_45060_1256# VGND.t6086 VGND.t6085 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6644 VPWR.t5080 a_5052_1592# a_4964_1636# VPWR.t5079 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6645 _450_.D _330_.A1.t23 VGND.t224 VGND.t223 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6646 VPWR.t6347 a_39324_19975# a_39236_20072# VPWR.t6346 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6647 VPWR.t654 a_1916_30951# a_1828_31048# VPWR.t653 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6648 VPWR.t3957 a_1468_29383# a_1380_29480# VPWR.t2015 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6649 VPWR.t6120 a_65084_1159# a_64996_1256# VPWR.t5361 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6650 a_50636_13703# a_50548_13800# VGND.t4184 VGND.t4183 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6651 VPWR.t5353 a_60828_26680# a_60740_26724# VPWR.t5352 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6652 a_66204_9432# a_66116_9476# VGND.t5739 VGND.t5738 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6653 a_67996_15704# a_67908_15748# VGND.t6052 VGND.t6051 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6654 a_23308_20408# a_23220_20452# VGND.t5921 VGND.t5920 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6655 _399_.ZN _399_.A1 a_49013_22805# VGND.t4077 nfet_06v0 ad=0.2015p pd=1.295u as=92.99999f ps=1.015u w=0.775u l=0.6u
X6656 a_63404_12135# a_63316_12232# VGND.t4272 VGND.t4271 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6657 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I VGND.t5420 VGND.t5419 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6658 VPWR.t658 a_1468_26247# a_1380_26344# VPWR.t657 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6659 a_66204_6296# a_66116_6340# VGND.t5925 VGND.t5924 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6660 a_18940_1592# a_18852_1636# VGND.t3164 VGND.t3163 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6661 a_47776_20893# a_47483_20569# VPWR.t3082 VPWR.t3081 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X6662 VGND.t39 _363_.Z.t8 _461_.D VGND.t38 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6663 a_38816_27555# a_38523_27967# VPWR.t1012 VPWR.t1011 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X6664 a_47732_22504# _416_.A3 VGND.t4316 VGND.t4315 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6665 VGND.t6322 _304_.A1.t13 _430_.ZN VGND.t6321 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X6666 a_62172_18407# a_62084_18504# VGND.t6180 VGND.t964 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6667 VPWR.t426 a_1468_23111# a_1380_23208# VPWR.t425 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6668 VPWR.t704 a_31820_23544# a_31732_23588# VPWR.t703 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6669 VGND.t1033 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I VGND.t1032 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6670 a_31088_30301# a_30795_29977# VPWR.t2284 VPWR.t2283 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X6671 a_48508_18407# a_48420_18504# VGND.t6182 VGND.t6181 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6672 a_30724_26020# _336_.Z VPWR.t4559 VPWR.t4558 pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X6673 a_42908_30951# a_42820_31048# VGND.t5304 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6674 VGND.t5511 _300_.ZN _432_.ZN VGND.t5510 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6675 VPWR.t5725 a_49852_14136# a_49764_14180# VPWR.t5724 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6676 VPWR.t710 a_20620_23544# a_20532_23588# VPWR.t709 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6677 VGND.t739 vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I VGND.t738 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6678 a_34396_15704# a_34308_15748# VGND.t4040 VGND.t4039 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6679 VPWR.t1910 _247_.ZN a_59796_29480# VPWR.t1909 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6680 a_59932_11000# a_59844_11044# VGND.t3020 VGND.t3019 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6681 a_34052_22137# a_32740_22504.t7 a_33708_22505# VPWR.t101 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X6682 VPWR.t6439 a_2812_29816# a_2724_29860# VPWR.t1607 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6683 VPWR.t1287 a_49852_11000# a_49764_11044# VPWR.t1286 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6684 VGND.t5644 _436_.B _436_.ZN VGND.t5643 nfet_06v0 ad=0.1209p pd=0.985u as=0.21175p ps=1.41u w=0.465u l=0.6u
X6685 VPWR.t927 a_4156_16839# a_4068_16936# VPWR.t926 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6686 VPWR.t3987 a_2812_26680# a_2724_26724# VPWR.t3028 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6687 vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN VPWR.t6253 VPWR.t6252 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6688 VPWR.t931 a_30812_16839# a_30724_16936# VPWR.t930 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6689 VPWR.t1108 a_65072_29860# _324_.C.t1 VPWR.t1107 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6690 a_67996_6296# a_67908_6340# VGND.t3371 VGND.t3370 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6691 VGND.t1014 _383_.A2 _383_.ZN VGND.t1013 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6692 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I VPWR.t4478 VPWR.t4477 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6693 vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I VPWR.t1638 VPWR.t1637 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6694 VGND.t4723 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6695 a_15132_1592# a_15044_1636# VGND.t3298 VGND.t3297 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6696 a_39100_1592# a_39012_1636# VGND.t5361 VGND.t3161 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6697 VGND.t1769 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t1768 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6698 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN VPWR.t3173 VPWR.t3172 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6699 a_1468_7864# a_1380_7908# VGND.t6183 VGND.t2439 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6700 a_67884_16839# a_67796_16936# VGND.t6185 VGND.t6184 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6701 _399_.A2 _397_.Z a_48308_23588# VPWR.t895 pfet_06v0 ad=0.2964p pd=1.66u as=0.5016p ps=3.16u w=1.14u l=0.5u
X6702 a_1468_4728# a_1380_4772# VGND.t2773 VGND.t2772 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6703 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I VGND.t2252 VGND.t2251 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6704 a_16588_25112# a_16500_25156# VGND.t2550 VGND.t2491 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6705 a_60059_28776# _229_.I.t12 _252_.B VGND.t6568 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6706 VPWR.t2629 a_11548_30951# a_11460_31048# VPWR.t2628 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6707 VPWR.t2454 a_53884_20408# a_53796_20452# VPWR.t2453 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6708 a_28556_29167# _373_.ZN a_28432_29535# VPWR.t1423 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X6709 _474_.Q a_48888_19243# VGND.t2760 VGND.t2759 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6710 VPWR.t5366 a_37196_23544# a_37108_23588# VPWR.t5365 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6711 uo_out[7].t5 a_40038_28720# VGND.t2984 VGND.t2983 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6712 VPWR.t917 a_12892_2727# a_12804_2824# VPWR.t916 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6713 a_34715_22137# a_33152_22091# a_34080_22461# VGND.t1394 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6714 a_41922_31073# _304_.B _495_.I VPWR.t4679 pfet_06v0 ad=0.55297p pd=2.105u as=0.31207p ps=1.665u w=1.095u l=0.5u
X6715 a_16588_21976# a_16500_22020# VGND.t4597 VGND.t1561 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6716 a_57220_29861# _268_.A2.t7 a_56596_29861# VPWR.t7064 pfet_06v0 ad=0.37665p pd=1.835u as=0.3402p ps=1.775u w=1.215u l=0.5u
X6717 a_48964_20204# _417_.A2.t12 a_48776_20204# VPWR.t136 pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X6718 VGND.t2167 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I VGND.t2082 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6719 VGND.t1101 _340_.ZN _342_.ZN VGND.t1100 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6720 a_20508_24679# a_20420_24776# VGND.t6187 VGND.t6186 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6721 VPWR.t1384 a_25436_24679# a_25348_24776# VPWR.t1383 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6722 VPWR.t6443 a_8188_29816# a_8100_29860# VPWR.t6442 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6723 _223_.I a_31088_30301# VPWR.t7137 VPWR.t7136 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6724 VPWR.t4256 a_49740_29383# a_49652_29480# VPWR.t4255 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6725 a_38768_27599# a_36548_27591.t6 a_38523_27967# VGND.t6326 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6726 a_59820_12135# a_59732_12232# VGND.t5889 VGND.t5888 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6727 VPWR.t4584 a_1020_12568# a_932_12612# VPWR.t4583 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6728 VPWR.t6487 _459_.CLK.t38 a_31508_29159.t0 VPWR.t6486 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X6729 VPWR.t4407 a_62844_9432# a_62756_9476# VPWR.t4406 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6730 a_20508_21543# a_20420_21640# VGND.t3775 VGND.t3774 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6731 VPWR.t4408 a_2812_17272# a_2724_17316# VPWR.t3166 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6732 VPWR.t428 a_52876_13703# a_52788_13800# VPWR.t427 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6733 VPWR.t6447 a_23644_29816# a_23556_29860# VPWR.t6446 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6734 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN VPWR.t4430 VPWR.t4429 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6735 VPWR.t630 a_47612_1159# a_47524_1256# VPWR.t629 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6736 a_58028_13703# a_57940_13800# VGND.t5772 VGND.t5771 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6737 VPWR.t6359 a_32156_19975# a_32068_20072# VPWR.t6358 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6738 a_37392_27967# a_36960_27912# VPWR.t5486 VPWR.t5485 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X6739 VPWR.t6451 a_12444_29816# a_12356_29860# VPWR.t1916 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6740 VPWR.t3900 a_34304_24029# a_34276_23705# VPWR.t3899 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X6741 VPWR.t1307 a_5388_10567# a_5300_10664# VPWR.t1306 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6742 a_43356_1592# a_43268_1636# VGND.t1972 VGND.t1971 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6743 VPWR.t5526 vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN VPWR.t5525 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6744 a_42778_21812# a_42154_21236# a_42610_21812# VPWR.t2504 pfet_06v0 ad=0.3852p pd=2.86u as=61.19999f ps=0.7u w=0.36u l=0.5u
X6745 a_41664_22020# _327_.A2 a_41460_22020# VPWR.t3397 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6746 a_29804_21976# a_29716_22020# VGND.t4492 VGND.t4491 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6747 VPWR.t5751 a_19724_21976# a_19636_22020# VPWR.t5750 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6748 a_67324_1592# a_67236_1636# VGND.t2999 VGND.t2998 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6749 a_58700_16839# a_58612_16936# VGND.t6749 VGND.t6748 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6750 a_38852_25156# _311_.A2.t11 a_38628_25156# VPWR.t6381 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6751 VPWR.t648 a_3260_9432# a_3172_9476# VPWR.t647 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6752 VPWR.t769 a_62620_1592# a_62532_1636# VPWR.t768 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6753 VPWR.t2418 a_16140_26247# a_16052_26344# VPWR.t2417 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6754 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I VPWR.t2276 VPWR.t2275 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6755 a_57468_1159# a_57380_1256# VGND.t1303 VGND.t1302 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6756 VPWR.t126 _281_.ZN.t9 a_46794_25156# VPWR.t125 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X6757 VPWR.t2420 a_24316_26247# a_24228_26344# VPWR.t2419 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6758 a_27676_26247# a_27588_26344# VGND.t4782 VGND.t4781 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6759 a_59260_26680# a_59172_26724# VGND.t5285 VGND.t5284 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6760 VPWR.t1309 a_57020_2727# a_56932_2824# VPWR.t1308 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6761 VPWR.t1311 a_46268_18407# a_46180_18504# VPWR.t1310 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6762 VPWR.t571 a_28012_23544# a_27924_23588# VPWR.t570 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6763 VPWR.t2421 a_47836_15271# a_47748_15368# VPWR.t1509 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6764 VGND.t5756 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I VGND.t5755 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6765 a_47500_16839# a_47412_16936# VGND.t6751 VGND.t6750 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6766 a_52756_29076# _274_.A2 VGND.t5674 VGND.t5673 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6767 VPWR.t2422 a_16140_23111# a_16052_23208# VPWR.t731 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6768 VPWR.t575 a_32380_1592# a_32292_1636# VPWR.t574 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6769 a_57500_30344# _272_.B1 _274_.A2 VGND.t325 nfet_06v0 ad=85.2f pd=0.95u as=0.21175p ps=1.41u w=0.71u l=0.6u
X6770 VPWR.t4590 a_55452_12568# a_55364_12612# VPWR.t4589 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6771 a_29575_28293# _370_.B a_29351_28293# VPWR.t5730 pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X6772 vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN VGND.t5303 VGND.t5302 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6773 a_31088_30301# a_30795_29977# VGND.t2177 VGND.t2052 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X6774 clkbuf_1_0__f_clk.I.t3 a_44296_24393.t38 VPWR.t292 VPWR.t291 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6775 VPWR.t4449 a_45088_29123# a_45080_29535# VPWR.t4448 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X6776 VPWR.t1138 a_39548_2727# a_39460_2824# VPWR.t1137 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6777 a_31040_30345# a_28820_30344.t5 a_30795_29977# VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6778 a_12892_29816# a_12804_29860# VGND.t6752 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6779 VPWR.t5302 a_34844_17272# a_34756_17316# VPWR.t5301 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6780 VPWR.t1144 a_54892_24679# a_54804_24776# VPWR.t1143 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6781 VPWR.t2613 a_51868_1159# a_51780_1256# VPWR.t2612 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6782 VPWR.t6455 a_1468_7864# a_1380_7908# VPWR.t6114 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6783 a_64412_17272# a_64324_17316# VGND.t2926 VGND.t1643 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6784 VPWR.t3345 _301_.A1 _434_.ZN VPWR.t3344 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X6785 VPWR.t3226 a_55900_14136# a_55812_14180# VPWR.t3225 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6786 VGND.t4005 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I VGND.t4004 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6787 VPWR.t5564 _327_.Z a_40244_18180# VPWR.t5563 pfet_06v0 ad=0.4268p pd=2.175u as=0.1391p ps=1.055u w=0.535u l=0.5u
X6788 a_40444_15704# a_40356_15748# VGND.t3578 VGND.t3577 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6789 a_53212_17272# a_53124_17316# VGND.t2068 VGND.t2067 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6790 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t5464 VGND.t5463 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6791 VPWR.t3195 a_55900_11000# a_55812_11044# VPWR.t3194 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6792 a_42236_2727# a_42148_2824# VGND.t310 VGND.t309 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6793 _252_.ZN _231_.ZN a_59397_26344# VPWR.t4365 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X6794 VPWR.t7072 a_45596_1159# a_45508_1256# VPWR.t5874 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6795 a_4156_12568# a_4068_12612# VGND.t2127 VGND.t2126 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6796 a_46716_9432# a_46628_9476# VGND.t2558 VGND.t2557 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6797 VPWR.t6434 a_39772_19975# a_39684_20072# VPWR.t5876 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6798 VGND.t6011 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN VGND.t6010 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6799 a_66204_2727# a_66116_2824# VGND.t822 VGND.t821 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6800 a_49316_23588# _279_.Z a_48308_23588# VPWR.t5586 pfet_06v0 ad=0.3534p pd=1.76u as=0.2964p ps=1.66u w=1.14u l=0.5u
X6801 VPWR.t3248 a_65308_4728# a_65220_4772# VPWR.t677 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6802 VPWR.t988 a_61276_2727# a_61188_2824# VPWR.t987 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6803 a_23756_20408# a_23668_20452# VGND.t5200 VGND.t5199 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6804 a_60276_26724# _252_.B _247_.B VPWR.t789 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6805 a_63852_12135# a_63764_12232# VGND.t3713 VGND.t3712 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6806 VPWR.t3723 a_4604_6296# a_4516_6340# VPWR.t3722 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6807 a_56124_27815# a_56036_27912# VGND.t3312 VGND.t3311 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6808 VPWR.t4375 a_4604_3160# a_4516_3204# VPWR.t4374 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6809 VPWR.t5029 a_61948_26247# a_61860_26344# VPWR.t5028 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6810 a_57120_31048# _474_.CLK.t54 VPWR.t6765 VPWR.t6764 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6811 _250_.B vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN a_63524_29098# VGND.t4722 nfet_06v0 ad=0.21175p pd=1.41u as=85.2f ps=0.95u w=0.71u l=0.6u
X6812 a_48956_18407# a_48868_18504# VGND.t2841 VGND.t2840 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6813 VPWR.t759 a_35068_1592# a_34980_1636# VPWR.t758 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6814 VPWR.t761 a_65644_23544# a_65556_23588# VPWR.t760 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6815 _404_.A1 _470_.Q VGND.t4064 VGND.t4063 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X6816 VGND.t2698 _407_.ZN a_51883_27508# VGND.t2697 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6817 a_5388_19975# a_5300_20072# VGND.t6756 VGND.t6755 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6818 VGND.t6213 _459_.CLK.t39 a_17060_28776.t1 VGND.t6212 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X6819 VPWR.t763 a_59036_1592# a_58948_1636# VPWR.t762 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6820 VPWR.t5986 a_21424_25987# a_21396_26399# VPWR.t5985 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X6821 VGND.t3190 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t3189 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6822 VGND.t5631 a_25936_25597# a_25888_25641# VGND.t5630 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X6823 VPWR.t554 a_54444_23544# a_54356_23588# VPWR.t553 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6824 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I VGND.t1073 VGND.t1072 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6825 VGND.t3129 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t3128 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6826 VPWR.t5804 a_52316_27815# a_52228_27912# VPWR.t5803 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6827 a_67996_2727# a_67908_2824# VGND.t5754 VGND.t5753 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6828 a_22636_25112# a_22548_25156# VGND.t2145 VGND.t2144 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6829 VPWR.t1677 a_22992_27555# a_22964_27967# VPWR.t1676 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X6830 a_62732_16839# a_62644_16936# VGND.t319 VGND.t318 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6831 VGND.t5013 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN VGND.t5012 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6832 a_58588_12568# a_58500_12612# VGND.t2105 VGND.t2104 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6833 a_22636_21976# a_22548_22020# VGND.t4425 VGND.t4424 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6834 a_33483_29535# a_31920_29480# a_32848_29123# VGND.t3138 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X6835 VPWR.t4313 _388_.B a_41922_31073# VPWR.t4312 pfet_06v0 ad=0.4818p pd=3.07u as=0.55297p ps=2.105u w=1.095u l=0.5u
X6836 a_44756_19001# _325_.ZN a_43888_19204# VPWR.t325 pfet_06v0 ad=54f pd=0.66u as=0.1872p ps=1.4u w=0.36u l=0.5u
X6837 a_26160_27165# a_25867_26841# VPWR.t3659 VPWR.t3658 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X6838 a_2812_15271# a_2724_15368# VGND.t2462 VGND.t2461 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6839 VPWR.t3824 a_1468_28248# a_1380_28292# VPWR.t3823 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6840 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN VPWR.t5073 VPWR.t5072 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6841 VPWR.t1979 a_45260_16839# a_45172_16936# VPWR.t1978 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6842 VGND.t4865 a_20672_30301# uio_out[5].t4 VGND.t71 nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X6843 VPWR.t5042 a_40668_15271# a_40580_15368# VPWR.t5041 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6844 VPWR.t6336 _288_.ZN.t10 a_36948_29860# VPWR.t6335 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6845 a_2812_12135# a_2724_12232# VGND.t2897 VGND.t2896 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6846 VPWR.t4418 a_1468_25112# a_1380_25156# VPWR.t4417 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6847 _287_.A1.t2 a_38472_30169# VPWR.t4963 VPWR.t4962 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6848 VPWR.t6594 _447_.Q.t17 _434_.ZN VPWR.t6593 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X6849 a_27228_26680# a_27140_26724# VGND.t5567 VGND.t5566 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6850 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN VGND.t3531 VGND.t3530 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6851 _436_.ZN _432_.ZN VGND.t5400 VGND.t5399 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X6852 VPWR.t6427 _451_.Q.t13 a_40244_18180# VPWR.t6426 pfet_06v0 ad=0.1391p pd=1.055u as=0.2354p ps=1.95u w=0.535u l=0.5u
X6853 _399_.A2 _279_.Z VGND.t5386 VGND.t5385 nfet_06v0 ad=0.1339p pd=1.035u as=0.23325p ps=1.48u w=0.515u l=0.6u
X6854 VPWR.t2112 a_4604_23544# a_4516_23588# VPWR.t2111 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6855 a_39264_18147# a_38971_18559# VPWR.t1797 VPWR.t1796 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X6856 VPWR.t1986 a_66540_18407# a_66452_18504# VPWR.t1985 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6857 a_28880_29167# a_28000_29480# a_28556_29167# VGND.t1838 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X6858 VPWR.t1988 a_3260_10567# a_3172_10664# VPWR.t1987 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6859 a_64188_2727# a_64100_2824# VGND.t5735 VGND.t980 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6860 a_36016_20893# a_35723_20569# VPWR.t4048 VPWR.t4047 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X6861 VGND.t5571 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I VGND.t5570 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6862 _252_.ZN _251_.A1.t34 a_59605_25962# VGND.t6705 nfet_06v0 ad=0.21175p pd=1.41u as=85.2f ps=0.95u w=0.71u l=0.6u
X6863 a_50412_18407# a_50324_18504# VGND.t4197 VGND.t4196 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6864 vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN VPWR.t2120 VPWR.t2119 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6865 a_3260_4295# a_3172_4392# VGND.t4014 VGND.t3294 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6866 VPWR.t1990 a_63516_18407# a_63428_18504# VPWR.t1989 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6867 VPWR.t1076 a_4156_18840# a_4068_18884# VPWR.t1075 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6868 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I VPWR.t2124 VPWR.t2123 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6869 _350_.A2.t0 _223_.ZN VPWR.t794 VPWR.t793 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X6870 VPWR.t1082 a_30812_18840# a_30724_18884# VPWR.t1081 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6871 VPWR.t1994 a_25884_24679# a_25796_24776# VPWR.t1993 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6872 VPWR.t5403 a_67772_21543# a_67684_21640# VPWR.t5402 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6873 a_20956_24679# a_20868_24776# VGND.t312 VGND.t311 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6874 a_27884_25641# _355_.ZN a_27716_25641# VGND.t2448 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X6875 VGND.t3838 _359_.ZN a_33188_25940# VGND.t3837 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X6876 VPWR.t2118 a_4156_15704# a_4068_15748# VPWR.t2117 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6877 VPWR.t5717 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I VPWR.t5716 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6878 VPWR.t1542 a_11100_1592# a_11012_1636# VPWR.t1541 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6879 VPWR.t1544 a_30812_15704# a_30724_15748# VPWR.t1543 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6880 VPWR.t5190 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I VPWR.t5189 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6881 VGND.t717 _427_.A2 a_52660_24072# VGND.t716 nfet_06v0 ad=0.23405p pd=1.555u as=58.39999f ps=0.685u w=0.365u l=0.6u
X6882 VPWR.t6489 _459_.CLK.t40 a_32180_25640.t0 VPWR.t6488 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X6883 a_49404_12568# a_49316_12612# VGND.t1761 VGND.t1760 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6884 _301_.A1 a_35008_22461# VGND.t5784 VGND.t5783 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6885 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I VGND.t1767 VGND.t1766 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6886 a_20956_21543# a_20868_21640# VGND.t2423 VGND.t2422 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6887 a_33724_23111# a_33636_23208# VGND.t2938 VGND.t2937 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6888 VGND.t1508 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t1507 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X6889 _452_.CLK.t26 a_42392_22825.t40 VGND.t6621 VGND.t6620 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X6890 VPWR.t4815 a_61500_12568# a_61412_12612# VPWR.t4814 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6891 hold2.I _260_.ZN a_42161_24776# VPWR.t3622 pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X6892 a_58476_13703# a_58388_13800# VGND.t3259 VGND.t3258 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6893 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t2446 VGND.t71 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X6894 VPWR.t826 a_43804_2727# a_43716_2824# VPWR.t825 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6895 a_7068_1159# a_6980_1256# VGND.t3373 VGND.t3372 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6896 a_56180_22137# _427_.ZN a_55312_22340# VPWR.t3784 pfet_06v0 ad=54f pd=0.66u as=0.1872p ps=1.4u w=0.36u l=0.5u
X6897 a_35188_22895# _304_.A1.t14 a_34980_22895# VGND.t6323 nfet_06v0 ad=58.39999f pd=0.685u as=0.1606p ps=1.61u w=0.365u l=0.6u
X6898 VPWR.t7071 a_12892_29816# a_12804_29860# VPWR.t1218 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6899 _365_.ZN a_35008_27533# VPWR.t2086 VPWR.t2085 pfet_06v0 ad=0.31207p pd=1.665u as=0.34437p ps=1.895u w=1.095u l=0.5u
X6900 a_23868_1592# a_23780_1636# VGND.t4126 VGND.t3228 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6901 _331_.ZN _451_.Q.t14 a_40416_18885# VPWR.t6428 pfet_06v0 ad=0.3159p pd=1.735u as=0.44955p ps=1.955u w=1.215u l=0.5u
X6902 a_23196_1159# a_23108_1256# VGND.t936 VGND.t935 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6903 VPWR.t4615 a_50300_12568# a_50212_12612# VPWR.t4614 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6904 VGND.t6215 _459_.CLK.t41 a_31508_29159.t1 VGND.t6214 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X6905 a_32308_29167# a_31508_29159.t7 VGND.t91 VGND.t90 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X6906 VPWR.t5621 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN VPWR.t5620 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6907 a_60156_27815# a_60068_27912# VGND.t344 VGND.t343 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6908 a_52924_20127# a_52408_19759# VPWR.t2740 VPWR.t2739 pfet_06v0 ad=43.2f pd=0.6u as=0.1044p ps=0.94u w=0.36u l=0.5u
X6909 a_26712_29977# a_24864_29931# a_26427_29977# VPWR.t4036 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X6910 VPWR.t830 a_65868_10567# a_65780_10664# VPWR.t829 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6911 a_39760_23588# _437_.A1.t12 a_39536_23588# VPWR.t5254 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6912 VPWR.t832 a_37532_2727# a_37444_2824# VPWR.t831 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6913 a_29788_30345# _370_.ZN a_29664_29977# VPWR.t1927 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X6914 a_17596_1592# a_17508_1636# VGND.t2494 VGND.t2493 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6915 VPWR.t1552 a_12892_1592# a_12804_1636# VPWR.t1551 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6916 clkbuf_1_0__f_clk.I.t19 a_44296_24393.t39 VGND.t291 VGND.t290 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X6917 VPWR.t808 a_54668_10567# a_54580_10664# VPWR.t807 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6918 VPWR.t1554 a_28460_23544# a_28372_23588# VPWR.t1553 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6919 a_61276_19975# a_61188_20072# VGND.t6758 VGND.t6757 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6920 a_37844_29860# _287_.A1.t32 uo_out[2].t2 VPWR.t6789 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X6921 VPWR.t1558 a_36860_1592# a_36772_1636# VPWR.t1557 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6922 a_47552_19715# a_47259_20127# VPWR.t2463 VPWR.t2462 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X6923 a_64412_7431# a_64324_7528# VGND.t3472 VGND.t3471 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6924 VPWR.t6295 a_24316_1159# a_24228_1256# VPWR.t6294 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6925 a_41392_27165# a_41099_26841# VPWR.t5463 VPWR.t5462 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X6926 VPWR.t1560 a_47388_15704# a_47300_15748# VPWR.t1559 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6927 VGND.t150 _294_.ZN.t10 uo_out[4].t8 VGND.t146 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X6928 VPWR.t2296 a_30924_20408# a_30836_20452# VPWR.t2295 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6929 VPWR.t4780 a_3708_21543# a_3620_21640# VPWR.t3089 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6930 clkbuf_1_0__f_clk.I.t2 a_44296_24393.t40 VPWR.t294 VPWR.t293 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X6931 a_25008_25597# a_24636_25641# VPWR.t4743 VPWR.t4742 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X6932 VPWR.t270 clkbuf_1_0__f_clk.I.t56 a_48272_25156.t1 VPWR.t269 pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X6933 a_64188_14136# a_64100_14180# VGND.t4148 VGND.t4147 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6934 VPWR.t1566 a_36188_15704# a_36100_15748# VPWR.t1565 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6935 VPWR.t445 a_57916_25112# a_57828_25156# VPWR.t444 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6936 VPWR.t447 a_57244_9432# a_57156_9476# VPWR.t446 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6937 a_5500_29816# a_5412_29860# VGND.t6759 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6938 VPWR.t7079 a_18044_1159# a_17956_1256# VPWR.t1186 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6939 _435_.A3 _451_.Q.t15 VPWR.t6430 VPWR.t6429 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X6940 _371_.A2 _337_.A3.t15 VPWR.t6413 VPWR.t6412 pfet_06v0 ad=0.2197p pd=1.365u as=0.4056p ps=1.805u w=0.845u l=0.5u
X6941 VPWR.t816 a_35628_16839# a_35540_16936# VPWR.t815 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6942 a_64188_11000# a_64100_11044# VGND.t4711 VGND.t4710 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6943 VPWR.t3903 a_45372_12135# a_45284_12232# VPWR.t3902 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6944 VGND.t6493 _287_.A1.t33 uo_out[6].t8 VGND.t6492 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X6945 VPWR.t2873 a_16140_28248# a_16052_28292# VPWR.t2872 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6946 a_64188_1159# a_64100_1256# VGND.t1275 VGND.t1274 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6947 VPWR.t1277 a_66316_13703# a_66228_13800# VPWR.t1276 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6948 a_55340_23544# a_55252_23588# VGND.t2407 VGND.t1329 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6949 a_44112_29167# a_43232_29480# a_43788_29167# VGND.t789 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X6950 VPWR.t607 vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN VPWR.t606 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6951 a_64860_17272# a_64772_17316# VGND.t1763 VGND.t1762 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6952 a_5052_25112# a_4964_25156# VGND.t4228 VGND.t4227 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6953 a_43296_28733# a_43003_28409# VPWR.t1652 VPWR.t1651 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X6954 VGND.t6128 _325_.A2.t11 a_43932_17800# VGND.t6127 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X6955 a_3260_19975# a_3172_20072# VGND.t6762 VGND.t5213 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6956 a_54192_22851# a_53744_22851.t7 a_54604_23263# VPWR.t28 pfet_06v0 ad=0.1872p pd=1.4u as=43.2f ps=0.6u w=0.36u l=0.5u
X6957 VPWR.t857 a_9980_2727# a_9892_2824# VPWR.t856 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6958 a_22748_2727# a_22660_2824# VGND.t1817 VGND.t1816 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6959 VPWR.t1279 a_55116_13703# a_55028_13800# VPWR.t1278 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6960 VPWR.t3616 a_16140_25112# a_16052_25156# VPWR.t3369 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6961 a_40892_15704# a_40804_15748# VGND.t2312 VGND.t2311 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6962 a_53660_17272# a_53572_17316# VGND.t2581 VGND.t2580 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6963 a_5052_21976# a_4964_22020# VGND.t4344 VGND.t4343 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6964 a_45012_29816# a_45456_30301.t5 a_45408_30345# VGND.t137 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X6965 a_46716_2727# a_46628_2824# VGND.t482 VGND.t481 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6966 VPWR.t5182 a_65756_5863# a_65668_5960# VPWR.t3689 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6967 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t2912 VPWR.t2271 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X6968 _435_.ZN _434_.ZN VGND.t1213 VGND.t1212 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X6969 _371_.A1.t4 _460_.Q VPWR.t3472 VPWR.t3471 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X6970 VPWR.t861 a_41788_2727# a_41700_2824# VPWR.t860 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6971 a_32604_18407# a_32516_18504# VGND.t5612 VGND.t4983 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6972 a_49764_23588# _398_.C VPWR.t3304 VPWR.t3303 pfet_06v0 ad=0.3534p pd=1.76u as=0.3534p ps=1.76u w=1.14u l=0.5u
X6973 _284_.B _397_.A1.t14 a_48560_26369# VPWR.t20 pfet_06v0 ad=0.2847p pd=1.615u as=0.33945p ps=1.715u w=1.095u l=0.5u
X6974 a_63068_15704# a_62980_15748# VGND.t2543 VGND.t2542 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6975 VPWR.t863 a_65756_2727# a_65668_2824# VPWR.t862 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6976 a_64636_12568# a_64548_12612# VGND.t2825 VGND.t2824 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6977 a_26720_30301# a_26427_29977# VPWR.t5219 VPWR.t5218 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X6978 VPWR.t3425 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I VPWR.t3424 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6979 VPWR.t2143 a_67324_14136# a_67236_14180# VPWR.t2142 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6980 a_31260_17272# a_31172_17316# VGND.t1940 VGND.t1939 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6981 a_50468_29977# _409_.ZN a_49600_30180# VPWR.t4911 pfet_06v0 ad=54f pd=0.66u as=0.1872p ps=1.4u w=0.36u l=0.5u
X6982 VPWR.t272 clkbuf_1_0__f_clk.I.t57 a_42392_22825.t0 VPWR.t271 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X6983 a_29828_26344# _336_.Z _358_.A2 VPWR.t4557 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X6984 VPWR.t6084 a_67324_11000# a_67236_11044# VPWR.t6083 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6985 a_28348_21543# a_28260_21640# VGND.t5927 VGND.t5926 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6986 VPWR.t5860 a_59484_2727# a_59396_2824# VPWR.t5859 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6987 a_60401_30300# _246_.B2 VGND.t5053 VGND.t1077 nfet_06v0 ad=93.59999f pd=0.88u as=0.2288p ps=1.58u w=0.36u l=0.6u
X6988 a_55004_14136# a_54916_14180# VGND.t447 VGND.t446 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6989 VPWR.t2104 a_39548_1592# a_39460_1636# VPWR.t2103 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6990 VPWR.t2866 a_3708_12135# a_3620_12232# VPWR.t2865 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6991 a_38816_27555# a_38523_27967# VGND.t985 VGND.t984 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X6992 VPWR.t34 _284_.A2.t8 a_44500_25156# VPWR.t33 pfet_06v0 ad=0.2847p pd=1.615u as=0.3942p ps=1.815u w=1.095u l=0.5u
X6993 VPWR.t2825 vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I VPWR.t2824 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X6994 a_55004_11000# a_54916_11044# VGND.t673 VGND.t672 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6995 VPWR.t5864 a_6172_2727# a_6084_2824# VPWR.t5863 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6996 VPWR.t2108 a_54892_23544# a_54804_23588# VPWR.t2107 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6997 VPWR.t5249 a_40040_17675# _452_.Q.t0 VPWR.t5248 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X6998 VPWR.t5443 a_52764_27815# a_52676_27912# VPWR.t5442 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6999 a_44700_1159# a_44612_1256# VGND.t904 VGND.t903 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7000 a_5052_15704# a_4964_15748# VGND.t2488 VGND.t2487 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7001 a_43392_19369# a_42392_19243# VGND.t586 VGND.t585 nfet_06v0 ad=43.2f pd=0.6u as=0.142p ps=1.14u w=0.36u l=0.6u
X7002 a_37084_25112# a_36996_25156# VGND.t1796 VGND.t1795 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7003 a_66652_9432# a_66564_9476# VGND.t1798 VGND.t1797 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7004 VGND.t4050 a_29184_25597# a_29136_25641# VGND.t4049 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X7005 VGND.t4958 vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN VGND.t4957 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7006 a_15132_29816# a_15044_29860# VGND.t6763 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7007 VGND.t5687 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN VGND.t5686 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7008 VPWR.t2098 a_18828_23544# a_18740_23588# VPWR.t2097 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7009 a_60405_30644# a_60285_30600# VGND.t349 VGND.t45 nfet_06v0 ad=43.8f pd=0.605u as=0.28262p ps=1.87u w=0.365u l=0.6u
X7010 a_66652_6296# a_66564_6340# VGND.t5315 VGND.t2594 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7011 VPWR.t2100 a_61276_1592# a_61188_1636# VPWR.t2099 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7012 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I VPWR.t5175 VPWR.t5174 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7013 uo_out[2].t4 _287_.A1.t34 VGND.t6494 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7014 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t2570 VPWR.t2569 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7015 a_5052_3160# a_4964_3204# VGND.t5118 VGND.t5117 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7016 VGND.t6412 vgaringosc.workerclkbuff_notouch_.I.t10 a_41048_29816.t4 VGND.t6409 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X7017 a_62060_20408# a_61972_20452# VGND.t5142 VGND.t5141 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7018 a_56836_27208# _241_.I0 VGND.t3737 VGND.t3736 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7019 a_27676_26680# a_27588_26724# VGND.t3186 VGND.t3185 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7020 VPWR.t6169 a_38316_20408# a_38228_20452# VPWR.t6168 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7021 a_3708_27815# a_3620_27912# VGND.t3010 VGND.t3009 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7022 a_1468_13703# a_1380_13800# VGND.t3723 VGND.t1764 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7023 _399_.A2 _398_.C VGND.t3150 VGND.t3149 nfet_06v0 ad=0.1339p pd=1.035u as=0.1339p ps=1.035u w=0.515u l=0.6u
X7024 VPWR.t6235 a_27116_20408# a_27028_20452# VPWR.t6234 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7025 VPWR.t595 a_55340_26680# a_55252_26724# VPWR.t594 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7026 VPWR.t3431 a_4156_29383# a_4068_29480# VPWR.t3430 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7027 a_53324_13703# a_53236_13800# VGND.t3116 VGND.t3115 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7028 VPWR.t2364 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN VPWR.t2363 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7029 _424_.ZN _424_.B1.t14 a_52436_18884# VPWR.t6619 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7030 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I VPWR.t3420 VPWR.t3066 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7031 a_49492_18840# a_49936_19325.t5 a_49888_19369# VGND.t125 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X7032 a_50860_18407# a_50772_18504# VGND.t1360 VGND.t1359 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7033 VPWR.t1225 a_48508_13703# a_48420_13800# VPWR.t1224 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7034 VPWR.t5106 a_63964_18407# a_63876_18504# VPWR.t58 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7035 VPWR.t1444 a_4156_26247# a_4068_26344# VPWR.t1443 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7036 VPWR.t4961 a_38472_30169# _287_.A1.t1 VPWR.t4960 pfet_06v0 ad=0.428p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7037 VPWR.t601 a_20172_25112# a_20084_25156# VPWR.t600 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7038 VGND.t2456 a_27668_31048# uio_out[1].t0 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7039 VPWR.t6173 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I VPWR.t6172 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7040 VPWR.t5108 a_60716_10567# a_60628_10664# VPWR.t5107 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7041 a_34980_22895# _304_.A1.t15 VPWR.t6608 VPWR.t6607 pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X7042 VPWR.t1446 a_4156_23111# a_4068_23208# VPWR.t1445 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7043 vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN VPWR.t5491 VPWR.t5490 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7044 _251_.A1.t0 a_63616_31128# VPWR.t6140 VPWR.t6139 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7045 a_15580_1592# a_15492_1636# VGND.t1548 VGND.t1272 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7046 a_48284_15704# a_48196_15748# VGND.t1550 VGND.t1549 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7047 a_2812_8999# a_2724_9096# VGND.t4075 VGND.t4074 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7048 a_49852_12568# a_49764_12612# VGND.t3998 VGND.t3997 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7049 VPWR.t4428 a_53436_18840# a_53348_18884# VPWR.t4427 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7050 _474_.CLK.t29 a_48272_25156.t43 VPWR.t6571 VPWR.t6570 pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X7051 _284_.B _381_.A2.t6 a_47636_25940# VGND.t6662 nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7052 a_9084_2727# a_8996_2824# VGND.t4624 VGND.t4623 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7053 a_62732_26680# a_62644_26724# VGND.t3291 VGND.t3290 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7054 a_37084_15704# a_36996_15748# VGND.t3743 VGND.t3742 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7055 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN VGND.t2401 VGND.t2400 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7056 a_2812_5863# a_2724_5960# VGND.t763 VGND.t762 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7057 a_58028_17272# a_57940_17316# VGND.t6044 VGND.t6043 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7058 a_2812_28248# a_2724_28292# VGND.t5936 VGND.t458 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7059 _455_.D _346_.ZN VGND.t4375 VGND.t4374 nfet_06v0 ad=0.2569p pd=1.56u as=0.2244p ps=1.9u w=0.51u l=0.6u
X7060 VPWR.t7078 a_5500_29816# a_5412_29860# VPWR.t7077 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7061 VPWR.t5083 a_61500_9432# a_61412_9476# VPWR.t5082 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7062 VPWR.t6994 _352_.A2.t28 a_27172_24328# VPWR.t6993 pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X7063 VPWR.t3553 a_22300_1159# a_22212_1256# VPWR.t3552 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7064 a_1020_20408# a_932_20452# VGND.t3840 VGND.t3839 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7065 _281_.ZN.t2 _476_.Q VPWR.t4321 VPWR.t4320 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X7066 a_48908_24080# _474_.Q _399_.A2 VGND.t4643 nfet_06v0 ad=93.59999f pd=1.02u as=0.2028p ps=1.3u w=0.78u l=0.6u
X7067 VPWR.t663 a_8188_1592# a_8100_1636# VPWR.t662 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7068 VPWR.t424 a_42236_15704# a_42148_15748# VPWR.t423 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7069 a_26954_28776# _455_.Q.t14 a_26750_28776# VGND.t6540 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7070 a_42368_28733# a_41996_28777# VGND.t2839 VGND.t2838 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X7071 VPWR.t418 a_33500_16839# a_33412_16936# VPWR.t417 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7072 VPWR.t1452 a_54108_15271# a_54020_15368# VPWR.t1451 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7073 VGND.t3427 _371_.A2 _371_.ZN VGND.t3426 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7074 a_42012_1592# a_41924_1636# VGND.t2164 VGND.t2163 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7075 a_37384_19624# _448_.Q.t13 a_37772_19759# VGND.t6579 nfet_06v0 ad=0.1606p pd=1.61u as=58.39999f ps=0.685u w=0.365u l=0.6u
X7076 VPWR.t923 a_58588_26247# a_58500_26344# VPWR.t922 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7077 a_49292_12135# a_49204_12232# VGND.t2702 VGND.t2701 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7078 _325_.ZN _325_.B VGND.t2627 VGND.t2626 nfet_06v0 ad=0.2569p pd=1.56u as=0.2244p ps=1.9u w=0.51u l=0.6u
X7079 VPWR.t714 a_63516_17272# a_63428_17316# VPWR.t713 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7080 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN VPWR.t536 VPWR.t535 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7081 VPWR.t404 a_18096_27165# uio_out[7].t2 VPWR.t403 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X7082 a_46268_12135# a_46180_12232# VGND.t3236 VGND.t2339 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7083 a_35068_15271# a_34980_15368# VGND.t3563 VGND.t3562 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7084 VPWR.t3986 a_1020_21976# a_932_22020# VPWR.t328 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7085 VGND.t6407 a_41048_29816.t19 _459_.CLK.t9 VGND.t6400 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X7086 VPWR.t741 a_52316_17272# a_52228_17316# VPWR.t740 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7087 VGND.t2722 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN VGND.t2721 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7088 VPWR.t2971 a_20508_2727# a_20420_2824# VPWR.t2970 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7089 VPWR.t929 a_36188_26247# a_36100_26344# VPWR.t928 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7090 a_19276_25112# a_19188_25156# VGND.t3975 VGND.t3974 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7091 a_44700_2727# a_44612_2824# VGND.t924 VGND.t923 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7092 a_39100_15704# a_39012_15748# VGND.t2256 VGND.t2255 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7093 a_36288_23208# _311_.Z a_36084_23208# VPWR.t4472 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7094 a_19276_21976# a_19188_22020# VGND.t4479 VGND.t4478 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7095 VGND.t1060 a_65072_29860# _324_.C.t4 VGND.t1059 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X7096 VPWR.t2975 a_63740_2727# a_63652_2824# VPWR.t2974 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7097 a_48508_1592# a_48420_1636# VGND.t2093 VGND.t2092 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7098 VPWR.t2410 a_43804_1592# a_43716_1636# VPWR.t2409 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7099 VPWR.t7074 a_5388_19975# a_5300_20072# VPWR.t7073 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7100 VPWR.t2977 a_14236_2727# a_14148_2824# VPWR.t2976 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7101 a_49740_13703# a_49652_13800# VGND.t1757 VGND.t1756 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7102 a_1020_14136# a_932_14180# VGND.t4618 VGND.t3193 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7103 VGND.t1926 _287_.A2 uo_out[6].t0 VGND.t1925 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7104 VPWR.t5320 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I VPWR.t5319 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7105 a_2812_18840# a_2724_18884# VGND.t3077 VGND.t3076 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7106 a_62560_25112# _251_.A1.t35 VPWR.t7026 VPWR.t7025 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7107 a_67772_1592# a_67684_1636# VGND.t2073 VGND.t2072 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7108 VPWR.t1448 a_66764_13703# a_66676_13800# VPWR.t1447 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7109 a_1020_11000# a_932_11044# VGND.t4373 VGND.t4372 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7110 a_46716_13703# a_46628_13800# VGND.t342 VGND.t341 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7111 VPWR.t4416 a_50524_1159# a_50436_1256# VPWR.t4415 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7112 VPWR.t1450 a_55564_13703# a_55476_13800# VPWR.t1449 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7113 VPWR.t6149 a_37532_26680# a_37444_26724# VPWR.t490 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7114 VPWR.t6893 _448_.Q.t14 _261_.ZN VPWR.t6892 pfet_06v0 ad=0.2561p pd=1.505u as=0.4016p ps=1.94u w=0.985u l=0.5u
X7115 a_30028_20408# a_29940_20452# VGND.t4736 VGND.t4735 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7116 _435_.ZN _437_.A1.t13 VGND.t6552 VGND.t6551 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7117 VPWR.t7081 a_15132_29816# a_15044_29860# VPWR.t3501 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7118 a_19724_23544# a_19636_23588# VGND.t1739 VGND.t1738 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7119 a_58252_18407# a_58164_18504# VGND.t4266 VGND.t4265 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7120 a_34592_20569# a_34160_20523# VPWR.t2899 VPWR.t2898 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X7121 VPWR.t937 _384_.A1 _398_.C VPWR.t936 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7122 VPWR.t5148 a_44252_1159# a_44164_1256# VPWR.t1251 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7123 VPWR.t4196 a_67772_14136# a_67684_14180# VPWR.t4195 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7124 a_62508_21976# a_62420_22020# VGND.t5155 VGND.t2638 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7125 VPWR.t2203 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN VPWR.t2202 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7126 VPWR.t3551 a_68108_10567# a_68020_10664# VPWR.t3550 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7127 VPWR.t2633 a_38652_15704# a_38564_15748# VPWR.t2632 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7128 a_30388_28776# _337_.ZN _350_.A2.t4 VGND.t4977 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7129 VPWR.t3032 a_67772_11000# a_67684_11044# VPWR.t3031 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7130 VPWR.t3555 a_39996_2727# a_39908_2824# VPWR.t3554 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7131 VPWR.t3034 a_3708_20408# a_3620_20452# VPWR.t3033 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7132 VPWR.t4564 a_51240_19624# _476_.Q VPWR.t4563 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7133 a_28796_21543# a_28708_21640# VGND.t3878 VGND.t3877 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7134 vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN VPWR.t3735 VPWR.t3734 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7135 a_55452_14136# a_55364_14180# VGND.t4769 VGND.t2159 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7136 VPWR.t3038 a_45372_14136# a_45284_14180# VPWR.t3037 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7137 VPWR.t1386 a_27004_23111# a_26916_23208# VPWR.t1385 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7138 VPWR.t5465 a_3708_4295# a_3620_4392# VPWR.t5464 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7139 a_2812_1159# a_2724_1256# VGND.t70 VGND.t69 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7140 VPWR.t5814 _301_.Z a_38576_22504# VPWR.t5813 pfet_06v0 ad=0.395p pd=2.02u as=0.156p ps=1.12u w=0.6u l=0.5u
X7141 a_23868_1159# a_23780_1256# VGND.t2833 VGND.t2832 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7142 a_55312_22340# a_54864_22461.t7 a_55724_22137# VPWR.t6598 pfet_06v0 ad=0.1872p pd=1.4u as=43.2f ps=0.6u w=0.36u l=0.5u
X7143 a_39796_22504# _301_.A1 _261_.ZN VGND.t3199 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7144 a_19164_26247# a_19076_26344# VGND.t3306 VGND.t3305 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7145 a_41264_30669# _388_.B a_41056_30669# VGND.t4150 nfet_06v0 ad=57.59999f pd=0.68u as=0.1584p ps=1.6u w=0.36u l=0.6u
X7146 VGND.t1848 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN VGND.t1847 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7147 a_25643_25273# a_23668_25640.t7 a_25008_25597# VPWR.t7030 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X7148 a_55452_11000# a_55364_11044# VGND.t4771 VGND.t4770 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7149 VPWR.t1305 a_39324_15271# a_39236_15368# VPWR.t1304 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7150 VGND.t6297 _350_.A2.t28 a_29371_30644# VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7151 VPWR.t3363 a_45372_11000# a_45284_11044# VPWR.t346 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7152 VPWR.t745 a_58140_12568# a_58052_12612# VPWR.t744 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7153 a_40264_30320# _285_.Z VPWR.t5930 VPWR.t5929 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X7154 a_62279_28293# _250_.C VPWR.t5059 VPWR.t5058 pfet_06v0 ad=0.37665p pd=1.835u as=0.5346p ps=3.31u w=1.215u l=0.5u
X7155 VPWR.t1374 a_3708_1159# a_3620_1256# VPWR.t649 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7156 a_19164_23111# a_19076_23208# VGND.t1529 VGND.t1528 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7157 VPWR.t3532 a_33776_29123# a_33768_29535# VPWR.t3531 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X7158 VPWR.t4333 a_24988_21543# a_24900_21640# VPWR.t4332 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7159 clkbuf_1_0__f_clk.I.t1 a_44296_24393.t41 VPWR.t296 VPWR.t295 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7160 VPWR.t2260 a_51576_25896# _397_.A1.t0 VPWR.t2259 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7161 a_59955_30600# a_60285_30600# a_60405_31198# VPWR.t358 pfet_06v0 ad=0.3456p pd=2.64u as=61.19999f ps=0.7u w=0.36u l=0.5u
X7162 input9.Z a_52639_30644# VGND.t3985 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.28262p ps=1.87u w=0.82u l=0.6u
X7163 VPWR.t971 a_60276_29032# _257_.B VPWR.t970 pfet_06v0 ad=0.389p pd=2.02u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7164 VPWR.t771 a_48732_17272# a_48644_17316# VPWR.t770 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7165 VGND.t3425 _371_.A2 _352_.A2.t4 VGND.t3424 nfet_06v0 ad=0.1326p pd=1.03u as=0.1326p ps=1.03u w=0.51u l=0.6u
X7166 a_66652_2727# a_66564_2824# VGND.t5204 VGND.t5203 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7167 a_46476_20937# _475_.D a_46308_20937# VGND.t4314 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X7168 a_2812_30951# a_2724_31048# VGND.t3112 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7169 a_17148_2727# a_17060_2824# VGND.t1137 VGND.t1136 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7170 VPWR.t6102 a_17168_27165# a_17140_26841# VPWR.t6101 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X7171 VPWR.t998 a_65756_4728# a_65668_4772# VPWR.t997 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7172 a_15580_29816# a_15492_29860# VGND.t72 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7173 VPWR.t573 a_37532_17272# a_37444_17316# VPWR.t572 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7174 a_20396_27815# a_20308_27912# VGND.t5596 VGND.t2654 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7175 a_36960_27912# a_36548_27591.t7 VGND.t6328 VGND.t6327 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X7176 VPWR.t577 a_45708_17272# a_45620_17316# VPWR.t576 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7177 VPWR.t5385 a_64188_27815# a_64100_27912# VPWR.t5384 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7178 VPWR.t1313 a_21292_30951# a_21204_31048# VPWR.t1312 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7179 VPWR.t726 a_36188_2727# a_36100_2824# VPWR.t725 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7180 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t1078 VPWR.t1077 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7181 a_54332_15704# a_54244_15748# VGND.t4547 VGND.t4546 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7182 a_2364_26247# a_2276_26344# VGND.t5331 VGND.t5330 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7183 a_67100_17272# a_67012_17316# VGND.t1974 VGND.t1973 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7184 VPWR.t6491 _459_.CLK.t42 a_18404_30344.t0 VPWR.t6490 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X7185 a_55900_12568# a_55812_12612# VGND.t3443 VGND.t3442 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7186 VPWR.t1689 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I VPWR.t1688 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7187 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I VPWR.t4482 VPWR.t4481 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7188 VPWR.t1132 a_10092_30951# a_10004_31048# VPWR.t1131 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7189 uio_out[7].t1 a_18096_27165# VPWR.t402 VPWR.t401 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7190 VGND.t2278 vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I VGND.t2277 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7191 a_19612_24679# a_19524_24776# VGND.t5337 VGND.t5336 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7192 VPWR.t3982 a_3708_14136# a_3620_14180# VPWR.t801 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7193 a_43132_15704# a_43044_15748# VGND.t2111 VGND.t2110 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7194 a_2364_23111# a_2276_23208# VGND.t2978 VGND.t2977 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7195 VPWR.t1529 _249_.A2 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I VPWR.t1528 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7196 VPWR.t3199 a_38764_20408# a_38676_20452# VPWR.t3198 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7197 a_64972_13703# a_64884_13800# VGND.t3029 VGND.t3028 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7198 VPWR.t1066 a_59484_1592# a_59396_1636# VPWR.t1065 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7199 VGND.t5028 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I VGND.t5027 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7200 a_19612_21543# a_19524_21640# VGND.t973 VGND.t972 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7201 VPWR.t3201 a_3708_11000# a_3620_11044# VPWR.t1026 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7202 a_4604_7864# a_4516_7908# VGND.t74 VGND.t73 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7203 VPWR.t3686 a_27564_20408# a_27476_20452# VPWR.t3685 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7204 _260_.A1 _327_.A2 VGND.t3246 VGND.t3245 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X7205 a_53772_13703# a_53684_13800# VGND.t3261 VGND.t3260 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7206 a_65308_3160# a_65220_3204# VGND.t3750 VGND.t670 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7207 VPWR.t7076 a_61276_19975# a_61188_20072# VPWR.t7075 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7208 a_4604_4728# a_4516_4772# VGND.t4179 VGND.t4178 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7209 a_51420_1159# a_51332_1256# VGND.t3733 VGND.t3732 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7210 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I VPWR.t3790 VPWR.t3789 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7211 a_44784_25987.t0 _474_.CLK.t55 VPWR.t6767 VPWR.t6766 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X7212 a_63516_15271# a_63428_15368# VGND.t3904 VGND.t3903 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7213 a_60909_30600# ui_in[3].t0 VPWR.t53 VPWR.t52 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X7214 a_43814_21236# a_42982_21730# a_43666_21812# VPWR.t5437 pfet_06v0 ad=0.3852p pd=2.86u as=61.19999f ps=0.7u w=0.36u l=0.5u
X7215 VPWR.t5739 a_56964_26724# _241_.Z VPWR.t5738 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X7216 VPWR.t4678 _304_.B a_41056_30669# VPWR.t4677 pfet_06v0 ad=0.34437p pd=1.895u as=0.1456p ps=1.08u w=0.56u l=0.5u
X7217 a_15244_20408# a_15156_20452# VGND.t1042 VGND.t1041 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7218 VGND.t4019 a_44752_18147# a_44704_18191# VGND.t4018 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X7219 VGND.t5711 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7220 VGND.t2946 _369_.ZN a_29835_28776# VGND.t2945 nfet_06v0 ad=0.3124p pd=2.3u as=85.2f ps=0.95u w=0.71u l=0.6u
X7221 a_2812_24679# a_2724_24776# VGND.t1399 VGND.t1398 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7222 VGND.t5084 a_40040_17675# _452_.Q.t2 VGND.t5083 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7223 a_31168_24419# a_30796_24463# VGND.t2973 VGND.t2972 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X7224 VGND.t1537 a_46198_27060# _330_.A1.t2 VGND.t1536 nfet_06v0 ad=0.2911p pd=1.53u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7225 a_62060_10567# a_61972_10664# VGND.t4212 VGND.t4211 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7226 a_41116_15271# a_41028_15368# VGND.t1336 VGND.t1335 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7227 a_34732_19975# a_34644_20072# VGND.t76 VGND.t75 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7228 VPWR.t1768 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN VPWR.t1767 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7229 a_2812_21543# a_2724_21640# VGND.t2209 VGND.t2208 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7230 a_38968_22504# _300_.A2 a_38784_22504# VGND.t937 nfet_06v0 ad=88.2f pd=0.84u as=67.2f ps=0.74u w=0.42u l=0.6u
X7231 VPWR.t5025 a_57132_23544# a_57044_23588# VPWR.t5024 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7232 a_58340_29860# _228_.ZN _272_.A2 VPWR.t323 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X7233 a_58476_17272# a_58388_17316# VGND.t3901 VGND.t3900 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7234 VGND.t1413 a_44160_29123# a_44112_29167# VGND.t1412 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X7235 VGND.t5742 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN VGND.t5741 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7236 a_65420_16839# a_65332_16936# VGND.t5078 VGND.t5077 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7237 a_31708_19975# a_31620_20072# VGND.t78 VGND.t77 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7238 VPWR.t5031 a_42684_15704# a_42596_15748# VPWR.t5030 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7239 a_2364_16839# a_2276_16936# VGND.t3512 VGND.t3511 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7240 a_36628_29535# a_35316_29159.t6 a_36284_29167# VPWR.t7055 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X7241 a_25324_21976# a_25236_22020# VGND.t5162 VGND.t5161 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7242 a_43908_26841# a_42596_27208.t6 a_43564_27209# VPWR.t142 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X7243 VPWR.t2468 a_15244_21976# a_15156_22020# VPWR.t338 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7244 a_34516_25940# _358_.A3 VGND.t467 VGND.t466 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7245 VPWR.t7080 a_3260_19975# a_3172_20072# VPWR.t5639 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7246 a_22524_1592# a_22436_1636# VGND.t5274 VGND.t5273 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7247 VPWR.t992 a_54556_15271# a_54468_15368# VPWR.t991 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7248 VPWR.t5432 a_6620_29383# a_6532_29480# VPWR.t5431 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7249 VPWR.t994 a_31036_23111# a_30948_23208# VPWR.t993 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7250 uo_out[4].t7 _287_.A1.t35 a_33812_29860# VPWR.t6790 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7251 a_60909_30600# ui_in[3].t1 VGND.t46 VGND.t45 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7252 VPWR.t485 a_4156_28248# a_4068_28292# VPWR.t484 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7253 a_50300_20408# a_50212_20452# VGND.t4506 VGND.t4505 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7254 a_35968_20937# a_33748_20936.t7 a_35723_20569# VGND.t44 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7255 VPWR.t487 a_40220_20408# a_40132_20452# VPWR.t486 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7256 VGND.t6217 _459_.CLK.t43 a_15828_27208.t1 VGND.t6216 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X7257 a_43020_16839# a_42932_16936# VGND.t1004 VGND.t1003 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7258 a_31348_25156# _358_.A2 a_31124_25156# VPWR.t4837 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7259 VGND.t5170 a_52848_25987# a_52744_26031# VGND.t5169 nfet_06v0 ad=0.2637p pd=1.825u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7260 VPWR.t581 a_48508_12568# a_48420_12612# VPWR.t580 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7261 VPWR.t556 a_63964_17272# a_63876_17316# VPWR.t555 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7262 a_23196_23111# a_23108_23208# VGND.t3352 VGND.t3351 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7263 VPWR.t558 a_4156_25112# a_4068_25156# VPWR.t557 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7264 a_25108_27508# _346_.A2 VGND.t3483 VGND.t3482 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7265 VPWR.t1134 a_61612_13703# a_61524_13800# VPWR.t1133 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7266 a_42252_20936# _452_.Q.t20 _304_.ZN.t9 VGND.t6646 nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X7267 VPWR.t1975 a_32156_15271# a_32068_15368# VPWR.t1974 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7268 a_60084_25640# vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN VGND.t4003 VGND.t4002 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7269 _252_.B _229_.I.t13 VPWR.t6878 VPWR.t6877 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X7270 a_41880_24072# _226_.ZN a_41696_24072# VGND.t2259 nfet_06v0 ad=88.2f pd=0.84u as=67.2f ps=0.74u w=0.42u l=0.6u
X7271 VPWR.t565 a_52764_17272# a_52676_17316# VPWR.t564 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7272 _293_.A2 _285_.Z VGND.t5705 VGND.t102 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X7273 VPWR.t2917 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN VPWR.t2916 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7274 VGND.t1662 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7275 a_1020_10567# a_932_10664# VGND.t3891 VGND.t3890 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7276 a_44459_18559# a_42484_18183.t7 a_43824_18147# VPWR.t7047 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X7277 a_6620_1159# a_6532_1256# VGND.t338 VGND.t337 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7278 a_27676_1159# a_27588_1256# VGND.t3350 VGND.t3349 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7279 _467_.D _355_.C.t18 VGND.t6393 VGND.t6392 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X7280 a_53100_18407# a_53012_18504# VGND.t1527 VGND.t1526 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7281 a_34844_24679# a_34756_24776# VGND.t2490 VGND.t2489 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7282 a_33768_29535# a_31920_29480# a_33483_29535# VPWR.t3290 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X7283 VPWR.t1982 a_1916_8999# a_1828_9096# VPWR.t1981 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7284 a_18940_2727# a_18852_2824# VGND.t3986 VGND.t3163 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7285 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN VGND.t5147 VGND.t5146 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7286 _300_.A2 _448_.Q.t15 VGND.t6581 VGND.t6580 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X7287 VPWR.t3733 a_33500_18840# a_33412_18884# VPWR.t2791 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7288 _427_.B1 a_52452_24072# VPWR.t5394 VPWR.t5393 pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X7289 a_23644_24679# a_23556_24776# VGND.t1901 VGND.t1900 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7290 VGND.t3280 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I VGND.t3279 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7291 VGND.t3481 _346_.A2 a_21868_27208# VGND.t3480 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7292 VPWR.t2804 a_37980_2727# a_37892_2824# VPWR.t2803 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7293 a_61500_14136# a_61412_14180# VGND.t4394 VGND.t4393 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7294 VPWR.t1347 a_33500_15704# a_33412_15748# VPWR.t1346 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7295 a_23644_21543# a_23556_21640# VGND.t4025 VGND.t4024 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7296 VGND.t3727 a_34448_25597# _460_.Q VGND.t3726 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7297 VPWR.t6493 _459_.CLK.t44 a_42820_29159.t1 VPWR.t6492 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X7298 a_61500_11000# a_61412_11044# VGND.t4398 VGND.t4397 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7299 VPWR.t81 a_4604_7864# a_4516_7908# VPWR.t80 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7300 a_50300_14136# a_50212_14180# VGND.t4399 VGND.t373 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7301 a_46171_27508# _324_.C.t32 _403_.ZN VGND.t233 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7302 a_48732_15271# a_48644_15368# VGND.t4706 VGND.t4705 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7303 a_64860_7431# a_64772_7528# VGND.t5979 VGND.t2699 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7304 _371_.A3 _223_.I VPWR.t7110 VPWR.t7109 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X7305 a_30476_20408# a_30388_20452# VGND.t4353 VGND.t4352 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7306 VPWR.t6948 a_49152_30301.t7 a_49112_29885# VPWR.t6947 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X7307 VPWR.t1074 a_20396_20408# a_20308_20452# VPWR.t1073 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7308 a_50300_11000# a_50212_11044# VGND.t4357 VGND.t4356 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7309 a_21404_2727# a_21316_2824# VGND.t3725 VGND.t3724 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7310 VPWR.t1662 a_24764_1159# a_24676_1256# VPWR.t1661 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7311 a_47297_25596# _279_.Z VGND.t5384 VGND.t5383 nfet_06v0 ad=93.59999f pd=0.88u as=0.2288p ps=1.58u w=0.36u l=0.6u
X7312 VPWR.t79 a_15580_29816# a_15492_29860# VPWR.t78 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7313 a_50748_1592# a_50660_1636# VGND.t4485 VGND.t4484 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7314 VPWR.t2806 a_47297_25596# _381_.A2.t0 VPWR.t2805 pfet_06v0 ad=0.38705p pd=2.08u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7315 VPWR.t5307 a_64412_5863# a_64324_5960# VPWR.t5306 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7316 VGND.t6190 a_43440_19325.t6 a_43400_18909# VGND.t6189 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X7317 a_38752_26344# _437_.A1.t14 VPWR.t6864 VPWR.t6863 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7318 a_35728_29480# a_35316_29159.t7 VPWR.t7057 VPWR.t7056 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X7319 VPWR.t2809 a_40444_2727# a_40356_2824# VPWR.t2808 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7320 _323_.A3 _319_.A3 VGND.t2568 VGND.t2567 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X7321 a_46084_19759# a_45284_19751.t5 VGND.t6714 VGND.t6713 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X7322 VPWR.t1538 a_36188_25112# a_36100_25156# VPWR.t1537 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7323 _311_.Z a_34980_22895# VPWR.t3224 VPWR.t3223 pfet_06v0 ad=0.5346p pd=3.31u as=0.40575p ps=2.055u w=1.215u l=0.5u
X7324 VPWR.t1546 a_57692_9432# a_57604_9476# VPWR.t1545 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7325 a_15132_2727# a_15044_2824# VGND.t3787 VGND.t3297 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7326 VPWR.t5417 a_16252_29383# a_16164_29480# VPWR.t5416 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7327 VPWR.t5664 a_18492_1159# a_18404_1256# VPWR.t1190 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7328 _342_.ZN _355_.C.t19 a_24304_29480# VPWR.t6680 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7329 a_40676_25640# _261_.ZN VGND.t3417 VGND.t3416 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7330 a_52428_10567# a_52340_10664# VGND.t3638 VGND.t3637 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7331 a_39100_2727# a_39012_2824# VGND.t3162 VGND.t3161 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7332 VGND.t4918 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN VGND.t4917 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7333 a_44028_25156# _284_.A2.t9 VPWR.t36 VPWR.t35 pfet_06v0 ad=0.4599p pd=1.935u as=0.3766p ps=1.815u w=1.095u l=0.5u
X7334 VPWR.t2817 a_34172_2727# a_34084_2824# VPWR.t2816 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7335 VPWR.t1283 a_63740_1592# a_63652_1636# VPWR.t1282 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7336 VPWR.t824 a_27452_23111# a_27364_23208# VPWR.t823 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7337 VPWR.t1285 a_14236_1592# a_14148_1636# VPWR.t1284 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7338 VGND.t6521 _325_.A1.t21 a_40452_22504# VGND.t6520 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7339 vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN VPWR.t4156 VPWR.t4155 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7340 a_1468_8999# a_1380_9096# VGND.t2440 VGND.t2439 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7341 a_63740_1159# a_63652_1256# VGND.t4799 VGND.t4798 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7342 VPWR.t1179 a_30476_21976# a_30388_22020# VPWR.t1178 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7343 a_29563_29535# a_28000_29480# a_28928_29123# VGND.t1837 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7344 a_67237_30644# a_67117_30600# VGND.t3176 VGND.t45 nfet_06v0 ad=43.8f pd=0.605u as=0.28262p ps=1.87u w=0.365u l=0.6u
X7345 VPWR.t868 a_58140_2727# a_58052_2824# VPWR.t867 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7346 VPWR.t828 a_39772_15271# a_39684_15368# VPWR.t827 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7347 a_3260_29383# a_3172_29480# VGND.t3602 VGND.t2767 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7348 VPWR.t636 a_38204_1592# a_38116_1636# VPWR.t635 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7349 VGND.t2376 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN VGND.t2375 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7350 VPWR.t22 _397_.A1.t15 _386_.A4 VPWR.t21 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7351 a_1468_5863# a_1380_5960# VGND.t3603 VGND.t2772 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7352 a_16588_26247# a_16500_26344# VGND.t2492 VGND.t2491 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7353 VPWR.t870 a_63180_16839# a_63092_16936# VPWR.t869 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7354 a_40636_18180# _452_.Q.t21 a_40452_18180# VGND.t6647 nfet_06v0 ad=79.8f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X7355 clkbuf_1_0__f_clk.I.t0 a_44296_24393.t42 VPWR.t298 VPWR.t297 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7356 VPWR.t6717 _324_.B.t33 _424_.A2.t0 VPWR.t6716 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7357 a_16588_23111# a_16500_23208# VGND.t1562 VGND.t1561 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7358 _422_.ZN _419_.Z VPWR.t4461 VPWR.t4460 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X7359 VPWR.t1025 a_22412_20408# a_22324_20452# VPWR.t1024 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7360 VPWR.t872 a_38316_16839# a_38228_16936# VPWR.t871 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7361 VPWR.t1556 a_37980_17272# a_37892_17316# VPWR.t1555 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7362 a_1916_25112# a_1828_25156# VGND.t1317 VGND.t1316 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7363 VPWR.t5451 a_48060_12135# a_47972_12232# VPWR.t4100 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7364 a_54780_15704# a_54692_15748# VGND.t2635 VGND.t2634 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7365 VPWR.t438 a_52024_20083# a_53380_20127# VPWR.t437 pfet_06v0 ad=0.4554p pd=3.25u as=54f ps=0.66u w=0.36u l=0.5u
X7366 a_1916_21976# a_1828_22020# VGND.t4473 VGND.t4185 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7367 _260_.ZN _260_.A1 VPWR.t3912 VPWR.t3911 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X7368 VPWR.t6695 a_41048_29816.t20 _459_.CLK.t1 VPWR.t6694 pfet_06v0 ad=0.367p pd=1.92u as=0.4392p ps=1.94u w=1.22u l=0.5u
X7369 VPWR.t4858 a_1020_27815# a_932_27912# VPWR.t697 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7370 a_1020_1159# a_932_1256# VGND.t1443 VGND.t1442 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7371 a_43580_15704# a_43492_15748# VGND.t2079 VGND.t2078 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7372 VGND.t775 _223_.ZN a_32476_28776# VGND.t774 nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7373 a_67548_7431# a_67460_7528# VGND.t1322 VGND.t1321 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7374 VGND.t2919 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN VGND.t2918 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7375 a_1468_17272# a_1380_17316# VGND.t5536 VGND.t3507 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7376 a_42168_22504# _305_.A2 _324_.B.t0 VGND.t2873 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7377 VPWR.t6495 _459_.CLK.t45 a_17060_28776.t0 VPWR.t6494 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X7378 a_43356_2727# a_43268_2824# VGND.t5378 VGND.t1971 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7379 a_67324_12568# a_67236_12612# VGND.t1628 VGND.t1627 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7380 VPWR.t4532 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN VPWR.t4531 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7381 a_31031_27208# _459_.Q.t16 a_30847_27208# VGND.t6661 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7382 a_63964_15271# a_63876_15368# VGND.t5108 VGND.t5107 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7383 vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN VPWR.t5188 VPWR.t5187 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7384 VPWR.t65 a_62396_2727# a_62308_2824# VPWR.t64 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7385 a_15692_20408# a_15604_20452# VGND.t4116 VGND.t3165 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7386 a_59380_27508# _243_.ZN VGND.t3887 VGND.t3886 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7387 a_35008_27533# _363_.Z.t9 VPWR.t47 VPWR.t46 pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X7388 VGND.t6781 a_49068_20408# _419_.Z VGND.t6780 nfet_06v0 ad=0.226p pd=1.515u as=0.3586p ps=2.51u w=0.815u l=0.6u
X7389 _319_.ZN _319_.A2 VGND.t1127 VGND.t1126 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7390 _452_.CLK.t27 a_42392_22825.t41 VPWR.t6938 VPWR.t6937 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7391 a_37084_2727# a_36996_2824# VGND.t3873 VGND.t3872 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7392 VPWR.t378 a_66428_1592# a_66340_1636# VPWR.t377 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7393 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I VGND.t3834 VGND.t3833 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7394 VGND.t6219 _459_.CLK.t46 a_27588_29159.t1 VGND.t6218 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X7395 a_28388_29167# a_27588_29159.t7 VGND.t6559 VGND.t6558 nfet_06v0 ad=43.2f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X7396 a_39996_1159# a_39908_1256# VGND.t4748 VGND.t4747 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7397 VPWR.t859 a_5276_30951# a_5188_31048# VPWR.t858 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7398 a_43246_24163# a_43126_24119# VGND.t3215 VGND.t3214 nfet_06v0 ad=43.8f pd=0.605u as=0.28262p ps=1.87u w=0.365u l=0.6u
X7399 a_41564_15271# a_41476_15368# VGND.t2509 VGND.t2508 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7400 VPWR.t1223 a_57580_23544# a_57492_23588# VPWR.t1222 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7401 a_44340_26183# a_44744_26355# a_44688_26399# VPWR.t6296 pfet_06v0 ad=0.1665p pd=1.285u as=50.4f ps=0.64u w=0.36u l=0.5u
X7402 a_1916_15704# a_1828_15748# VGND.t1938 VGND.t1937 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7403 VPWR.t4499 vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I VPWR.t4498 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7404 a_40973_24776# _436_.B a_40357_24776# VPWR.t5868 pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X7405 VPWR.t226 _324_.C.t33 _393_.A3 VPWR.t225 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7406 a_25772_21976# a_25684_22020# VGND.t4677 VGND.t4676 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7407 VPWR.t6137 a_15692_21976# a_15604_22020# VPWR.t5546 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7408 a_40468_25157# _260_.A1 _264_.B VPWR.t3910 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X7409 a_44795_29535# a_43232_29480# a_44160_29123# VGND.t788 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7410 VPWR.t69 a_1020_18407# a_932_18504# VPWR.t68 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7411 VPWR.t5862 a_31484_23111# a_31396_23208# VPWR.t5861 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7412 _399_.ZN _399_.A2 a_48321_23208# VPWR.t1472 pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X7413 a_4828_29383# a_4740_29480# VGND.t3049 VGND.t3048 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7414 VPWR.t5497 a_41228_27815# a_41140_27912# VPWR.t5496 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7415 VPWR.t73 a_50188_10567# a_50100_10664# VPWR.t72 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7416 VPWR.t75 a_16700_2727# a_16612_2824# VPWR.t74 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7417 VPWR.t6610 _304_.A1.t16 a_36148_21976# VPWR.t6609 pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X7418 a_63292_9432# a_63204_9476# VGND.t2720 VGND.t2719 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7419 VPWR.t5627 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I VPWR.t5626 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7420 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN VGND.t5710 VGND.t71 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7421 VPWR.t5591 _284_.B _284_.ZN.t16 VPWR.t5590 pfet_06v0 ad=0.3766p pd=1.815u as=0.2561p ps=1.505u w=0.985u l=0.5u
X7422 VPWR.t3396 _327_.A2 a_41188_18840# VPWR.t3395 pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X7423 VPWR.t1562 a_48956_12568# a_48868_12612# VPWR.t1561 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7424 VGND.t6378 _452_.CLK.t58 a_36996_18183.t1 VGND.t6377 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X7425 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I _274_.A1 VPWR.t2653 VPWR.t2652 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7426 VPWR.t7084 a_53548_16839# a_53460_16936# VPWR.t7083 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7427 VPWR.t6461 a_43440_19325.t7 a_43400_18909# VPWR.t6460 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X7428 a_67212_13703# a_67124_13800# VGND.t4757 VGND.t4756 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7429 a_4156_13703# a_4068_13800# VGND.t5052 VGND.t2126 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7430 a_27552_24397# _336_.A2.t13 VGND.t170 VGND.t169 nfet_06v0 ad=57.59999f pd=0.68u as=0.218p ps=1.52u w=0.36u l=0.6u
X7431 a_56012_13703# a_55924_13800# VGND.t2166 VGND.t2165 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7432 a_47504_19759# a_45284_19751.t6 a_47259_20127# VGND.t6715 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7433 a_1020_29816# a_932_29860# VGND.t79 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7434 VPWR.t5173 a_60268_12135# a_60180_12232# VPWR.t5172 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7435 VGND.t6221 _459_.CLK.t47 a_41028_28776.t1 VGND.t6220 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X7436 a_7628_30951# a_7540_31048# VGND.t1626 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7437 a_61724_18407# a_61636_18504# VGND.t3916 VGND.t3915 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7438 a_18372_28409# a_17060_28776.t7 a_18028_28777# VPWR.t6908 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X7439 _360_.ZN _460_.Q a_33396_26344# VPWR.t3470 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7440 VPWR.t7086 a_63404_10567# a_63316_10664# VPWR.t7085 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7441 a_42460_1592# a_42372_1636# VGND.t1753 VGND.t1752 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7442 _459_.CLK.t8 a_41048_29816.t21 VGND.t6408 VGND.t6400 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X7443 a_33948_15704# a_33860_15748# VGND.t1914 VGND.t1132 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7444 _427_.ZN _427_.B1 a_52660_21640# VPWR.t3960 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7445 _459_.CLK.t0 a_41048_29816.t22 VPWR.t6697 VPWR.t6696 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7446 a_36860_23111# a_36772_23208# VGND.t1586 VGND.t1585 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7447 VPWR.t1315 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t1314 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7448 a_59036_26247# a_58948_26344# VGND.t2460 VGND.t2459 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7449 a_2364_26680# a_2276_26724# VGND.t4205 VGND.t4204 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7450 a_48508_1159# a_48420_1256# VGND.t2667 VGND.t2666 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7451 VPWR.t5098 a_67100_8999# a_67012_9096# VPWR.t1579 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7452 VPWR.t5100 a_22300_23111# a_22212_23208# VPWR.t5099 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7453 VPWR.t7087 a_3708_16839# a_3620_16936# VPWR.t5242 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7454 VPWR.t1119 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN VPWR.t1118 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7455 VPWR.t7089 a_14796_24679# a_14708_24776# VPWR.t3600 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7456 VPWR.t7088 a_33052_18407# a_32964_18504# VPWR.t4712 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7457 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN VPWR.t3423 VPWR.t3422 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7458 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN VGND.t1661 VGND.t34 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7459 VGND.t6248 _284_.ZN.t36 uo_out[1].t2 VGND.t6247 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7460 a_38584_28292# _437_.A1.t15 VGND.t6554 VGND.t6553 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X7461 VPWR.t5105 a_34620_15271# a_34532_15368# VPWR.t5104 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7462 VPWR.t7091 a_20956_2727# a_20868_2824# VPWR.t7090 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7463 a_29184_25597# a_28891_25273# VGND.t455 VGND.t454 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X7464 VGND.t6290 a_48272_25156.t44 _474_.CLK.t30 VGND.t6289 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X7465 a_39536_26795# a_39124_27208.t6 VPWR.t223 VPWR.t222 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X7466 a_1916_1592# a_1828_1636# VGND.t1225 VGND.t1224 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7467 a_24988_1592# a_24900_1636# VGND.t1227 VGND.t1226 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7468 a_50012_29977# a_49496_30345# VPWR.t880 VPWR.t879 pfet_06v0 ad=43.2f pd=0.6u as=0.1044p ps=0.94u w=0.36u l=0.5u
X7469 a_33312_28776# _335_.ZN.t27 a_30388_28776# VGND.t6679 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7470 a_63516_18840# a_63428_18884# VGND.t4135 VGND.t2842 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7471 a_48956_1592# a_48868_1636# VGND.t1801 VGND.t1354 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7472 a_66787_30600# a_67117_30600# a_67237_31198# VPWR.t3324 pfet_06v0 ad=0.3456p pd=2.64u as=61.19999f ps=0.7u w=0.36u l=0.5u
X7473 VGND.t947 a_60276_29032# _257_.B VGND.t946 nfet_06v0 ad=0.224p pd=1.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7474 a_43214_21812# a_42778_21812# a_42982_21730# VPWR.t5046 pfet_06v0 ad=61.19999f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X7475 VPWR.t7093 a_14684_2727# a_14596_2824# VPWR.t7092 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7476 a_52876_10567# a_52788_10664# VGND.t3188 VGND.t3187 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7477 a_1020_23544# a_932_23588# VGND.t1802 VGND.t766 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7478 VGND.t2511 _424_.B2 a_52228_19368# VGND.t2510 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7479 VPWR.t661 a_66204_17272# a_66116_17316# VPWR.t660 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7480 a_30912_27508# _350_.A1.t13 _352_.A2.t14 VGND.t6341 nfet_06v0 ad=98.39999f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7481 VPWR.t2538 hold2.I _284_.ZN.t4 VPWR.t2537 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X7482 _428_.Z a_51240_23340# VGND.t430 VGND.t429 nfet_06v0 ad=0.3608p pd=2.52u as=0.218p ps=1.52u w=0.82u l=0.6u
X7483 _223_.ZN _223_.I VGND.t6789 VGND.t6788 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X7484 VPWR.t1454 a_36748_23544# a_36660_23588# VPWR.t1453 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7485 VPWR.t5867 a_50972_1159# a_50884_1256# VPWR.t5866 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7486 a_10428_1159# a_10340_1256# VGND.t4628 VGND.t4627 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7487 VPWR.t7114 a_65308_7431# a_65220_7528# VPWR.t3454 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7488 VGND.t1463 _249_.A2 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I VGND.t1462 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7489 VPWR.t4630 a_15244_27815# a_15156_27912# VPWR.t1165 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7490 VPWR.t2829 vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I VPWR.t2828 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7491 a_44688_26399# a_43736_25896# VPWR.t4110 VPWR.t4109 pfet_06v0 ad=50.4f pd=0.64u as=0.23p ps=1.54u w=0.36u l=0.5u
X7492 a_52292_29480# _268_.A2.t8 a_52068_29480# VPWR.t7065 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7493 VPWR.t5055 a_22860_20408# a_22772_20452# VPWR.t5054 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7494 VPWR.t2911 a_49404_1159# a_49316_1256# VPWR.t2910 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7495 a_35936_19001# a_35504_18955# VPWR.t1329 VPWR.t1328 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X7496 a_41340_2727# a_41252_2824# VGND.t3817 VGND.t3816 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7497 VPWR.t7116 a_38764_16839# a_38676_16936# VPWR.t7115 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7498 a_66316_20408# a_66228_20452# VGND.t4434 VGND.t4433 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7499 VPWR.t5057 a_60492_28248# a_60404_28292# VPWR.t5056 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7500 a_45820_9432# a_45732_9476# VGND.t5116 VGND.t1154 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7501 VPWR.t83 a_34732_19975# a_34644_20072# VPWR.t82 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7502 a_21740_20408# a_21652_20452# VGND.t4441 VGND.t4440 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7503 VGND.t6445 _268_.A1.t9 _274_.A3 VGND.t108 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7504 VPWR.t2929 a_64412_4728# a_64324_4772# VPWR.t2495 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7505 VPWR.t7120 a_60380_2727# a_60292_2824# VPWR.t7119 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7506 a_45148_1592# a_45060_1636# VGND.t4783 VGND.t3517 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7507 _442_.ZN _436_.ZN VGND.t570 VGND.t569 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7508 a_41344_27209# a_39124_27208.t7 a_41099_26841# VGND.t229 nfet_06v0 ad=43.2f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7509 VGND.t5301 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN VGND.t5300 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7510 VPWR.t85 a_31708_19975# a_31620_20072# VPWR.t84 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7511 VGND.t174 a_44784_25987.t6 a_44744_26355# VGND.t173 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X7512 VPWR.t2406 a_5052_9432# a_4964_9476# VPWR.t2405 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7513 VGND.t1672 a_36016_20893# a_35968_20937# VGND.t1671 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X7514 _274_.ZN _268_.A2.t9 a_52964_29480# VPWR.t7066 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7515 VPWR.t7124 a_59820_10567# a_59732_10664# VPWR.t7123 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7516 a_20003_29611# uio_out[5].t13 VGND.t6587 VGND.t6586 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X7517 VPWR.t4524 a_61500_27815# a_61412_27912# VPWR.t4523 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7518 a_31820_25112# a_31732_25156# VGND.t1554 VGND.t1553 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7519 a_23868_2727# a_23780_2824# VGND.t3229 VGND.t3228 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7520 VPWR.t913 a_34172_1592# a_34084_1636# VPWR.t912 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7521 VGND.t4360 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN VGND.t4359 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7522 _335_.ZN.t1 _334_.A1 VPWR.t2349 VPWR.t2348 pfet_06v0 ad=0.2197p pd=1.365u as=0.4056p ps=1.805u w=0.845u l=0.5u
X7523 VGND.t912 a_28256_25597# a_28208_25641# VGND.t911 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X7524 a_67772_12568# a_67684_12612# VGND.t1566 VGND.t1565 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7525 a_39648_19435# _451_.Q.t16 VGND.t6159 VGND.t6158 nfet_06v0 ad=57.59999f pd=0.68u as=0.218p ps=1.52u w=0.36u l=0.6u
X7526 a_31820_21976# a_31732_22020# VGND.t4744 VGND.t4743 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7527 a_20620_25112# a_20532_25156# VGND.t5563 VGND.t5562 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7528 VPWR.t915 a_58140_1592# a_58052_1636# VPWR.t914 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7529 VGND.t6380 _452_.CLK.t59 a_32964_24072.t1 VGND.t6379 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X7530 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN VPWR.t5934 VPWR.t5933 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7531 VGND.t5824 a_61297_30300# _246_.B2 VGND.t71 nfet_06v0 ad=0.2288p pd=1.58u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7532 a_20620_21976# a_20532_22020# VGND.t4750 VGND.t4749 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7533 a_17596_2727# a_17508_2824# VGND.t6005 VGND.t2493 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7534 VPWR.t6244 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t6243 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7535 VGND.t1775 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN VGND.t1774 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7536 a_19744_30301# a_19372_30345# VGND.t1285 VGND.t137 nfet_06v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X7537 _452_.CLK.t28 a_42392_22825.t42 VPWR.t6940 VPWR.t6939 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7538 VGND.t5462 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN VGND.t5461 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7539 a_45372_12568# a_45284_12612# VGND.t5451 VGND.t613 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7540 vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN VPWR.t1102 VPWR.t1101 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7541 VPWR.t4033 a_48060_14136# a_47972_14180# VPWR.t3566 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7542 _473_.Q a_47552_19715# VPWR.t1922 VPWR.t1921 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7543 _455_.D _455_.Q.t15 a_21600_26725# VPWR.t6856 pfet_06v0 ad=0.3159p pd=1.735u as=0.44955p ps=1.955u w=1.215u l=0.5u
X7544 VGND.t512 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I VGND.t511 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7545 a_41432_17801# a_41048_17341# a_40644_17272# VGND.t4864 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7546 _395_.A1 _397_.A2.t20 a_49637_28776# VGND.t6228 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7547 a_58140_11000# a_58052_11044# VGND.t4450 VGND.t4449 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7548 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I VPWR.t4832 VPWR.t4831 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7549 VPWR.t5195 a_48060_11000# a_47972_11044# VPWR.t4169 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7550 VPWR.t87 a_1020_29816# a_932_29860# VPWR.t86 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7551 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I VGND.t2917 VGND.t2916 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7552 VPWR.t5459 a_1020_26680# a_932_26724# VPWR.t2281 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7553 _441_.ZN _441_.A3 a_39780_22805# VGND.t1678 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X7554 a_39480_28776# _402_.A1.t23 _285_.Z VGND.t6441 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7555 a_65756_3160# a_65668_3204# VGND.t4038 VGND.t464 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7556 VPWR.t2554 _349_.A4 a_24952_29032# VPWR.t2553 pfet_06v0 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X7557 VPWR.t720 a_43356_30951# a_43268_31048# VPWR.t719 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7558 a_48508_9432# a_48420_9476# VGND.t5513 VGND.t5512 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7559 a_39873_21236# _438_.A2 a_39669_21236# VGND.t4961 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7560 a_63292_2727# a_63204_2824# VGND.t4046 VGND.t4045 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7561 a_55340_24679# a_55252_24776# VGND.t1330 VGND.t1329 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7562 a_46252_19759# _416_.ZN a_46084_19759# VGND.t1064 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X7563 VPWR.t7130 a_5388_24679# a_5300_24776# VPWR.t7129 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7564 VGND.t6664 _381_.A2.t7 a_50084_24328# VGND.t6663 nfet_06v0 ad=0.104p pd=0.92u as=0.14p ps=1.1u w=0.4u l=0.6u
X7565 VPWR.t1866 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t1865 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7566 VPWR.t2207 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I VPWR.t2206 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7567 a_3708_12568# a_3620_12612# VGND.t3778 VGND.t782 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7568 a_66092_16839# a_66004_16936# VGND.t1826 VGND.t1825 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7569 VPWR.t7132 a_53996_16839# a_53908_16936# VPWR.t7131 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7570 VPWR.t5600 _432_.ZN a_40973_24776# VPWR.t5599 pfet_06v0 ad=0.5346p pd=3.31u as=0.37665p ps=1.835u w=1.215u l=0.5u
X7571 a_67660_13703# a_67572_13800# VGND.t1782 VGND.t1781 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7572 a_51016_25940# _397_.A1.t16 _412_.B2 VGND.t18 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7573 VPWR.t6880 _229_.I.t14 a_63336_29480# VPWR.t6879 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X7574 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN VPWR.t5950 VPWR.t5949 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7575 VPWR.t2347 _334_.A1 _335_.ZN.t0 VPWR.t2346 pfet_06v0 ad=0.4056p pd=1.805u as=0.2197p ps=1.365u w=0.845u l=0.5u
X7576 VGND.t6623 a_42392_22825.t43 _452_.CLK.t29 VGND.t6622 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X7577 a_56460_13703# a_56372_13800# VGND.t2577 VGND.t2576 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7578 VGND.t127 a_49936_19325.t6 a_49896_18909# VGND.t126 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X7579 VPWR.t1006 a_19052_20408# a_18964_20452# VPWR.t1005 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7580 VPWR.t4850 a_40332_21543# a_40244_21640# VPWR.t4849 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7581 a_22972_1592# a_22884_1636# VGND.t3811 VGND.t3810 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7582 a_22748_1159# a_22660_1256# VGND.t357 VGND.t356 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7583 a_14236_1159# a_14148_1256# VGND.t4437 VGND.t4436 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7584 VPWR.t7141 a_63852_10567# a_63764_10664# VPWR.t7140 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7585 a_37644_23544# a_37556_23588# VGND.t3441 VGND.t3440 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7586 a_55004_15271# a_54916_15368# VGND.t5069 VGND.t446 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7587 VPWR.t3634 _346_.A2 a_23284_26724# VPWR.t3633 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7588 a_46940_1592# a_46852_1636# VGND.t4626 VGND.t4625 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7589 VPWR.t1062 a_1020_17272# a_932_17316# VPWR.t1061 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7590 VPWR.t3547 a_51084_13703# a_50996_13800# VPWR.t3546 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7591 VPWR.t1146 a_16700_1592# a_16612_1636# VPWR.t1145 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7592 VPWR.t1125 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN VPWR.t1124 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7593 VPWR.t2998 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN VPWR.t2997 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7594 VPWR.t4720 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_59226_25156# VPWR.t4719 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X7595 VPWR.t515 a_56124_23111# a_56036_23208# VPWR.t514 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7596 a_15244_23544# a_15156_23588# VGND.t5941 VGND.t1249 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7597 a_41776_18504# _331_.ZN a_41572_18504# VPWR.t3724 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7598 _430_.ZN _301_.A1 VGND.t3198 VGND.t3197 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X7599 VPWR.t6003 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I VPWR.t6002 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7600 VPWR.t2320 a_63292_14136# a_63204_14180# VPWR.t2319 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7601 VPWR.t1148 a_45372_15704# a_45284_15748# VPWR.t1147 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7602 VGND.t1139 _290_.ZN uo_out[5].t0 VGND.t1138 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7603 VPWR.t517 a_5388_15271# a_5300_15368# VPWR.t516 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7604 a_28012_21976# a_27924_22020# VGND.t4553 VGND.t4552 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7605 VGND.t4307 _419_.Z a_52136_20936# VGND.t4306 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7606 a_37084_26247# a_36996_26344# VGND.t5999 VGND.t1795 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7607 _386_.A4 _397_.A1.t17 a_46837_29076# VGND.t19 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7608 VPWR.t6348 a_44812_16839# a_44724_16936# VPWR.t3976 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7609 VGND.t2758 a_48888_19243# _474_.Q VGND.t2757 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7610 VPWR.t3856 a_63292_11000# a_63204_11044# VPWR.t3855 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7611 VPWR.t3608 a_52092_14136# a_52004_14180# VPWR.t3607 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7612 VPWR.t3609 a_60268_14136# a_60180_14180# VPWR.t590 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7613 a_48508_14136# a_48420_14180# VGND.t4558 VGND.t4557 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7614 a_63964_18840# a_63876_18884# VGND.t50 VGND.t49 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7615 uo_out[2].t1 _287_.A1.t36 a_36500_29860# VPWR.t6791 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7616 VGND.t6570 _229_.I.t15 _243_.A1 VGND.t6569 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X7617 _365_.ZN _334_.A1 a_35660_27508# VGND.t2238 nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7618 VPWR.t3220 a_29856_29123# a_29848_29535# VPWR.t3219 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X7619 VPWR.t521 a_46044_15271# a_45956_15368# VPWR.t520 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7620 VPWR.t2300 a_52092_11000# a_52004_11044# VPWR.t2299 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7621 a_48508_11000# a_48420_11044# VGND.t4567 VGND.t1814 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7622 _424_.ZN _424_.A1 a_52228_19368# VGND.t303 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7623 VPWR.t7135 a_31088_30301# a_31080_29977# VPWR.t7134 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X7624 VGND.t2445 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7625 VPWR.t5027 a_66652_17272# a_66564_17316# VPWR.t5026 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7626 a_25300_26344# _355_.C.t20 _351_.ZN VPWR.t6681 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7627 VPWR.t4875 a_51532_12135# a_51444_12232# VPWR.t4874 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7628 _441_.ZN _441_.B VPWR.t5255 VPWR.t5254 pfet_06v0 ad=0.4012p pd=1.85u as=0.4972p ps=3.14u w=1.13u l=0.5u
X7629 VPWR.t724 a_64300_13703# a_64212_13800# VPWR.t723 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7630 a_55060_23263# _478_.D a_54192_22851# VPWR.t6069 pfet_06v0 ad=54f pd=0.66u as=0.1872p ps=1.4u w=0.36u l=0.5u
X7631 _324_.C.t0 a_65072_29860# VPWR.t1106 VPWR.t1105 pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X7632 a_28672_31048# _371_.ZN VPWR.t5832 VPWR.t5831 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7633 VPWR.t6351 a_2812_10567# a_2724_10664# VPWR.t3955 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7634 _393_.A1 _383_.ZN VGND.t2545 VGND.t2544 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7635 uo_out[7].t0 a_40038_28720# VPWR.t3139 VPWR.t3138 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7636 a_55228_1159# a_55140_1256# VGND.t2549 VGND.t2548 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7637 _474_.CLK.t31 a_48272_25156.t45 VPWR.t6573 VPWR.t6572 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7638 VPWR.t1904 a_17372_30951# a_17284_31048# VPWR.t1903 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7639 VPWR.t5799 a_3708_18840# a_3620_18884# VPWR.t5798 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7640 VGND.t293 a_44296_24393.t43 clkbuf_1_0__f_clk.I.t18 VGND.t292 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X7641 VPWR.t4755 a_15692_27815# a_15604_27912# VPWR.t2620 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7642 VPWR.t1824 a_29916_1159# a_29828_1256# VPWR.t1823 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7643 a_21852_2727# a_21764_2824# VGND.t3141 VGND.t3140 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7644 uo_out[0].t8 _284_.ZN.t37 VGND.t6249 VGND.t1138 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7645 VGND.t1150 a_8627_30644# a_8627_30644# VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7646 a_20672_30301# a_20379_29977# VPWR.t1947 VPWR.t1946 pfet_06v0 ad=0.2457p pd=1.465u as=0.2619p ps=1.685u w=0.945u l=0.5u
X7647 VPWR.t1971 a_3708_15704# a_3620_15748# VPWR.t1970 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7648 VPWR.t5038 a_33052_17272# a_32964_17316# VPWR.t3696 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7649 a_66764_20408# a_66676_20452# VGND.t4661 VGND.t4660 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7650 VPWR.t1973 a_14796_23544# a_14708_23588# VPWR.t1972 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7651 VPWR.t4757 a_64860_5863# a_64772_5960# VPWR.t2839 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7652 VPWR.t6353 a_40892_2727# a_40804_2824# VPWR.t6352 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7653 VGND.t6223 _459_.CLK.t48 a_29828_24455.t1 VGND.t6222 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X7654 VPWR.t1129 _237_.A1 _238_.I VPWR.t1128 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7655 a_37532_21543# a_37444_21640# VGND.t5583 VGND.t5582 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7656 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN VPWR.t1687 VPWR.t1686 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7657 a_15580_2727# a_15492_2824# VGND.t1273 VGND.t1272 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7658 VGND.t2982 a_40038_28720# uo_out[7].t4 VGND.t2981 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7659 a_29232_29931# a_28820_30344.t6 VPWR.t6368 VPWR.t6367 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X7660 a_19388_1592# a_19300_1636# VGND.t1944 VGND.t1943 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7661 VPWR.t1980 a_14684_1592# a_14596_1636# VPWR.t1484 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7662 a_36204_21327# _317_.A2 VGND.t2450 VGND.t2449 nfet_06v0 ad=58.39999f pd=0.685u as=0.23405p ps=1.555u w=0.365u l=0.6u
X7663 VPWR.t4542 a_33724_21543# a_33636_21640# VPWR.t4541 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7664 a_33164_20408# a_33076_20452# VGND.t4464 VGND.t4463 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7665 VPWR.t6354 a_17036_24679# a_16948_24776# VPWR.t5901 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7666 VPWR.t1984 a_38652_1592# a_38564_1636# VPWR.t1983 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7667 a_18028_28777# _378_.ZN a_17904_28409# VPWR.t3448 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X7668 a_66204_7431# a_66116_7528# VGND.t5990 VGND.t5924 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7669 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I _249_.A2 VGND.t1461 VGND.t1460 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7670 VPWR.t1343 a_65308_9432# a_65220_9476# VPWR.t1342 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7671 VPWR.t7139 a_26108_1159# a_26020_1256# VPWR.t7138 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7672 a_22560_30288# _459_.CLK.t49 VGND.t6225 VGND.t6224 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X7673 a_62060_12135# a_61972_12232# VGND.t4793 VGND.t4792 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7674 _304_.B a_54432_31128# VGND.t4515 VGND.t4514 nfet_06v0 ad=0.1183p pd=0.975u as=0.1183p ps=0.975u w=0.455u l=0.6u
X7675 a_54444_25112# a_54356_25156# VGND.t3108 VGND.t3107 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7676 a_66316_10567# a_66228_10664# VGND.t3231 VGND.t3230 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7677 VGND.t4347 vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I VGND.t4346 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7678 a_30476_23544# a_30388_23588# VGND.t4843 VGND.t4842 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7679 VPWR.t2467 a_15244_26680# a_15156_26724# VPWR.t2466 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7680 VPWR.t6357 a_3260_24679# a_3172_24776# VPWR.t3497 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7681 a_55116_10567# a_55028_10664# VGND.t1197 VGND.t1196 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7682 a_47164_18407# a_47076_18504# VGND.t4371 VGND.t4370 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7683 VPWR.t1349 a_59036_9432# a_58948_9476# VPWR.t1348 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7684 a_27884_25641# _355_.ZN a_27760_25273# VPWR.t2574 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X7685 a_52240_22504# _476_.Q a_52036_22504# VGND.t4158 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X7686 VPWR.t1992 a_41116_1592# a_41028_1636# VPWR.t1991 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7687 _324_.B.t6 _304_.B a_42168_22504# VGND.t4522 nfet_06v0 ad=0.30965p pd=1.685u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7688 VGND.t6495 _287_.A1.t37 uo_out[4].t3 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7689 VPWR.t128 a_49936_19325.t7 a_49896_18909# VPWR.t127 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X7690 a_47259_20127# a_45284_19751.t7 a_46624_19715# VPWR.t7034 pfet_06v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X7691 a_65084_1592# a_64996_1636# VGND.t5188 VGND.t564 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7692 a_44296_24393.t13 clk.t13 VPWR.t6845 VPWR.t6844 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X7693 a_38628_25156# _416_.A1.t15 _444_.D VPWR.t206 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7694 VPWR.t822 a_60380_1592# a_60292_1636# VPWR.t821 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7695 a_26556_1159# a_26468_1256# VGND.t6162 VGND.t6161 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7696 a_18044_1159# a_17956_1256# VGND.t6761 VGND.t6760 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7697 a_30128_27508# _350_.A1.t14 _352_.A2.t12 VGND.t6342 nfet_06v0 ad=98.39999f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7698 VPWR.t2811 a_61276_15271# a_61188_15368# VPWR.t2810 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7699 VGND.t267 clkbuf_1_0__f_clk.I.t58 a_48272_25156.t8 VGND.t266 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X7700 a_52744_26031# a_52400_25987.t7 a_51956_26183# VPWR.t6372 pfet_06v0 ad=0.1791p pd=1.355u as=0.1665p ps=1.285u w=0.36u l=0.5u
X7701 a_41968_17801# a_41432_17801# VGND.t1515 VGND.t1514 nfet_06v0 ad=43.2f pd=0.6u as=0.2637p ps=1.825u w=0.36u l=0.6u
X7702 VPWR.t2782 a_32096_24419# a_32088_24831# VPWR.t2781 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X7703 VPWR.t2311 a_4828_1159# a_4740_1256# VPWR.t2310 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7704 VPWR.t5037 a_66428_12568# a_66340_12612# VPWR.t5036 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7705 VGND.t302 _424_.A1 a_53003_22504# VGND.t301 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7706 VPWR.t3747 a_25100_20408# a_25012_20452# VPWR.t3746 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7707 a_48508_2727# a_48420_2824# VGND.t4125 VGND.t2092 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7708 VPWR.t4445 a_67548_5863# a_67460_5960# VPWR.t4213 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7709 VGND.t4941 a_43824_18147# a_43776_18191# VGND.t4940 nfet_06v0 ad=0.2637p pd=1.825u as=43.2f ps=0.6u w=0.36u l=0.6u
X7710 a_1020_15271# a_932_15368# VGND.t3194 VGND.t3193 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7711 _411_.A2.t4 _470_.Q VPWR.t4221 VPWR.t4220 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X7712 a_33584_22137# a_33152_22091# VPWR.t1468 VPWR.t1467 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X7713 a_4604_25112# a_4516_25156# VGND.t2268 VGND.t2267 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7714 a_2812_19975# a_2724_20072# VGND.t6163 VGND.t3076 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7715 VPWR.t6360 a_67548_2727# a_67460_2824# VPWR.t1175 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7716 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN VGND.t1773 VGND.t1772 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7717 VGND.t6674 _352_.A2.t29 _351_.ZN VGND.t6673 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7718 a_1020_12135# a_932_12232# VGND.t5237 VGND.t4372 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7719 a_4604_21976# a_4516_22020# VGND.t2536 VGND.t2535 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7720 VGND.t2199 a_25652_31048# uio_out[2].t0 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7721 VPWR.t5448 a_62620_18840# a_62532_18884# VPWR.t3859 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7722 VPWR.t1620 a_46198_27060# _330_.A1.t0 VPWR.t1619 pfet_06v0 ad=0.4941p pd=2.03u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7723 VGND.t2228 _316_.A3 _316_.ZN VGND.t2227 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7724 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I VPWR.t2915 VPWR.t2914 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7725 VPWR.t834 a_66876_1592# a_66788_1636# VPWR.t833 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7726 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I VGND.t510 VGND.t509 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7727 a_29848_29535# a_28000_29480# a_29563_29535# VPWR.t1928 pfet_06v0 ad=50.4f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X7728 VPWR.t810 a_62620_15704# a_62532_15748# VPWR.t809 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7729 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN VPWR.t5990 VPWR.t5989 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7730 a_4156_17272# a_4068_17316# VGND.t2195 VGND.t2194 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7731 a_48859_29076# _384_.ZN _392_.A2 VGND.t3022 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7732 a_47776_20893# a_47483_20569# VGND.t2930 VGND.t2929 nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X7733 a_52452_21236# _427_.B1 VGND.t3813 VGND.t3812 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7734 a_41564_24679# a_41476_24776# VGND.t1697 VGND.t1696 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7735 a_30812_17272# a_30724_17316# VGND.t2198 VGND.t1400 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7736 VGND.t6625 a_42392_22825.t44 _452_.CLK.t30 VGND.t6624 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X7737 VPWR.t874 a_3260_15271# a_3172_15368# VPWR.t873 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7738 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN VGND.t604 VGND.t603 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7739 VPWR.t812 a_51420_15704# a_51332_15748# VPWR.t811 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7740 a_62508_23111# a_62420_23208# VGND.t2639 VGND.t2638 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7741 VPWR.t728 _427_.A2 a_52452_24072# VPWR.t727 pfet_06v0 ad=0.40575p pd=2.055u as=0.156p ps=1.12u w=0.6u l=0.5u
X7742 VGND.t5608 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN VGND.t5607 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7743 VPWR.t4270 a_40780_21543# a_40692_21640# VPWR.t4269 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7744 VPWR.t6364 a_24092_24679# a_24004_24776# VPWR.t6363 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7745 a_59036_1159# a_58948_1256# VGND.t5310 VGND.t5309 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7746 a_67548_1159# a_67460_1256# VGND.t2013 VGND.t2012 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7747 VPWR.t4273 a_56572_29383# a_56484_29480# VPWR.t4272 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7748 VPWR.t814 a_7292_1592# a_7204_1636# VPWR.t813 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7749 a_43008_26795# a_42596_27208.t7 VPWR.t144 VPWR.t143 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X7750 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN VGND.t2940 VGND.t2939 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7751 a_55452_15271# a_55364_15368# VGND.t2160 VGND.t2159 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7752 a_53003_22504# _427_.B2 _395_.A3 VGND.t3784 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7753 a_33476_27912# _287_.A1.t38 uo_out[6].t7 VPWR.t6792 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X7754 VPWR.t3278 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN VPWR.t3277 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7755 a_52016_19759# a_51240_19624# VGND.t4417 VGND.t4416 nfet_06v0 ad=43.2f pd=0.6u as=0.142p ps=1.14u w=0.36u l=0.6u
X7756 a_49405_22805# _399_.A1 _399_.ZN VGND.t4076 nfet_06v0 ad=92.99999f pd=1.015u as=0.2015p ps=1.295u w=0.775u l=0.6u
X7757 VPWR.t3901 a_2364_6296# a_2276_6340# VPWR.t3104 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7758 VPWR.t370 a_61500_17272# a_61412_17316# VPWR.t369 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7759 VPWR.t855 a_63068_1592# a_62980_1636# VPWR.t854 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7760 a_35140_26680# _362_.B.t19 a_35756_27216# VGND.t6258 nfet_06v0 ad=0.1672p pd=1.64u as=60.8f ps=0.7u w=0.38u l=0.6u
X7761 VGND.t787 _400_.ZN a_45577_27509# VGND.t786 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X7762 a_4604_15704# a_4516_15748# VGND.t1660 VGND.t1659 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7763 VPWR.t876 a_56572_23111# a_56484_23208# VPWR.t875 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7764 a_33052_15271# a_32964_15368# VGND.t1876 VGND.t1875 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7765 VPWR.t63 a_64748_23111# a_64660_23208# VPWR.t62 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7766 a_15692_23544# a_15604_23588# VGND.t2744 VGND.t2743 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7767 a_36636_25112# a_36548_25156# VGND.t5961 VGND.t5240 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7768 VPWR.t1540 a_2364_3160# a_2276_3204# VPWR.t1539 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7769 a_52428_12135# a_52340_12232# VGND.t4764 VGND.t4763 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7770 VGND.t5 ui_in[2].t1 a_61860_30736# VGND.t4 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X7771 a_48508_10567# a_48420_10664# VGND.t5867 VGND.t5512 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7772 a_28460_21976# a_28372_22020# VGND.t3461 VGND.t3460 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7773 a_36048_24831# a_35616_24776# VPWR.t1666 VPWR.t1665 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X7774 VPWR.t2376 a_18380_21976# a_18292_22020# VPWR.t2375 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7775 VGND.t4521 _304_.B a_42252_20936# VGND.t4520 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7776 a_47388_17272# a_47300_17316# VGND.t2694 VGND.t2693 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7777 a_7516_29383# a_7428_29480# VGND.t5019 VGND.t5018 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7778 a_48956_14136# a_48868_14180# VGND.t3464 VGND.t3463 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7779 a_61612_20408# a_61524_20452# VGND.t544 VGND.t543 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7780 VPWR.t67 a_46492_15271# a_46404_15368# VPWR.t66 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7781 VPWR.t301 _424_.A1 a_51428_20452# VPWR.t300 pfet_06v0 ad=0.4005p pd=2.12u as=0.1456p ps=1.08u w=0.56u l=0.5u
X7782 VGND.t2399 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I VGND.t2398 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7783 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN VPWR.t3680 VPWR.t3679 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7784 VPWR.t6436 a_67436_16839# a_67348_16936# VPWR.t6435 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7785 a_36188_17272# a_36100_17316# VGND.t2043 VGND.t2042 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7786 a_48956_11000# a_48868_11044# VGND.t548 VGND.t547 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7787 VPWR.t3576 _371_.A2 a_28596_27916.t4 VPWR.t3575 pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X7788 VPWR.t6438 a_13340_2727# a_13252_2824# VPWR.t6437 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7789 VPWR.t676 a_51980_12135# a_51892_12232# VPWR.t675 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7790 a_44340_26183# a_44784_25987.t7 a_44736_26031# VGND.t175 nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X7791 a_51308_16839# a_51220_16936# VGND.t504 VGND.t503 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7792 a_52871_31198# a_52415_31220# a_52639_30644# VPWR.t5969 pfet_06v0 ad=61.19999f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X7793 _383_.ZN _381_.Z VGND.t3801 VGND.t3800 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7794 VPWR.t3698 a_56124_28248# a_56036_28292# VPWR.t3456 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7795 a_22560_30288# _459_.CLK.t50 VPWR.t6497 VPWR.t6496 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X7796 VPWR.t4286 a_3708_29383# a_3620_29480# VPWR.t4285 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7797 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN VGND.t4118 VGND.t4117 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7798 _399_.A2 _474_.Q a_48308_23588# VPWR.t4791 pfet_06v0 ad=0.2964p pd=1.66u as=0.3078p ps=1.68u w=1.14u l=0.5u
X7799 a_40108_16839# a_40020_16936# VGND.t1439 VGND.t1438 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7800 a_65308_4295# a_65220_4392# VGND.t671 VGND.t670 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7801 VPWR.t71 a_3708_26247# a_3620_26344# VPWR.t70 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7802 VPWR.t4959 a_38472_30169# _287_.A1.t0 VPWR.t4958 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7803 VGND.t1305 a_11091_30644# a_11091_30644# VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7804 a_64412_18407# a_64324_18504# VGND.t1644 VGND.t1643 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7805 VPWR.t7082 a_3708_23111# a_3620_23208# VPWR.t5196 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7806 a_47700_28292# _470_.Q a_47476_28292# VPWR.t4219 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7807 a_47836_15704# a_47748_15748# VGND.t1445 VGND.t1444 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7808 VPWR.t947 a_26160_27165# a_26152_26841# VPWR.t946 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X7809 VGND.t758 _282_.ZN a_47636_25940# VGND.t757 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7810 a_40684_19368# _451_.Q.t17 _331_.ZN VGND.t6160 nfet_06v0 ad=0.1312p pd=1.14u as=0.2569p ps=1.56u w=0.82u l=0.6u
X7811 a_36636_15704# a_36548_15748# VGND.t1648 VGND.t1647 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7812 VGND.t2980 a_40038_28720# uo_out[7].t3 VGND.t2979 nfet_06v0 ad=0.2911p pd=1.53u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7813 _395_.A3 _427_.B2 VPWR.t3931 VPWR.t3930 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X7814 VPWR.t5810 _272_.B1 a_57220_29861# VPWR.t5809 pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X7815 a_5052_26680# a_4964_26724# VGND.t4753 VGND.t4752 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7816 a_24860_27209# _351_.ZN a_24736_26841# VPWR.t2301 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X7817 _342_.ZN _355_.C.t21 VGND.t6395 VGND.t6394 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7818 VPWR.t6440 a_17484_24679# a_17396_24776# VPWR.t1476 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7819 a_39748_31048# _284_.ZN.t38 uo_out[0].t5 VPWR.t6524 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X7820 VGND.t6397 _355_.C.t22 _454_.D VGND.t6396 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X7821 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I VPWR.t4530 VPWR.t4529 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7822 a_19948_20408# a_19860_20452# VGND.t1727 VGND.t1726 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7823 _470_.D _403_.ZN a_45169_27509# VGND.t3589 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X7824 VPWR.t4366 a_2812_4295# a_2724_4392# VPWR.t3039 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7825 a_40780_27815# a_40692_27912# VGND.t5008 VGND.t5007 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7826 VPWR.t6441 a_65756_7431# a_65668_7528# VPWR.t5819 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7827 a_54892_25112# a_54804_25156# VGND.t2055 VGND.t2054 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7828 VPWR.t77 a_2812_1159# a_2724_1256# VPWR.t76 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7829 a_66764_10567# a_66676_10664# VGND.t5469 VGND.t5468 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7830 VGND.t943 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I VGND.t942 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X7831 a_66988_18407# a_66900_18504# VGND.t2410 VGND.t2409 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7832 a_66204_18840# a_66116_18884# VGND.t1990 VGND.t1989 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7833 VPWR.t4746 a_49852_1159# a_49764_1256# VPWR.t4146 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7834 VPWR.t2286 a_53300_23047# a_52920_22760# VPWR.t2285 pfet_06v0 ad=0.23p pd=1.54u as=0.352p ps=2.48u w=0.8u l=0.5u
X7835 a_17148_29383# a_17060_29480# VGND.t2921 VGND.t2920 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7836 a_55564_10567# a_55476_10664# VGND.t1598 VGND.t1597 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7837 VPWR.t5103 a_21628_1592# a_21540_1636# VPWR.t5102 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7838 a_16252_2727# a_16164_2824# VGND.t5455 VGND.t5454 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7839 VGND.t4453 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].I VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7840 VPWR.t6181 a_64860_4728# a_64772_4772# VPWR.t3116 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7841 a_32592_25227# a_32180_25640.t7 VGND.t33 VGND.t32 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X7842 a_45596_1592# a_45508_1636# VGND.t5652 VGND.t5429 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7843 VPWR.t6445 a_49292_10567# a_49204_10664# VPWR.t6444 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7844 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I VPWR.t4497 VPWR.t4496 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7845 _433_.ZN _226_.ZN a_41664_22020# VPWR.t2377 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7846 a_18828_25112# a_18740_25156# VGND.t5952 VGND.t5951 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7847 a_41160_29083# _495_.I VPWR.t1691 VPWR.t1690 pfet_06v0 ad=0.2542p pd=1.44u as=0.428p ps=2.02u w=0.82u l=0.5u
X7848 VPWR.t1323 _397_.A4 _403_.ZN VPWR.t1322 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X7849 a_39536_23588# _435_.A3 a_39332_23588# VPWR.t972 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7850 VPWR.t6449 a_35292_2727# a_35204_2824# VPWR.t6448 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7851 VPWR.t3071 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN VPWR.t3070 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X7852 a_18828_21976# a_18740_22020# VGND.t598 VGND.t597 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7853 VPWR.t6450 a_46268_10567# a_46180_10664# VPWR.t2464 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7854 VGND.t295 a_44296_24393.t44 clkbuf_1_0__f_clk.I.t17 VGND.t294 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X7855 VPWR.t6093 a_52316_1159# a_52228_1256# VPWR.t6092 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7856 VPWR.t1229 a_66876_12568# a_66788_12612# VPWR.t1228 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7857 _325_.A1.t2 a_42392_19243# VGND.t584 VGND.t583 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7858 a_48384_26724# _474_.CLK.t56 VGND.t6464 VGND.t6463 nfet_06v0 ad=0.2662p pd=2.09u as=0.2662p ps=2.09u w=0.605u l=0.6u
X7859 VPWR.t416 a_17036_23544# a_16948_23588# VPWR.t415 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7860 VPWR.t4108 a_43736_25896# _402_.A1.t0 VPWR.t4107 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7861 a_32240_31048# _223_.I VPWR.t7108 VPWR.t7107 pfet_06v0 ad=0.44955p pd=1.955u as=0.5346p ps=3.31u w=1.215u l=0.5u
X7862 a_58020_27508# _243_.A1 _243_.ZN VGND.t5787 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7863 a_36524_16839# a_36436_16936# VGND.t3574 VGND.t3573 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7864 a_41948_17433# a_41432_17801# VPWR.t1598 VPWR.t1597 pfet_06v0 ad=43.2f pd=0.6u as=0.1044p ps=0.94u w=0.36u l=0.5u
X7865 a_30240_24776# a_29828_24455.t7 VPWR.t6389 VPWR.t6388 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X7866 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN VPWR.t5625 VPWR.t5624 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7867 _370_.ZN _352_.A2.t30 a_29575_28293# VPWR.t6995 pfet_06v0 ad=0.3159p pd=1.735u as=0.37665p ps=1.835u w=1.215u l=0.5u
X7868 a_37084_26680# a_36996_26724# VGND.t386 VGND.t385 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7869 a_64412_3160# a_64324_3204# VGND.t5885 VGND.t4548 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7870 uo_out[4].t2 _287_.A1.t39 VGND.t6496 VGND.t146 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X7871 VPWR.t2236 a_46044_1159# a_45956_1256# VPWR.t2235 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7872 VPWR.t5482 a_59372_12135# a_59284_12232# VPWR.t5481 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7873 a_33776_29123# a_33483_29535# VPWR.t3530 VPWR.t3529 pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
X7874 a_61029_31220# a_60909_30600# a_60285_30600# VPWR.t1436 pfet_06v0 ad=61.19999f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X7875 a_48272_25156.t0 clkbuf_1_0__f_clk.I.t59 VPWR.t274 VPWR.t273 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X7876 a_50300_15271# a_50212_15368# VGND.t374 VGND.t373 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7877 VPWR.t422 a_3260_23544# a_3172_23588# VPWR.t421 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7878 a_6172_30951# a_6084_31048# VGND.t4176 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7879 a_54780_26247# a_54692_26344# VGND.t4421 VGND.t4420 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7880 a_33276_1159# a_33188_1256# VGND.t5484 VGND.t5483 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7881 a_41788_1159# a_41700_1256# VGND.t4583 VGND.t4582 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7882 a_51868_15704# a_51780_15748# VGND.t5522 VGND.t5521 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7883 _335_.ZN.t19 _459_.Q.t17 VPWR.t6978 VPWR.t6977 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X7884 VPWR.t7118 a_40220_26247# a_40132_26344# VPWR.t7117 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7885 a_30388_28776# _371_.A1.t19 _350_.A2.t15 VGND.t6236 nfet_06v0 ad=0.2132p pd=1.34u as=0.30965p ps=1.685u w=0.82u l=0.6u
X7886 a_34532_27208# _362_.B.t20 a_34348_27208# VGND.t6259 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7887 VPWR.t6452 a_62172_18407# a_62084_18504# VPWR.t4621 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7888 a_62956_23111# a_62868_23208# VGND.t3651 VGND.t3650 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7889 a_45260_17272# a_45172_17316# VGND.t5174 VGND.t5173 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7890 a_30036_25940# _352_.A2.t31 VGND.t6676 VGND.t6675 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7891 _223_.I a_31088_30301# VGND.t6811 VGND.t71 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7892 VPWR.t6454 a_48508_18407# a_48420_18504# VPWR.t6453 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7893 a_1916_9432# a_1828_9476# VGND.t3340 VGND.t3339 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7894 _304_.ZN.t7 _304_.A1.t17 a_42728_20452# VPWR.t6611 pfet_06v0 ad=0.2847p pd=1.615u as=0.33945p ps=1.715u w=1.095u l=0.5u
X7895 _441_.B _430_.ZN VPWR.t4820 VPWR.t4819 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X7896 a_32380_26247# a_32292_26344# VGND.t5996 VGND.t5995 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7897 VPWR.t7122 a_52540_15271# a_52452_15368# VPWR.t7121 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7898 a_18716_26247# a_18628_26344# VGND.t5998 VGND.t5997 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7899 a_37408_18504# a_36996_18183.t7 VPWR.t6944 VPWR.t6943 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X7900 a_1916_6296# a_1828_6340# VGND.t734 VGND.t0 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7901 a_48060_12568# a_47972_12612# VGND.t3949 VGND.t3571 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7902 VPWR.t2135 a_36432_19325# a_36404_19001# VPWR.t2134 pfet_06v0 ad=0.1044p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X7903 a_61029_30644# a_60909_30600# a_60285_30600# VGND.t45 nfet_06v0 ad=43.2f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X7904 VGND.t5045 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN VGND.t5044 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7905 a_32380_23111# a_32292_23208# VGND.t1856 VGND.t1855 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7906 VPWR.t4741 a_67548_4728# a_67460_4772# VPWR.t3377 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7907 VGND.t5591 a_38816_27555# a_38768_27599# VGND.t5590 nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X7908 VPWR.t5489 _395_.A3 a_50732_23233# VPWR.t5488 pfet_06v0 ad=0.5913p pd=3.27u as=0.2847p ps=1.615u w=1.095u l=0.5u
X7909 a_33024_25273# a_32592_25227# VPWR.t5912 VPWR.t5911 pfet_06v0 ad=54f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X7910 a_18716_23111# a_18628_23208# VGND.t5099 VGND.t5098 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7911 _452_.CLK.t31 a_42392_22825.t45 VGND.t6627 VGND.t6626 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X7912 a_1020_28248# a_932_28292# VGND.t687 VGND.t686 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7913 VPWR.t5343 a_52848_25987# a_52744_26031# VPWR.t5342 pfet_06v0 ad=0.1044p pd=0.94u as=0.1791p ps=1.355u w=0.36u l=0.5u
X7914 _268_.A2.t1 a_50436_30689# VGND.t2011 VGND.t2010 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X7915 _386_.ZN _386_.A4 VGND.t643 VGND.t642 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X7916 a_46576_19759# a_45696_20072# a_46252_19759# VGND.t2469 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X7917 _340_.A2 _350_.A1.t15 VPWR.t6628 VPWR.t6627 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X7918 a_52876_12135# a_52788_12232# VGND.t4379 VGND.t4378 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7919 a_4940_26247# a_4852_26344# VGND.t1903 VGND.t1902 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7920 VPWR.t4597 a_19164_21543# a_19076_21640# VPWR.t4596 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7921 _373_.ZN _355_.C.t23 VGND.t6399 VGND.t6398 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X7922 VPWR.t7061 a_45456_30301.t6 a_45416_29885# VPWR.t7060 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X7923 a_49652_20936# _473_.Q a_49448_20936# VGND.t4991 nfet_06v0 ad=88.2f pd=0.84u as=88.2f ps=0.84u w=0.42u l=0.6u
X7924 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I VGND.t5164 VGND.t5163 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7925 a_4940_23111# a_4852_23208# VGND.t3137 VGND.t3136 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7926 VPWR.t7128 a_46044_30951# a_45956_31048# VPWR.t7127 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7927 a_1916_26247# a_1828_26344# VGND.t3000 VGND.t1316 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7928 a_29232_29931# a_28820_30344.t7 VGND.t6095 VGND.t139 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X7929 a_7964_29383# a_7876_29480# VGND.t4322 VGND.t4321 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7930 a_59172_27912# _252_.B _247_.ZN VPWR.t788 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X7931 a_30520_27508# _350_.A2.t29 VGND.t6299 VGND.t6298 nfet_06v0 ad=98.39999f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X7932 uio_out[7].t0 a_18096_27165# VPWR.t400 VPWR.t399 pfet_06v0 ad=0.4392p pd=1.94u as=0.38575p ps=1.92u w=1.22u l=0.5u
X7933 a_1916_23111# a_1828_23208# VGND.t4186 VGND.t4185 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7934 a_25420_30345# _342_.ZN a_25296_29977# VPWR.t4296 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X7935 VPWR.t6457 a_67884_16839# a_67796_16936# VPWR.t6456 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7936 a_20496_26344# a_20084_26023.t7 VPWR.t7007 VPWR.t7006 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X7937 VPWR.t6499 _459_.CLK.t51 a_41028_28776.t0 VPWR.t6498 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X7938 _238_.I _237_.A1 a_58709_29076# VGND.t1076 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7939 a_51756_16839# a_51668_16936# VGND.t2566 VGND.t2565 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7940 VPWR.t718 a_32268_23544# a_32180_23588# VPWR.t717 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7941 _474_.D _424_.B1.t15 a_50196_21640# VPWR.t6620 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X7942 VPWR.t5928 _285_.Z a_37386_31048# VPWR.t5927 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X7943 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN VPWR.t842 VPWR.t841 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7944 a_55004_21543# a_54916_21640# VGND.t5002 VGND.t5001 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7945 _327_.A2 a_44752_18147# VGND.t4017 VGND.t4016 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7946 VPWR.t642 a_2364_21543# a_2276_21640# VPWR.t641 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7947 a_40556_16839# a_40468_16936# VGND.t1964 VGND.t1963 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7948 VPWR.t722 a_21068_23544# a_20980_23588# VPWR.t721 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7949 VPWR.t6459 a_20508_24679# a_20420_24776# VPWR.t6458 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7950 a_51414_22504# _475_.Q a_51220_22504# VGND.t4854 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X7951 _335_.ZN.t8 _460_.Q VPWR.t3469 VPWR.t3468 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X7952 a_64860_18407# a_64772_18504# VGND.t2146 VGND.t1762 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7953 VPWR.t4335 a_58140_26680# a_58052_26724# VPWR.t4334 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7954 a_46476_20937# _475_.D a_46352_20569# VPWR.t2077 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X7955 a_41012_23208# _438_.ZN VPWR.t2649 VPWR.t2648 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7956 _371_.A1.t3 _334_.A1 a_33940_27208# VGND.t2237 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7957 _350_.A1.t0 a_29856_29123# VPWR.t3218 VPWR.t3217 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7958 a_1020_18840# a_932_18884# VGND.t623 VGND.t622 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7959 _409_.ZN _407_.A1 a_50276_27912# VPWR.t522 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X7960 a_41536_17636# a_41048_17341# a_41968_17801# VGND.t4863 nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X7961 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN VGND.t1650 VGND.t1649 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7962 a_61612_10567# a_61524_10664# VGND.t2123 VGND.t2122 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7963 _441_.B _439_.ZN VPWR.t6108 VPWR.t6107 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X7964 VGND.t886 _395_.A1 _383_.ZN VGND.t885 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X7965 a_52436_18884# _424_.B2 VPWR.t2647 VPWR.t2646 pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X7966 VGND.t6351 _230_.I.t15 _243_.B2 VGND.t6350 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X7967 a_4940_16839# a_4852_16936# VGND.t2716 VGND.t2715 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7968 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I VGND.t3314 VGND.t3313 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X7969 _316_.A3 _311_.Z VGND.t4324 VGND.t4323 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X7970 a_1916_16839# a_1828_16936# VGND.t2822 VGND.t1937 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7971 a_31260_18407# a_31172_18504# VGND.t2823 VGND.t1939 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7972 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN VPWR.t5693 VPWR.t5692 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X7973 VGND.t2414 hold2.I a_42376_25640# VGND.t2413 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7974 VPWR.t6433 a_2812_19975# a_2724_20072# VPWR.t4260 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7975 a_18044_1592# a_17956_1636# VGND.t1129 VGND.t1128 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7976 VPWR.t7068 a_58700_16839# a_58612_16936# VPWR.t7067 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7977 a_63292_12568# a_63204_12612# VGND.t2348 VGND.t2347 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7978 VPWR.t513 a_13340_1592# a_13252_1636# VPWR.t512 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7979 VGND.t241 _304_.ZN.t17 a_42376_22504# VGND.t240 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X7980 VPWR.t3649 a_3708_28248# a_3620_28292# VPWR.t3428 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7981 VPWR.t7070 a_47500_16839# a_47412_16936# VPWR.t7069 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7982 a_52092_12568# a_52004_12612# VGND.t488 VGND.t487 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7983 a_66652_18840# a_66564_18884# VGND.t630 VGND.t629 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7984 a_37964_18191# _330_.ZN a_37840_18559# VPWR.t6310 pfet_06v0 ad=0.1872p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X7985 a_22748_23111# a_22660_23208# VGND.t3908 VGND.t3907 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7986 VPWR.t1140 a_3708_25112# a_3620_25156# VPWR.t1139 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7987 VGND.t6743 a_45456_30301.t7 a_46828_30345# VGND.t137 nfet_06v0 ad=0.1584p pd=1.6u as=43.2f ps=0.6u w=0.36u l=0.6u
X7988 VPWR.t5364 a_20060_1159# a_19972_1256# VPWR.t5363 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7989 VPWR.t1090 a_65420_12135# a_65332_12232# VPWR.t1089 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7990 VPWR.t7142 a_31708_15271# a_31620_15368# VPWR.t1495 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7991 a_37084_1159# a_36996_1256# VGND.t837 VGND.t836 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7992 a_45596_1159# a_45508_1256# VGND.t6754 VGND.t6753 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7993 VPWR.t55 a_2364_12135# a_2276_12232# VPWR.t54 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7994 VPWR.t4718 a_34396_21543# a_34308_21640# VPWR.t4717 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7995 VPWR.t6345 a_3708_8999# a_3620_9096# VPWR.t3406 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7996 _454_.D _345_.A2 VGND.t3071 VGND.t3070 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X7997 VPWR.t61 a_54220_12135# a_54132_12232# VPWR.t60 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X7998 a_33940_27208# _362_.B.t21 a_33764_27208# VGND.t6260 nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X7999 a_50524_30345# _409_.ZN a_49600_30180# VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X8000 a_42340_28409# a_41028_28776.t7 a_41996_28777# VPWR.t7099 pfet_06v0 ad=43.2f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X8001 a_60940_15704# a_60852_15748# VGND.t5625 VGND.t5624 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8002 VPWR.t4728 a_23196_21543# a_23108_21640# VPWR.t4727 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X8003 _435_.ZN _438_.A2 a_39760_23588# VPWR.t5116 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X8004 VPWR.t4729 a_13788_29383# a_13700_29480# VPWR.t3785 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X8005 VPWR.t1714 a_32828_1159# a_32740_1256# VPWR.t1702 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X8006 VPWR.t519 a_19836_1592# a_19748_1636# VPWR.t518 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X8007 a_33052_18840# a_32964_18884# VGND.t4554 VGND.t3353 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8008 VGND.t297 a_44296_24393.t45 clkbuf_1_0__f_clk.I.t16 VGND.t296 nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X8009 a_51620_19911# a_52064_19715.t7 a_52016_19759# VGND nfet_06v0 ad=93.59999f pd=0.88u as=43.2f ps=0.6u w=0.36u l=0.6u
X8010 VGND.t4519 _304_.B a_41264_30669# VGND.t4150 nfet_06v0 ad=0.218p pd=1.52u as=57.59999f ps=0.68u w=0.36u l=0.6u
X8011 VPWR.t4005 a_22352_25987# a_22344_26399# VPWR.t4004 pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X8012 a_1020_30951# a_932_31048# VGND.t4079 VGND.t34 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8013 VPWR.t882 a_26556_27815# a_26468_27912# VPWR.t881 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X8014 VPWR.t6350 a_24988_23111# a_24900_23208# VPWR.t6349 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X8015 a_66652_7431# a_66564_7528# VGND.t2595 VGND.t2594 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8016 a_36972_16839# a_36884_16936# VGND.t2186 VGND.t2185 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X8017 VPWR.t1902 a_17484_23544# a_17396_23588# VPWR.t1901 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X8018 a_58020_27508# _243_.B2 VGND.t5289 VGND.t5288 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8019 VPWR.t990 a_65756_9432# a_65668_9476# VPWR.t989 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X8020 a_28256_25597# a_27884_25641# VPWR.t2967 VPWR.t2966 pfet_06v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X8021 VPWR.t6432 a_26556_1159# a_26468_1256# VPWR.t6431 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X8022 a_43600_25640# hold2.I VGND.t2412 VGND.t2411 nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X8023 a_46336_30345# a_45800_30345# VGND.t5092 VGND.t137 nfet_06v0 ad=43.2f pd=0.6u as=0.2637p ps=1.825u w=0.36u l=0.6u
X8024 a_47412_23588# _397_.A2.t21 a_47172_23588# VPWR.t6507 pfet_06v0 ad=0.1736p pd=1.18u as=0.196p ps=1.26u w=0.56u l=0.5u
R0 VPWR.t3355 VPWR.t4669 988.418
R1 VPWR.n392 VPWR.t1113 986.607
R2 VPWR.t5565 VPWR.t6941 968.213
R3 VPWR.t6748 VPWR.t4137 947.876
R4 VPWR.t3324 VPWR.t3323 880.309
R5 VPWR.t1436 VPWR.t358 880.309
R6 VPWR.t5521 VPWR.t3241 880.309
R7 VPWR.t5969 VPWR.t5454 880.309
R8 VPWR.t1163 VPWR.t2760 864.865
R9 VPWR.t4153 VPWR.t2584 864.865
R10 VPWR.t1659 VPWR.t6199 864.865
R11 VPWR.t5350 VPWR.t545 864.865
R12 VPWR.t847 VPWR.t5350 864.865
R13 VPWR.t1312 VPWR.t847 864.865
R14 VPWR.t2081 VPWR.t2293 864.865
R15 VPWR.t2293 VPWR.t3107 864.865
R16 VPWR.t3107 VPWR.t1903 864.865
R17 VPWR.t543 VPWR.t1840 864.865
R18 VPWR.t1407 VPWR.t2445 864.865
R19 VPWR.t1131 VPWR.t3940 864.865
R20 VPWR.t1028 VPWR.t1704 864.865
R21 VPWR.t3765 VPWR.t4342 864.865
R22 VPWR.t858 VPWR.t3765 864.865
R23 VPWR.t5634 VPWR.t858 864.865
R24 VPWR.t6116 VPWR.t5400 864.865
R25 VPWR.t5400 VPWR.t350 864.865
R26 VPWR.t350 VPWR.t2289 864.865
R27 VPWR.t2289 VPWR.t4892 864.865
R28 VPWR.t4892 VPWR.t653 864.865
R29 VPWR.t653 VPWR.t2834 864.865
R30 VPWR.t2834 VPWR.t4242 864.865
R31 VPWR.t1151 VPWR.t3064 864.865
R32 VPWR.t3064 VPWR.t2968 864.865
R33 VPWR.t2968 VPWR.t5529 864.865
R34 VPWR.t5529 VPWR.t5429 864.865
R35 VPWR.t5429 VPWR.t5297 864.865
R36 VPWR.t5297 VPWR.t1952 864.865
R37 VPWR.t1952 VPWR.t5548 864.865
R38 VPWR.t622 VPWR.t7127 864.865
R39 VPWR.t4283 VPWR.t622 864.865
R40 VPWR.t3281 VPWR.t4283 864.865
R41 VPWR.t5980 VPWR.t3281 864.865
R42 VPWR.t5917 VPWR.t5980 864.865
R43 VPWR.t719 VPWR.t5917 864.865
R44 VPWR.t5494 VPWR.t719 864.865
R45 VPWR.t2855 VPWR.t691 864.865
R46 VPWR.t4406 VPWR.t2855 864.865
R47 VPWR.t1577 VPWR.t4406 864.865
R48 VPWR.t3793 VPWR.t1577 864.865
R49 VPWR.t5082 VPWR.t3793 864.865
R50 VPWR.t5580 VPWR.t5082 864.865
R51 VPWR.t5811 VPWR.t5580 864.865
R52 VPWR.t551 VPWR.t4376 864.865
R53 VPWR.t1348 VPWR.t551 864.865
R54 VPWR.t2087 VPWR.t1348 864.865
R55 VPWR.t4859 VPWR.t2087 864.865
R56 VPWR.t1545 VPWR.t4859 864.865
R57 VPWR.t446 VPWR.t1545 864.865
R58 VPWR.t3521 VPWR.t446 864.865
R59 VPWR.t4077 VPWR.t1093 864.865
R60 VPWR.t4975 VPWR.t4077 864.865
R61 VPWR.t5374 VPWR.t4975 864.865
R62 VPWR.t5786 VPWR.t5374 864.865
R63 VPWR.t6121 VPWR.t5786 864.865
R64 VPWR.t1497 VPWR.t6121 864.865
R65 VPWR.t3938 VPWR.t1497 864.865
R66 VPWR.t5065 VPWR.t1938 864.865
R67 VPWR.t5648 VPWR.t5065 864.865
R68 VPWR.t1802 VPWR.t5648 864.865
R69 VPWR.t3293 VPWR.t1802 864.865
R70 VPWR.t6236 VPWR.t3293 864.865
R71 VPWR.t6272 VPWR.t6236 864.865
R72 VPWR.t4363 VPWR.t6272 864.865
R73 VPWR.t2459 VPWR.t5714 864.865
R74 VPWR.t5838 VPWR.t2459 864.865
R75 VPWR.t5279 VPWR.t5838 864.865
R76 VPWR.t2692 VPWR.t5279 864.865
R77 VPWR.t6050 VPWR.t2692 864.865
R78 VPWR.t5285 VPWR.t6050 864.865
R79 VPWR.t1829 VPWR.t5285 864.865
R80 VPWR.t6299 VPWR.t566 864.865
R81 VPWR.t4516 VPWR.t6299 864.865
R82 VPWR.t3244 VPWR.t4516 864.865
R83 VPWR.t3685 VPWR.t3244 864.865
R84 VPWR.t6234 VPWR.t3685 864.865
R85 VPWR.t5947 VPWR.t6234 864.865
R86 VPWR.t3740 VPWR.t5947 864.865
R87 VPWR.t3746 VPWR.t1499 864.865
R88 VPWR.t1892 VPWR.t3746 864.865
R89 VPWR.t3844 VPWR.t1892 864.865
R90 VPWR.t5372 VPWR.t3844 864.865
R91 VPWR.t6182 VPWR.t5372 864.865
R92 VPWR.t5054 VPWR.t6182 864.865
R93 VPWR.t1024 VPWR.t5054 864.865
R94 VPWR.t1808 VPWR.t4586 864.865
R95 VPWR.t2883 VPWR.t1808 864.865
R96 VPWR.t1073 VPWR.t2883 864.865
R97 VPWR.t1817 VPWR.t1073 864.865
R98 VPWR.t2469 VPWR.t1817 864.865
R99 VPWR.t1005 VPWR.t2469 864.865
R100 VPWR.t864 VPWR.t1005 864.865
R101 VPWR.t3687 VPWR.t3527 864.865
R102 VPWR.t2129 VPWR.t3687 864.865
R103 VPWR.t4338 VPWR.t2129 864.865
R104 VPWR.t2308 VPWR.t4338 864.865
R105 VPWR.t4276 VPWR.t2308 864.865
R106 VPWR.t1087 VPWR.t4276 864.865
R107 VPWR.t3926 VPWR.t1087 864.865
R108 VPWR.t2974 VPWR.t4197 864.865
R109 VPWR.t4197 VPWR.t2667 864.865
R110 VPWR.t2667 VPWR.t64 864.865
R111 VPWR.t64 VPWR.t3383 864.865
R112 VPWR.t4952 VPWR.t987 864.865
R113 VPWR.t7119 VPWR.t4952 864.865
R114 VPWR.t4623 VPWR.t7119 864.865
R115 VPWR.t5859 VPWR.t4623 864.865
R116 VPWR.t1439 VPWR.t5859 864.865
R117 VPWR.t625 VPWR.t1439 864.865
R118 VPWR.t867 VPWR.t625 864.865
R119 VPWR.t1308 VPWR.t4372 864.865
R120 VPWR.t1239 VPWR.t1308 864.865
R121 VPWR.t4452 VPWR.t1239 864.865
R122 VPWR.t2927 VPWR.t4452 864.865
R123 VPWR.t5198 VPWR.t2927 864.865
R124 VPWR.t452 VPWR.t5198 864.865
R125 VPWR.t5170 VPWR.t452 864.865
R126 VPWR.t4657 VPWR.t3738 864.865
R127 VPWR.t3738 VPWR.t5893 864.865
R128 VPWR.t5893 VPWR.t2696 864.865
R129 VPWR.t2696 VPWR.t1038 864.865
R130 VPWR.t1038 VPWR.t2934 864.865
R131 VPWR.t2934 VPWR.t2748 864.865
R132 VPWR.t2748 VPWR.t6322 864.865
R133 VPWR.t6013 VPWR.t1962 864.865
R134 VPWR.t1962 VPWR.t1571 864.865
R135 VPWR.t1571 VPWR.t4288 864.865
R136 VPWR.t4288 VPWR.t3319 864.865
R137 VPWR.t3319 VPWR.t5690 864.865
R138 VPWR.t5690 VPWR.t5853 864.865
R139 VPWR.t5853 VPWR.t5129 864.865
R140 VPWR.t1116 VPWR.t639 864.865
R141 VPWR.t1015 VPWR.t1116 864.865
R142 VPWR.t500 VPWR.t1015 864.865
R143 VPWR.t3132 VPWR.t500 864.865
R144 VPWR.t825 VPWR.t3132 864.865
R145 VPWR.t5577 VPWR.t825 864.865
R146 VPWR.t4788 VPWR.t5577 864.865
R147 VPWR.t860 VPWR.t318 864.865
R148 VPWR.t3160 VPWR.t860 864.865
R149 VPWR.t6352 VPWR.t3160 864.865
R150 VPWR.t2808 VPWR.t6352 864.865
R151 VPWR.t3554 VPWR.t2808 864.865
R152 VPWR.t1137 VPWR.t3554 864.865
R153 VPWR.t1775 VPWR.t1137 864.865
R154 VPWR.t2083 VPWR.t2803 864.865
R155 VPWR.t2803 VPWR.t831 864.865
R156 VPWR.t831 VPWR.t4028 864.865
R157 VPWR.t4028 VPWR.t4896 864.865
R158 VPWR.t4896 VPWR.t725 864.865
R159 VPWR.t725 VPWR.t2101 864.865
R160 VPWR.t2101 VPWR.t6448 864.865
R161 VPWR.t4810 VPWR.t2816 864.865
R162 VPWR.t2816 VPWR.t3811 864.865
R163 VPWR.t3811 VPWR.t748 864.865
R164 VPWR.t748 VPWR.t2005 864.865
R165 VPWR.t2005 VPWR.t379 864.865
R166 VPWR.t379 VPWR.t3486 864.865
R167 VPWR.t3486 VPWR.t4535 864.865
R168 VPWR.t3327 VPWR.t2333 864.865
R169 VPWR.t2265 VPWR.t3327 864.865
R170 VPWR.t3275 VPWR.t2265 864.865
R171 VPWR.t596 VPWR.t3275 864.865
R172 VPWR.t4344 VPWR.t596 864.865
R173 VPWR.t5792 VPWR.t4344 864.865
R174 VPWR.t2154 VPWR.t5792 864.865
R175 VPWR.t6222 VPWR.t4946 864.865
R176 VPWR.t2688 VPWR.t6222 864.865
R177 VPWR.t3758 VPWR.t2688 864.865
R178 VPWR.t5734 VPWR.t3758 864.865
R179 VPWR.t2567 VPWR.t5734 864.865
R180 VPWR.t3438 VPWR.t2567 864.865
R181 VPWR.t3375 VPWR.t3438 864.865
R182 VPWR.t3681 VPWR.t784 864.865
R183 VPWR.t784 VPWR.t3503 864.865
R184 VPWR.t3503 VPWR.t4240 864.865
R185 VPWR.t4240 VPWR.t3866 864.865
R186 VPWR.t3866 VPWR.t7090 864.865
R187 VPWR.t7090 VPWR.t2970 864.865
R188 VPWR.t2970 VPWR.t3699 864.865
R189 VPWR.t3605 VPWR.t6118 864.865
R190 VPWR.t5266 VPWR.t3605 864.865
R191 VPWR.t5388 VPWR.t5266 864.865
R192 VPWR.t3778 VPWR.t5388 864.865
R193 VPWR.t1198 VPWR.t3778 864.865
R194 VPWR.t74 VPWR.t1198 864.865
R195 VPWR.t5650 VPWR.t74 864.865
R196 VPWR.t3134 VPWR.t5517 864.865
R197 VPWR.t7092 VPWR.t3134 864.865
R198 VPWR.t2976 VPWR.t7092 864.865
R199 VPWR.t560 VPWR.t2976 864.865
R200 VPWR.t6437 VPWR.t560 864.865
R201 VPWR.t916 VPWR.t6437 864.865
R202 VPWR.t2423 VPWR.t916 864.865
R203 VPWR.t1821 VPWR.t954 864.865
R204 VPWR.t5378 VPWR.t1821 864.865
R205 VPWR.t2987 VPWR.t5378 864.865
R206 VPWR.t856 VPWR.t2987 864.865
R207 VPWR.t1434 VPWR.t856 864.865
R208 VPWR.t4776 VPWR.t1434 864.865
R209 VPWR.t1091 VPWR.t4776 864.865
R210 VPWR.t5501 VPWR.t6184 864.865
R211 VPWR.t6184 VPWR.t2630 864.865
R212 VPWR.t2630 VPWR.t4732 864.865
R213 VPWR.t4732 VPWR.t5863 864.865
R214 VPWR.t6622 VPWR.t6627 859.073
R215 VPWR.t340 VPWR.t2921 837.838
R216 VPWR.t2590 VPWR 789.576
R217 VPWR.n1522 VPWR.t3660 745.174
R218 VPWR.n1535 VPWR.t1220 743.244
R219 VPWR.n1572 VPWR.t6899 725.87
R220 VPWR.n946 VPWR.t6772 709.163
R221 VPWR.n928 VPWR.t6329 709.163
R222 VPWR.n114 VPWR.t2750 709.163
R223 VPWR.n1782 VPWR.t1537 709.163
R224 VPWR.n2879 VPWR.t5703 709.163
R225 VPWR.t4886 VPWR.n2955 707.163
R226 VPWR.t5863 VPWR.n3685 707.163
R227 VPWR.n1525 VPWR.t2580 706.564
R228 VPWR.n141 VPWR.t4040 705.179
R229 VPWR.n2880 VPWR.t685 705.179
R230 VPWR.n175 VPWR.t4541 705.179
R231 VPWR.n2952 VPWR.t82 705.179
R232 VPWR.n1059 VPWR.t1739 694.981
R233 VPWR.t1206 VPWR 662.163
R234 VPWR VPWR.t4312 662.163
R235 VPWR.t778 VPWR.n1525 648.649
R236 VPWR.n1542 VPWR.t6116 648.649
R237 VPWR.t5283 VPWR.n1059 648.649
R238 VPWR.n1022 VPWR.t1151 648.649
R239 VPWR.t7127 VPWR.n1507 648.649
R240 VPWR.t4376 VPWR.n2327 648.649
R241 VPWR.t1093 VPWR.n2328 648.649
R242 VPWR.t1938 VPWR.n2329 648.649
R243 VPWR.t5714 VPWR.n2330 648.649
R244 VPWR.t566 VPWR.n2956 648.649
R245 VPWR.t1499 VPWR.n2957 648.649
R246 VPWR.t4586 VPWR.n2958 648.649
R247 VPWR.t3527 VPWR.n2959 648.649
R248 VPWR.t987 VPWR.n2480 648.649
R249 VPWR.t4372 VPWR.n2481 648.649
R250 VPWR.n2482 VPWR.t4657 648.649
R251 VPWR.n257 VPWR.t6013 648.649
R252 VPWR.t639 VPWR.n2620 648.649
R253 VPWR.t318 VPWR.n2621 648.649
R254 VPWR.n2623 VPWR.t2083 648.649
R255 VPWR.n2622 VPWR.t4810 648.649
R256 VPWR.t2333 VPWR.n5 648.649
R257 VPWR.t4946 VPWR.n6 648.649
R258 VPWR.n39 VPWR.t3681 648.649
R259 VPWR.t6118 VPWR.n57 648.649
R260 VPWR.t5517 VPWR.n58 648.649
R261 VPWR.t954 VPWR.n59 648.649
R262 VPWR.n3686 VPWR.t5501 648.649
R263 VPWR.t2360 VPWR 642.857
R264 VPWR.t6771 VPWR 642.857
R265 VPWR VPWR.t7021 642.857
R266 VPWR.t1379 VPWR.t3325 637.067
R267 VPWR.t359 VPWR.t340 637.067
R268 VPWR.t2921 VPWR.t5519 637.067
R269 VPWR.t4137 VPWR.t5970 637.067
R270 VPWR.t5386 VPWR 623.553
R271 VPWR VPWR.t2770 623.553
R272 VPWR VPWR.t1381 610.039
R273 VPWR VPWR.t320 610.039
R274 VPWR VPWR.t2291 610.039
R275 VPWR VPWR.t7107 604.247
R276 VPWR VPWR.t6621 592.664
R277 VPWR VPWR.t6972 592.664
R278 VPWR.t6141 VPWR 592.664
R279 VPWR VPWR.t2113 592.664
R280 VPWR.t2529 VPWR 577.221
R281 VPWR.t5652 VPWR 577.221
R282 VPWR VPWR.t2306 573.36
R283 VPWR VPWR.t2148 573.36
R284 VPWR VPWR.t5303 573.36
R285 VPWR VPWR.t5872 573.36
R286 VPWR VPWR.t4123 573.36
R287 VPWR.t2760 VPWR 565.638
R288 VPWR.t2287 VPWR 565.638
R289 VPWR.t1232 VPWR 565.638
R290 VPWR.t2584 VPWR 565.638
R291 VPWR.t6199 VPWR 565.638
R292 VPWR.t5317 VPWR 565.638
R293 VPWR.t545 VPWR 565.638
R294 VPWR VPWR.t4580 565.638
R295 VPWR VPWR.t2081 565.638
R296 VPWR VPWR.t2317 565.638
R297 VPWR.t1840 VPWR 565.638
R298 VPWR.t2445 VPWR 565.638
R299 VPWR.t2628 VPWR 565.638
R300 VPWR.t3940 VPWR 565.638
R301 VPWR.t2758 VPWR 565.638
R302 VPWR.t1704 VPWR 565.638
R303 VPWR.t4342 VPWR 565.638
R304 VPWR VPWR.t4828 565.638
R305 VPWR.t4312 VPWR.t4679 527.356
R306 VPWR.t3428 VPWR.t484 518.519
R307 VPWR.t2885 VPWR.t3428 518.519
R308 VPWR.t2822 VPWR.t2885 518.519
R309 VPWR.t2642 VPWR.t2822 518.519
R310 VPWR.t3269 VPWR.t2642 518.519
R311 VPWR.t3823 VPWR.t3269 518.519
R312 VPWR.t697 VPWR.t3823 518.519
R313 VPWR.t70 VPWR.t1443 518.519
R314 VPWR.t2185 VPWR.t70 518.519
R315 VPWR.t3028 VPWR.t2185 518.519
R316 VPWR.t4369 VPWR.t3028 518.519
R317 VPWR.t962 VPWR.t4369 518.519
R318 VPWR.t657 VPWR.t962 518.519
R319 VPWR.t2281 VPWR.t657 518.519
R320 VPWR.t1139 VPWR.t557 518.519
R321 VPWR.t3497 VPWR.t1139 518.519
R322 VPWR.t1358 VPWR.t3497 518.519
R323 VPWR.t620 VPWR.t1358 518.519
R324 VPWR.t1397 VPWR.t620 518.519
R325 VPWR.t4417 VPWR.t1397 518.519
R326 VPWR.t1013 VPWR.t4417 518.519
R327 VPWR.t5196 VPWR.t1445 518.519
R328 VPWR.t421 VPWR.t5196 518.519
R329 VPWR.t3099 VPWR.t421 518.519
R330 VPWR.t3965 VPWR.t3099 518.519
R331 VPWR.t2669 VPWR.t3965 518.519
R332 VPWR.t425 VPWR.t2669 518.519
R333 VPWR.t1899 VPWR.t425 518.519
R334 VPWR.t3089 VPWR.t2007 518.519
R335 VPWR.t3819 VPWR.t3089 518.519
R336 VPWR.t1298 VPWR.t3819 518.519
R337 VPWR.t641 VPWR.t1298 518.519
R338 VPWR.t3288 VPWR.t641 518.519
R339 VPWR.t4760 VPWR.t3288 518.519
R340 VPWR.t328 VPWR.t4760 518.519
R341 VPWR.t3033 VPWR.t2338 518.519
R342 VPWR.t5639 VPWR.t3033 518.519
R343 VPWR.t4260 VPWR.t5639 518.519
R344 VPWR.t316 VPWR.t4260 518.519
R345 VPWR.t1141 VPWR.t316 518.519
R346 VPWR.t2297 VPWR.t1141 518.519
R347 VPWR.t3540 VPWR.t2297 518.519
R348 VPWR.t5798 VPWR.t1075 518.519
R349 VPWR.t1813 VPWR.t5798 518.519
R350 VPWR.t365 VPWR.t1813 518.519
R351 VPWR.t2513 VPWR.t365 518.519
R352 VPWR.t2896 VPWR.t2513 518.519
R353 VPWR.t1393 VPWR.t2896 518.519
R354 VPWR.t68 VPWR.t1393 518.519
R355 VPWR.t5242 VPWR.t926 518.519
R356 VPWR.t2179 VPWR.t5242 518.519
R357 VPWR.t3166 VPWR.t2179 518.519
R358 VPWR.t5711 VPWR.t3166 518.519
R359 VPWR.t2961 VPWR.t5711 518.519
R360 VPWR.t2413 VPWR.t2961 518.519
R361 VPWR.t1061 VPWR.t2413 518.519
R362 VPWR.t1970 VPWR.t2117 518.519
R363 VPWR.t873 VPWR.t1970 518.519
R364 VPWR.t1567 VPWR.t873 518.519
R365 VPWR.t1085 VPWR.t1567 518.519
R366 VPWR.t2039 VPWR.t1085 518.519
R367 VPWR.t1241 VPWR.t2039 518.519
R368 VPWR.t3340 VPWR.t1241 518.519
R369 VPWR.t801 VPWR.t3052 518.519
R370 VPWR.t3756 VPWR.t801 518.519
R371 VPWR.t3908 VPWR.t3756 518.519
R372 VPWR.t693 VPWR.t3908 518.519
R373 VPWR.t1290 VPWR.t693 518.519
R374 VPWR.t2216 VPWR.t1290 518.519
R375 VPWR.t2109 VPWR.t2216 518.519
R376 VPWR.t2865 VPWR.t2233 518.519
R377 VPWR.t2390 VPWR.t2865 518.519
R378 VPWR.t3047 VPWR.t2390 518.519
R379 VPWR.t54 VPWR.t3047 518.519
R380 VPWR.t2698 VPWR.t54 518.519
R381 VPWR.t1857 VPWR.t2698 518.519
R382 VPWR.t4583 VPWR.t1857 518.519
R383 VPWR.t1026 VPWR.t2943 518.519
R384 VPWR.t1987 VPWR.t1026 518.519
R385 VPWR.t3955 VPWR.t1987 518.519
R386 VPWR.t1352 VPWR.t3955 518.519
R387 VPWR.t1800 VPWR.t1352 518.519
R388 VPWR.t1897 VPWR.t1800 518.519
R389 VPWR.t3594 VPWR.t1897 518.519
R390 VPWR.t3406 VPWR.t3188 518.519
R391 VPWR.t647 VPWR.t3406 518.519
R392 VPWR.t2725 VPWR.t647 518.519
R393 VPWR.t4000 VPWR.t2725 518.519
R394 VPWR.t1981 VPWR.t4000 518.519
R395 VPWR.t2564 VPWR.t1981 518.519
R396 VPWR.t4883 VPWR.t2564 518.519
R397 VPWR.t4244 VPWR.t742 518.519
R398 VPWR.t373 VPWR.t4244 518.519
R399 VPWR.t5345 VPWR.t373 518.519
R400 VPWR.t791 VPWR.t5345 518.519
R401 VPWR.t2 VPWR.t791 518.519
R402 VPWR.t6114 VPWR.t2 518.519
R403 VPWR.t482 VPWR.t6114 518.519
R404 VPWR.t1188 VPWR.t2582 518.519
R405 VPWR.t2754 VPWR.t1188 518.519
R406 VPWR.t780 VPWR.t2754 518.519
R407 VPWR.t3104 VPWR.t780 518.519
R408 VPWR.t746 VPWR.t3104 518.519
R409 VPWR.t3744 VPWR.t746 518.519
R410 VPWR.t2610 VPWR.t3744 518.519
R411 VPWR.t5464 VPWR.t1377 518.519
R412 VPWR.t4167 VPWR.t5464 518.519
R413 VPWR.t3039 VPWR.t4167 518.519
R414 VPWR.t383 VPWR.t3039 518.519
R415 VPWR.t1362 VPWR.t383 518.519
R416 VPWR.t1459 VPWR.t1362 518.519
R417 VPWR.t1757 VPWR.t1459 518.519
R418 VPWR.t6361 VPWR.t3074 518.519
R419 VPWR.t78 VPWR.t3501 518.519
R420 VPWR.t3501 VPWR.t655 518.519
R421 VPWR.t655 VPWR.t1547 518.519
R422 VPWR.t1547 VPWR.t3785 518.519
R423 VPWR.t3785 VPWR.t5572 518.519
R424 VPWR.t5572 VPWR.t1218 518.519
R425 VPWR.t1218 VPWR.t1916 518.519
R426 VPWR.t4285 VPWR.t3430 518.519
R427 VPWR.t3742 VPWR.t4285 518.519
R428 VPWR.t1607 VPWR.t3742 518.519
R429 VPWR.t2663 VPWR.t1607 518.519
R430 VPWR.t1999 VPWR.t2663 518.519
R431 VPWR.t2015 VPWR.t1999 518.519
R432 VPWR.t86 VPWR.t2015 518.519
R433 VPWR.t2620 VPWR.t2872 518.519
R434 VPWR.t1165 VPWR.t2620 518.519
R435 VPWR.t4177 VPWR.t1165 518.519
R436 VPWR.t1149 VPWR.t2521 518.519
R437 VPWR.t1936 VPWR.t2466 518.519
R438 VPWR.t490 VPWR.t397 518.519
R439 VPWR.t1573 VPWR.t928 518.519
R440 VPWR.t4994 VPWR.t361 518.519
R441 VPWR.t1476 VPWR.t2127 518.519
R442 VPWR.t5901 VPWR.t1476 518.519
R443 VPWR.t1237 VPWR.t5901 518.519
R444 VPWR.t3369 VPWR.t1237 518.519
R445 VPWR.t2991 VPWR.t3369 518.519
R446 VPWR.t666 VPWR.t2991 518.519
R447 VPWR.t3600 VPWR.t666 518.519
R448 VPWR.t1143 VPWR.t1441 518.519
R449 VPWR.t1441 VPWR.t502 518.519
R450 VPWR.t1901 VPWR.t2491 518.519
R451 VPWR.t415 VPWR.t1901 518.519
R452 VPWR.t1643 VPWR.t415 518.519
R453 VPWR.t731 VPWR.t1643 518.519
R454 VPWR.t1735 VPWR.t731 518.519
R455 VPWR.t3803 VPWR.t1735 518.519
R456 VPWR.t1972 VPWR.t3803 518.519
R457 VPWR.t1036 VPWR.t4409 518.519
R458 VPWR.t5291 VPWR.t1036 518.519
R459 VPWR.t1721 VPWR.t2247 518.519
R460 VPWR.t58 VPWR.t1721 518.519
R461 VPWR.t1989 VPWR.t58 518.519
R462 VPWR.t4066 VPWR.t1989 518.519
R463 VPWR.t3859 VPWR.t4066 518.519
R464 VPWR.t4621 VPWR.t3859 518.519
R465 VPWR.t2791 VPWR.t2941 518.519
R466 VPWR.t4712 VPWR.t2791 518.519
R467 VPWR.t1253 VPWR.t4712 518.519
R468 VPWR.t4443 VPWR.t1253 518.519
R469 VPWR.t3511 VPWR.t4443 518.519
R470 VPWR.t2963 VPWR.t3511 518.519
R471 VPWR.t1081 VPWR.t2963 518.519
R472 VPWR.t590 VPWR.t3787 518.519
R473 VPWR.t3787 VPWR.t4307 518.519
R474 VPWR.t4307 VPWR.t1781 518.519
R475 VPWR.t3566 VPWR.t1224 518.519
R476 VPWR.t1044 VPWR.t3566 518.519
R477 VPWR.t975 VPWR.t1044 518.519
R478 VPWR.t348 VPWR.t975 518.519
R479 VPWR.t393 VPWR.t348 518.519
R480 VPWR.t3204 VPWR.t393 518.519
R481 VPWR.t3037 VPWR.t3204 518.519
R482 VPWR.t4100 VPWR.t580 518.519
R483 VPWR.t1391 VPWR.t4100 518.519
R484 VPWR.t1335 VPWR.t1391 518.519
R485 VPWR.t2527 VPWR.t1335 518.519
R486 VPWR.t3385 VPWR.t2527 518.519
R487 VPWR.t3980 VPWR.t3385 518.519
R488 VPWR.t3902 VPWR.t3980 518.519
R489 VPWR.t5034 VPWR.t1401 518.519
R490 VPWR.t2731 VPWR.t5034 518.519
R491 VPWR.t1615 VPWR.t2731 518.519
R492 VPWR.t5819 VPWR.t1615 518.519
R493 VPWR.t3454 VPWR.t5819 518.519
R494 VPWR.t3432 VPWR.t3454 518.519
R495 VPWR.t2340 VPWR.t3432 518.519
R496 VPWR.t995 VPWR.t4213 518.519
R497 VPWR.t5505 VPWR.t995 518.519
R498 VPWR.t1208 VPWR.t5505 518.519
R499 VPWR.t3689 VPWR.t1208 518.519
R500 VPWR.t3102 VPWR.t3689 518.519
R501 VPWR.t2839 VPWR.t3102 518.519
R502 VPWR.t5306 VPWR.t2839 518.519
R503 VPWR.t4054 VPWR.t3377 518.519
R504 VPWR.t3436 VPWR.t4054 518.519
R505 VPWR.t891 VPWR.t3436 518.519
R506 VPWR.t997 VPWR.t891 518.519
R507 VPWR.t677 VPWR.t997 518.519
R508 VPWR.t3116 VPWR.t677 518.519
R509 VPWR.t2495 VPWR.t3116 518.519
R510 VPWR.t4169 VPWR.t4725 518.519
R511 VPWR.t1052 VPWR.t4169 518.519
R512 VPWR.t3381 VPWR.t1052 518.519
R513 VPWR.t1419 VPWR.t3381 518.519
R514 VPWR.t2464 VPWR.t1419 518.519
R515 VPWR.t1226 VPWR.t2464 518.519
R516 VPWR.t346 VPWR.t1226 518.519
R517 VPWR.t1579 VPWR.t4010 518.519
R518 VPWR.t578 VPWR.t1579 518.519
R519 VPWR.t883 VPWR.t578 518.519
R520 VPWR.t989 VPWR.t883 518.519
R521 VPWR.t1342 VPWR.t989 518.519
R522 VPWR.t3967 VPWR.t1342 518.519
R523 VPWR.t5077 VPWR.t3967 518.519
R524 VPWR.t417 VPWR.t651 518.519
R525 VPWR.t3696 VPWR.t417 518.519
R526 VPWR.t4764 VPWR.t3696 518.519
R527 VPWR.t2905 VPWR.t4764 518.519
R528 VPWR.t1934 VPWR.t2905 518.519
R529 VPWR.t766 VPWR.t1934 518.519
R530 VPWR.t930 VPWR.t766 518.519
R531 VPWR.t1978 VPWR.t576 518.519
R532 VPWR.t3976 VPWR.t1978 518.519
R533 VPWR.t326 VPWR.t3976 518.519
R534 VPWR.t5274 VPWR.t1871 518.519
R535 VPWR.t1611 VPWR.t5274 518.519
R536 VPWR.t2676 VPWR.t1611 518.519
R537 VPWR.t809 VPWR.t2676 518.519
R538 VPWR.t940 VPWR.t809 518.519
R539 VPWR.t4852 VPWR.t1806 518.519
R540 VPWR.t1631 VPWR.t4852 518.519
R541 VPWR.t1509 VPWR.t1631 518.519
R542 VPWR.t1559 VPWR.t1509 518.519
R543 VPWR.t4305 VPWR.t1559 518.519
R544 VPWR.t66 VPWR.t4305 518.519
R545 VPWR.t3640 VPWR.t1147 518.519
R546 VPWR.t1894 VPWR.t3640 518.519
R547 VPWR.t3703 VPWR.t1894 518.519
R548 VPWR.t699 VPWR.t3703 518.519
R549 VPWR.t450 VPWR.t699 518.519
R550 VPWR.t5030 VPWR.t450 518.519
R551 VPWR.t423 VPWR.t5030 518.519
R552 VPWR.t1346 VPWR.t2011 518.519
R553 VPWR.t1968 VPWR.t1346 518.519
R554 VPWR.t3951 VPWR.t1968 518.519
R555 VPWR.t1974 VPWR.t3951 518.519
R556 VPWR.t1495 VPWR.t1974 518.519
R557 VPWR.t1569 VPWR.t1495 518.519
R558 VPWR.t1543 VPWR.t1569 518.519
R559 VPWR.t1696 VPWR.t381 518.519
R560 VPWR.t2489 VPWR.t1696 518.519
R561 VPWR.t893 VPWR.t2489 518.519
R562 VPWR.t2982 VPWR.t893 518.519
R563 VPWR.t5546 VPWR.t2982 518.519
R564 VPWR.t338 VPWR.t5546 518.519
R565 VPWR.t1657 VPWR.t338 518.519
R566 VPWR.t486 VPWR.t5876 518.519
R567 VPWR.t3110 VPWR.t4130 518.519
R568 VPWR.t1243 VPWR.t3110 518.519
R569 VPWR.t1296 VPWR.t1243 518.519
R570 VPWR.t1539 VPWR.t1296 518.519
R571 VPWR.t964 VPWR.t1539 518.519
R572 VPWR.t529 VPWR.t964 518.519
R573 VPWR.t3076 VPWR.t529 518.519
R574 VPWR.t689 VPWR.t2509 518.519
R575 VPWR.t2509 VPWR.t5244 518.519
R576 VPWR.t5244 VPWR.t862 518.519
R577 VPWR.t1097 VPWR.t5361 518.519
R578 VPWR.t1009 VPWR.t1097 518.519
R579 VPWR.t1282 VPWR.t1009 518.519
R580 VPWR.t2099 VPWR.t1771 518.519
R581 VPWR.t1771 VPWR.t821 518.519
R582 VPWR.t821 VPWR.t2551 518.519
R583 VPWR.t2551 VPWR.t1065 518.519
R584 VPWR.t1065 VPWR.t762 518.519
R585 VPWR.t762 VPWR.t456 518.519
R586 VPWR.t456 VPWR.t914 518.519
R587 VPWR.t2936 VPWR.t2945 518.519
R588 VPWR.t2910 VPWR.t4146 518.519
R589 VPWR.t3085 VPWR.t2910 518.519
R590 VPWR.t2194 VPWR.t3085 518.519
R591 VPWR.t3127 VPWR.t2194 518.519
R592 VPWR.t5874 VPWR.t2235 518.519
R593 VPWR.t4931 VPWR.t5874 518.519
R594 VPWR.t924 VPWR.t4931 518.519
R595 VPWR.t1251 VPWR.t924 518.519
R596 VPWR.t2409 VPWR.t1251 518.519
R597 VPWR.t2072 VPWR.t2409 518.519
R598 VPWR.t5308 VPWR.t2072 518.519
R599 VPWR.t912 VPWR.t2314 518.519
R600 VPWR.t673 VPWR.t912 518.519
R601 VPWR.t4300 VPWR.t673 518.519
R602 VPWR.t1702 VPWR.t4300 518.519
R603 VPWR.t574 VPWR.t1702 518.519
R604 VPWR.t1700 VPWR.t1114 518.519
R605 VPWR.t1823 VPWR.t1700 518.519
R606 VPWR.t2690 VPWR.t1823 518.519
R607 VPWR.t4262 VPWR.t2690 518.519
R608 VPWR.t3691 VPWR.t4262 518.519
R609 VPWR.t3136 VPWR.t3691 518.519
R610 VPWR.t5972 VPWR.t3136 518.519
R611 VPWR.t4612 VPWR.t2042 518.519
R612 VPWR.t1190 VPWR.t4612 518.519
R613 VPWR.t1186 VPWR.t1190 518.519
R614 VPWR.t2624 VPWR.t1186 518.519
R615 VPWR.t952 VPWR.t2624 518.519
R616 VPWR.t1145 VPWR.t952 518.519
R617 VPWR.t1629 VPWR.t2606 518.519
R618 VPWR.t2606 VPWR.t1484 518.519
R619 VPWR.t1484 VPWR.t1284 518.519
R620 VPWR.t1284 VPWR.t389 518.519
R621 VPWR.t389 VPWR.t512 518.519
R622 VPWR.t512 VPWR.t1551 518.519
R623 VPWR.t1551 VPWR.t549 518.519
R624 VPWR.t649 VPWR.t4249 518.519
R625 VPWR.t2279 VPWR.t649 518.519
R626 VPWR.t76 VPWR.t2279 518.519
R627 VPWR.t356 VPWR.t76 518.519
R628 VPWR.t1300 VPWR.t356 518.519
R629 VPWR.t1364 VPWR.t1300 518.519
R630 VPWR.t1507 VPWR.t1364 518.519
R631 VPWR.n1572 VPWR 515.444
R632 VPWR VPWR.n1534 515.444
R633 VPWR.n1029 VPWR 515.444
R634 VPWR.t6227 VPWR.t4677 501.932
R635 VPWR VPWR.t1379 501.932
R636 VPWR.t7050 VPWR.t6145 501.932
R637 VPWR.t4671 VPWR.t10 501.932
R638 VPWR.t691 VPWR.n2326 490.947
R639 VPWR.n266 VPWR.t2974 490.947
R640 VPWR.t6897 VPWR 482.625
R641 VPWR.t1739 VPWR.t1737 482.625
R642 VPWR.t7107 VPWR.t2356 478.764
R643 VPWR.t23 VPWR.t2529 478.764
R644 VPWR.t6 VPWR.t5652 478.764
R645 VPWR.t6521 VPWR.t6514 471.043
R646 VPWR.t3664 VPWR.t3662 471.043
R647 VPWR.t6524 VPWR.t6516 471.043
R648 VPWR.t6786 VPWR.t6785 471.043
R649 VPWR.t1202 VPWR.t1204 471.043
R650 VPWR.t6782 VPWR.t6781 471.043
R651 VPWR.t2113 VPWR.t88 463.32
R652 VPWR.n953 VPWR.t2553 462.151
R653 VPWR.t5931 VPWR.t2360 451.738
R654 VPWR.t6621 VPWR.t5927 451.738
R655 VPWR.t3559 VPWR.t6771 451.738
R656 VPWR.t6972 VPWR.t108 451.738
R657 VPWR.t5831 VPWR.t6622 451.738
R658 VPWR.t6899 VPWR.t6672 451.738
R659 VPWR.t7021 VPWR.t6764 451.738
R660 VPWR.t222 VPWR.t4148 446.76
R661 VPWR.t127 VPWR.t4264 446.76
R662 VPWR.t2417 VPWR.t5615 442.13
R663 VPWR.t2892 VPWR.t6453 442.13
R664 VPWR.t985 VPWR.t5252 442.13
R665 VPWR.t871 VPWR.t215 435.185
R666 VPWR.t3321 VPWR.t6817 432.433
R667 VPWR.t6139 VPWR.t6141 432.433
R668 VPWR.t6143 VPWR.t6139 432.433
R669 VPWR.t6145 VPWR.t6143 432.433
R670 VPWR.t7052 VPWR.t7050 432.433
R671 VPWR.t52 VPWR.t1437 432.433
R672 VPWR.t3239 VPWR.t7048 432.433
R673 VPWR.t4669 VPWR.t4673 432.433
R674 VPWR.t4673 VPWR.t4675 432.433
R675 VPWR.t4675 VPWR.t4671 432.433
R676 VPWR.t10 VPWR.t8 432.433
R677 VPWR.t5455 VPWR.t179 432.433
R678 VPWR.t5599 VPWR 418.981
R679 VPWR.t1747 VPWR.t3251 418.981
R680 VPWR.t470 VPWR.t3118 416.668
R681 VPWR.t4679 VPWR.t6227 413.127
R682 VPWR.t2439 VPWR.t5049 402.779
R683 VPWR.t207 VPWR 396.991
R684 VPWR.t195 VPWR 396.991
R685 VPWR.t6189 VPWR.t1360 395.834
R686 VPWR.t4677 VPWR.t4314 393.822
R687 VPWR.t3666 VPWR.t6521 393.822
R688 VPWR.t6514 VPWR.t3664 393.822
R689 VPWR.t3662 VPWR.t6524 393.822
R690 VPWR.t6516 VPWR.t3660 393.822
R691 VPWR.t6785 VPWR.t1206 393.822
R692 VPWR.t1204 VPWR.t6786 393.822
R693 VPWR.t6781 VPWR.t1202 393.822
R694 VPWR.t1200 VPWR.t6782 393.822
R695 VPWR.t2356 VPWR.t45 393.822
R696 VPWR.t6627 VPWR.t6578 393.822
R697 VPWR.t6903 VPWR.t6897 393.822
R698 VPWR.n798 VPWR.n749 393.091
R699 VPWR.n1439 VPWR.n1397 389.106
R700 VPWR.n907 VPWR.n827 389.106
R701 VPWR.n2795 VPWR.n2748 389.106
R702 VPWR.t3430 VPWR.n3435 388.889
R703 VPWR.t2901 VPWR.t3315 388.889
R704 VPWR.t1234 VPWR.t3434 388.889
R705 VPWR.t2415 VPWR.t4052 388.889
R706 VPWR.t5498 VPWR.t3202 388.889
R707 VPWR.t1413 VPWR.t3945 388.889
R708 VPWR.t5775 VPWR.t1593 388.889
R709 VPWR.t600 VPWR.t6458 388.889
R710 VPWR.t5281 VPWR.t2431 388.889
R711 VPWR.t4127 VPWR.t5531 388.889
R712 VPWR.t6210 VPWR.t4592 388.889
R713 VPWR.t5861 VPWR.t703 388.889
R714 VPWR.t993 VPWR.t2947 388.889
R715 VPWR.t4935 VPWR.t4954 388.889
R716 VPWR.t4340 VPWR.t4888 388.889
R717 VPWR.t1712 VPWR.t570 388.889
R718 VPWR.t823 VPWR.t4097 388.889
R719 VPWR.t1385 VPWR.t2678 388.889
R720 VPWR.t5299 VPWR.t6349 388.889
R721 VPWR.t3644 VPWR.t4391 388.889
R722 VPWR.t5636 VPWR.t1851 388.889
R723 VPWR.t4485 VPWR.t2385 388.889
R724 VPWR.t330 VPWR.t3499 388.889
R725 VPWR.t5780 VPWR.t4058 388.889
R726 VPWR.t2531 VPWR.t5099 388.889
R727 VPWR.t721 VPWR.t5414 388.889
R728 VPWR.t709 VPWR.t1395 388.889
R729 VPWR.t1505 VPWR.t1960 388.889
R730 VPWR.t1827 VPWR.t701 388.889
R731 VPWR.t4943 VPWR.t3921 388.889
R732 VPWR.t2097 VPWR.t1605 388.889
R733 VPWR.t3387 VPWR.t875 388.889
R734 VPWR.t631 VPWR.t2535 388.889
R735 VPWR.t2089 VPWR.t1985 388.889
R736 VPWR.t4926 VPWR.n1937 388.889
R737 VPWR.t2853 VPWR.t4739 388.889
R738 VPWR.t2515 VPWR.n2861 388.889
R739 VPWR.t1879 VPWR.t2142 388.889
R740 VPWR.t4906 VPWR.t604 388.889
R741 VPWR.t1447 VPWR.t1171 388.889
R742 VPWR.t1276 VPWR.t1773 388.889
R743 VPWR.t4357 VPWR.t3515 388.889
R744 VPWR.t2756 VPWR.t5678 388.889
R745 VPWR.t5768 VPWR.t723 388.889
R746 VPWR.t2517 VPWR.t4367 388.889
R747 VPWR.t2319 VPWR.t2429 388.889
R748 VPWR.t5699 VPWR.t6193 388.889
R749 VPWR.t6000 VPWR.t756 388.889
R750 VPWR.t2009 VPWR.t1133 388.889
R751 VPWR.t4539 VPWR.t4969 388.889
R752 VPWR.t3225 VPWR.t1449 388.889
R753 VPWR.t4918 VPWR.t1278 388.889
R754 VPWR.t458 VPWR.t4361 388.889
R755 VPWR.t5770 VPWR.t3246 388.889
R756 VPWR.t4162 VPWR.t4031 388.889
R757 VPWR.t1844 VPWR.t3262 388.889
R758 VPWR.t494 VPWR.t427 388.889
R759 VPWR.t5709 VPWR.t2661 388.889
R760 VPWR.t4238 VPWR.t6282 388.889
R761 VPWR.t3186 VPWR.t3546 388.889
R762 VPWR.t4545 VPWR.t4353 388.889
R763 VPWR.t5724 VPWR.t681 388.889
R764 VPWR.t6159 VPWR.t1474 388.889
R765 VPWR.t4189 VPWR.t1706 388.889
R766 VPWR.t2132 VPWR.t1228 388.889
R767 VPWR.t1007 VPWR.t5036 388.889
R768 VPWR.t5840 VPWR.t4758 388.889
R769 VPWR.t2888 VPWR.t2200 388.889
R770 VPWR.t1089 VPWR.t4766 388.889
R771 VPWR.t3190 VPWR.t3093 388.889
R772 VPWR.t3815 VPWR.t782 388.889
R773 VPWR.t2471 VPWR.t3774 388.889
R774 VPWR.t2493 VPWR.t3364 388.889
R775 VPWR.t5452 VPWR.t4940 388.889
R776 VPWR.t3886 VPWR.t944 388.889
R777 VPWR.t4814 VPWR.t4253 388.889
R778 VPWR.t1765 VPWR.t5541 388.889
R779 VPWR.t4861 VPWR.t6150 388.889
R780 VPWR.t4706 VPWR.t5481 388.889
R781 VPWR.t2212 VPWR.t2056 388.889
R782 VPWR.t744 VPWR.t1421 388.889
R783 VPWR.t6109 VPWR.t3588 388.889
R784 VPWR.t5060 VPWR.t3213 388.889
R785 VPWR.t4008 VPWR.t3626 388.889
R786 VPWR.t5630 VPWR.t3596 388.889
R787 VPWR.t4351 VPWR.t4589 388.889
R788 VPWR.t6218 VPWR.t4454 388.889
R789 VPWR.t60 VPWR.t6208 388.889
R790 VPWR.t3725 VPWR.t3807 388.889
R791 VPWR.t1654 VPWR.t4024 388.889
R792 VPWR.t3817 VPWR.t4525 388.889
R793 VPWR.t2626 VPWR.t675 388.889
R794 VPWR.t6191 VPWR.t4874 388.889
R795 VPWR.t4490 VPWR.t3353 388.889
R796 VPWR.t4614 VPWR.t6053 388.889
R797 VPWR.t4151 VPWR.t3168 388.889
R798 VPWR.t1853 VPWR.t5272 388.889
R799 VPWR.t6083 VPWR.t1670 388.889
R800 VPWR.t1249 VPWR.t2923 388.889
R801 VPWR.t472 VPWR.t5668 388.889
R802 VPWR.t3451 VPWR.t3379 388.889
R803 VPWR.t3947 VPWR.t829 388.889
R804 VPWR.t2060 VPWR.t4640 388.889
R805 VPWR.t498 VPWR.t2449 388.889
R806 VPWR.t7085 VPWR.t492 388.889
R807 VPWR.t391 VPWR.t3855 388.889
R808 VPWR.t4929 VPWR.t1194 388.889
R809 VPWR.t5955 VPWR.t1925 388.889
R810 VPWR.t2229 VPWR.t2192 388.889
R811 VPWR.t2407 VPWR.t4543 388.889
R812 VPWR.t1417 VPWR.t5107 388.889
R813 VPWR.t3466 VPWR.t7123 388.889
R814 VPWR.t4806 VPWR.t3333 388.889
R815 VPWR.t5359 VPWR.t4458 388.889
R816 VPWR.t4594 VPWR.t4636 388.889
R817 VPWR.t3035 VPWR.t2249 388.889
R818 VPWR.t6085 VPWR.t2425 388.889
R819 VPWR.t1247 VPWR.t5766 388.889
R820 VPWR.t3194 VPWR.t1678 388.889
R821 VPWR.t4920 VPWR.t1274 388.889
R822 VPWR.t679 VPWR.t807 388.889
R823 VPWR.t2451 VPWR.t4643 388.889
R824 VPWR.t5943 VPWR.t2017 388.889
R825 VPWR.t533 VPWR.t3537 388.889
R826 VPWR.t2473 VPWR.t5555 388.889
R827 VPWR.t5605 VPWR.t5449 388.889
R828 VPWR.t1183 VPWR.t5509 388.889
R829 VPWR.t3443 VPWR.t3673 388.889
R830 VPWR.t4504 VPWR.t1680 388.889
R831 VPWR.t1286 VPWR.t72 388.889
R832 VPWR.t1409 VPWR.t6307 388.889
R833 VPWR.t1555 VPWR.t871 388.889
R834 VPWR.t2441 VPWR.t5759 388.889
R835 VPWR.t592 VPWR.t2190 388.889
R836 VPWR.t2146 VPWR.t3714 388.889
R837 VPWR.t1482 VPWR.t2105 388.889
R838 VPWR.t4571 VPWR.t815 388.889
R839 VPWR.t5301 VPWR.t4119 388.889
R840 VPWR.t5026 VPWR.t1815 388.889
R841 VPWR.t660 VPWR.t3249 388.889
R842 VPWR.t1344 VPWR.t4121 388.889
R843 VPWR.t2156 VPWR.t1888 388.889
R844 VPWR.t2382 VPWR.t555 388.889
R845 VPWR.t869 VPWR.t713 388.889
R846 VPWR.t312 VPWR.t5755 388.889
R847 VPWR.t4845 VPWR.t5937 388.889
R848 VPWR.t5367 VPWR.t369 388.889
R849 VPWR.t564 VPWR.t4663 388.889
R850 VPWR.t740 VPWR.t3418 388.889
R851 VPWR.t6105 VPWR.t5903 388.889
R852 VPWR.t6017 VPWR.t2700 388.889
R853 VPWR.t1501 VPWR.t1884 388.889
R854 VPWR.t6324 VPWR.t5503 388.889
R855 VPWR.t1059 VPWR.t4336 388.889
R856 VPWR.t3953 VPWR.t5333 388.889
R857 VPWR.t1122 VPWR.t770 388.889
R858 VPWR.t1641 VPWR.t5537 388.889
R859 VPWR.t7069 VPWR.t3062 388.889
R860 VPWR.t4518 VPWR.t2832 388.889
R861 VPWR.t602 VPWR.t6103 388.889
R862 VPWR.t1871 VPWR.n2065 388.889
R863 VPWR.t387 VPWR.n199 388.889
R864 VPWR.t1806 VPWR.n201 388.889
R865 VPWR.t2011 VPWR.n207 388.889
R866 VPWR.t4894 VPWR.t4073 388.889
R867 VPWR.t2079 VPWR.t1001 388.889
R868 VPWR.t2908 VPWR.t3846 388.889
R869 VPWR.t4647 VPWR.t2136 388.889
R870 VPWR.t2938 VPWR.t1370 388.889
R871 VPWR.t3614 VPWR.t4034 388.889
R872 VPWR.t4710 VPWR.t6187 388.889
R873 VPWR.t3458 VPWR.t2214 388.889
R874 VPWR.t5644 VPWR.t3043 388.889
R875 VPWR.t5953 VPWR.t4950 388.889
R876 VPWR.t2221 VPWR.t2025 388.889
R877 VPWR.t4332 VPWR.t5335 388.889
R878 VPWR.t2251 VPWR.t3509 388.889
R879 VPWR.t4424 VPWR.t2443 388.889
R880 VPWR.t4179 VPWR.t2723 388.889
R881 VPWR.t4727 VPWR.t1647 388.889
R882 VPWR.t1798 VPWR.t2819 388.889
R883 VPWR.t1715 VPWR.t3210 388.889
R884 VPWR.t4199 VPWR.t3556 388.889
R885 VPWR.t4900 VPWR.t2549 388.889
R886 VPWR.t2013 VPWR.t3917 388.889
R887 VPWR.t5750 VPWR.t5731 388.889
R888 VPWR.t4632 VPWR.t1003 388.889
R889 VPWR.t598 VPWR.t4596 388.889
R890 VPWR.t4616 VPWR.t6133 388.889
R891 VPWR.t3009 VPWR.t3864 388.889
R892 VPWR.t2984 VPWR.t2720 388.889
R893 VPWR.t5681 VPWR.t6358 388.889
R894 VPWR.t2327 VPWR.t84 388.889
R895 VPWR.t2295 VPWR.t4022 388.889
R896 VPWR.t7075 VPWR.t3620 388.889
R897 VPWR.t3548 VPWR.t3776 388.889
R898 VPWR.t5361 VPWR.n2427 388.889
R899 VPWR.n2429 VPWR.t2099 388.889
R900 VPWR.n261 VPWR.t2685 388.889
R901 VPWR.t4146 VPWR.n2536 388.889
R902 VPWR.t2235 VPWR.n2538 388.889
R903 VPWR.t2103 VPWR.n2540 388.889
R904 VPWR.t2314 VPWR.n1 388.889
R905 VPWR.t1114 VPWR.n31 388.889
R906 VPWR.t2972 VPWR.n33 388.889
R907 VPWR.t2042 VPWR.n35 388.889
R908 VPWR.t4249 VPWR.n88 388.889
R909 VPWR VPWR.t6885 385.418
R910 VPWR VPWR.t3848 369.214
R911 VPWR.t3223 VPWR 369.214
R912 VPWR VPWR.t5716 366.899
R913 VPWR VPWR.t6057 366.899
R914 VPWR VPWR.t206 366.899
R915 VPWR.t2523 VPWR 366.899
R916 VPWR.t537 VPWR 366.899
R917 VPWR VPWR.t1515 366.899
R918 VPWR.t1710 VPWR 366.899
R919 VPWR.t5835 VPWR.t6671 361.111
R920 VPWR.n151 VPWR.t5855 358.796
R921 VPWR.t5248 VPWR.t2064 358.796
R922 VPWR VPWR.t205 355.325
R923 VPWR.t3003 VPWR 355.325
R924 VPWR.n1523 VPWR 349.421
R925 VPWR.n1524 VPWR 349.421
R926 VPWR VPWR.n1524 349.421
R927 VPWR.n1526 VPWR 349.421
R928 VPWR VPWR.n1571 349.421
R929 VPWR.n1534 VPWR 349.421
R930 VPWR.n1542 VPWR 349.421
R931 VPWR.n1064 VPWR 349.421
R932 VPWR.n1064 VPWR 349.421
R933 VPWR VPWR.n1029 349.421
R934 VPWR VPWR.n1026 349.421
R935 VPWR.n1026 VPWR 349.421
R936 VPWR VPWR.n1022 349.421
R937 VPWR.n1507 VPWR 349.421
R938 VPWR.n1508 VPWR 349.421
R939 VPWR.n2327 VPWR 349.421
R940 VPWR.n2328 VPWR 349.421
R941 VPWR.n2329 VPWR 349.421
R942 VPWR.n2330 VPWR 349.421
R943 VPWR.n2956 VPWR 349.421
R944 VPWR.n2957 VPWR 349.421
R945 VPWR.n2958 VPWR 349.421
R946 VPWR.n2959 VPWR 349.421
R947 VPWR.n2480 VPWR 349.421
R948 VPWR.n2481 VPWR 349.421
R949 VPWR.n2482 VPWR 349.421
R950 VPWR VPWR.n257 349.421
R951 VPWR.n2620 VPWR 349.421
R952 VPWR.n2621 VPWR 349.421
R953 VPWR.n2623 VPWR 349.421
R954 VPWR VPWR.n2622 349.421
R955 VPWR VPWR.n5 349.421
R956 VPWR.n6 VPWR 349.421
R957 VPWR.n39 VPWR 349.421
R958 VPWR.n57 VPWR 349.421
R959 VPWR.n58 VPWR 349.421
R960 VPWR.n59 VPWR 349.421
R961 VPWR.n3686 VPWR 349.421
R962 VPWR.t1617 VPWR.t6865 346.065
R963 VPWR.t6398 VPWR.t5642 346.065
R964 VPWR.t1956 VPWR.t3564 344.908
R965 VPWR VPWR.t1424 343.75
R966 VPWR VPWR.t1838 339.12
R967 VPWR.t484 VPWR 339.12
R968 VPWR VPWR.t4904 339.12
R969 VPWR.t1443 VPWR 339.12
R970 VPWR VPWR.t4385 339.12
R971 VPWR.t557 VPWR 339.12
R972 VPWR VPWR.t4627 339.12
R973 VPWR.t1445 VPWR 339.12
R974 VPWR VPWR.t4492 339.12
R975 VPWR.t2007 VPWR 339.12
R976 VPWR VPWR.t4113 339.12
R977 VPWR.t2338 VPWR 339.12
R978 VPWR VPWR.t2665 339.12
R979 VPWR.t1075 VPWR 339.12
R980 VPWR VPWR.t1745 339.12
R981 VPWR.t926 VPWR 339.12
R982 VPWR VPWR.t2616 339.12
R983 VPWR.t2117 VPWR 339.12
R984 VPWR VPWR.t3464 339.12
R985 VPWR.t3052 VPWR 339.12
R986 VPWR VPWR.t1783 339.12
R987 VPWR.t2233 VPWR 339.12
R988 VPWR VPWR.t3260 339.12
R989 VPWR.t2943 VPWR 339.12
R990 VPWR VPWR.t2405 339.12
R991 VPWR.t3188 VPWR 339.12
R992 VPWR VPWR.t6075 339.12
R993 VPWR.t742 VPWR 339.12
R994 VPWR VPWR.t5533 339.12
R995 VPWR.t2582 VPWR 339.12
R996 VPWR VPWR.t5550 339.12
R997 VPWR.t1377 VPWR 339.12
R998 VPWR VPWR.t2403 339.12
R999 VPWR VPWR.t78 339.12
R1000 VPWR.t633 VPWR 339.12
R1001 VPWR.t2872 VPWR 339.12
R1002 VPWR.t3456 VPWR 339.12
R1003 VPWR.t2521 VPWR 339.12
R1004 VPWR.t3748 VPWR 339.12
R1005 VPWR.t2466 VPWR 339.12
R1006 VPWR.t2795 VPWR 339.12
R1007 VPWR.t5028 VPWR 339.12
R1008 VPWR VPWR.t4334 339.12
R1009 VPWR.t3170 VPWR 339.12
R1010 VPWR VPWR.t490 339.12
R1011 VPWR VPWR.t1573 339.12
R1012 VPWR VPWR.t3646 339.12
R1013 VPWR.t361 VPWR 339.12
R1014 VPWR.t5433 VPWR 339.12
R1015 VPWR.t2127 VPWR 339.12
R1016 VPWR VPWR.t4537 339.12
R1017 VPWR VPWR.t1609 339.12
R1018 VPWR VPWR.t1143 339.12
R1019 VPWR.t4667 VPWR 339.12
R1020 VPWR VPWR.t1553 339.12
R1021 VPWR VPWR.t1159 339.12
R1022 VPWR VPWR.t6241 339.12
R1023 VPWR.t1755 VPWR 339.12
R1024 VPWR.t2491 VPWR 339.12
R1025 VPWR.t1663 VPWR 339.12
R1026 VPWR.t62 VPWR 339.12
R1027 VPWR.t4409 VPWR 339.12
R1028 VPWR.t2497 VPWR 339.12
R1029 VPWR.t1222 VPWR 339.12
R1030 VPWR.t1674 VPWR 339.12
R1031 VPWR.t3056 VPWR 339.12
R1032 VPWR.t2247 VPWR 339.12
R1033 VPWR.t5323 VPWR 339.12
R1034 VPWR.t4645 VPWR 339.12
R1035 VPWR VPWR.t5558 339.12
R1036 VPWR.t2941 VPWR 339.12
R1037 VPWR VPWR.t4195 339.12
R1038 VPWR VPWR.t4847 339.12
R1039 VPWR VPWR.t590 339.12
R1040 VPWR VPWR.t4018 339.12
R1041 VPWR VPWR.t2144 339.12
R1042 VPWR VPWR.t2269 339.12
R1043 VPWR.t3607 VPWR 339.12
R1044 VPWR.t1224 VPWR 339.12
R1045 VPWR VPWR.t1645 339.12
R1046 VPWR VPWR.t3853 339.12
R1047 VPWR.t4297 VPWR 339.12
R1048 VPWR.t6088 VPWR 339.12
R1049 VPWR.t488 VPWR 339.12
R1050 VPWR.t580 VPWR 339.12
R1051 VPWR.t1401 VPWR 339.12
R1052 VPWR.t4213 VPWR 339.12
R1053 VPWR.t3377 VPWR 339.12
R1054 VPWR.t3031 VPWR 339.12
R1055 VPWR.t7140 VPWR 339.12
R1056 VPWR.t3176 VPWR 339.12
R1057 VPWR VPWR.t1759 339.12
R1058 VPWR.t2299 VPWR 339.12
R1059 VPWR.t4725 VPWR 339.12
R1060 VPWR.t4010 VPWR 339.12
R1061 VPWR.t4267 VPWR 339.12
R1062 VPWR.t572 VPWR 339.12
R1063 VPWR.t651 VPWR 339.12
R1064 VPWR.t2074 VPWR 339.12
R1065 VPWR.t2411 VPWR 339.12
R1066 VPWR.t2172 VPWR 339.12
R1067 VPWR.t3760 VPWR 339.12
R1068 VPWR.t576 VPWR 339.12
R1069 VPWR VPWR.t2255 339.12
R1070 VPWR.t2709 VPWR 339.12
R1071 VPWR.t1147 VPWR 339.12
R1072 VPWR.t5561 VPWR 339.12
R1073 VPWR.t1890 VPWR 339.12
R1074 VPWR.t5945 VPWR 339.12
R1075 VPWR.t381 VPWR 339.12
R1076 VPWR.n181 VPWR 339.12
R1077 VPWR VPWR.t1831 339.12
R1078 VPWR VPWR.t486 339.12
R1079 VPWR.t2814 VPWR 339.12
R1080 VPWR.t4130 VPWR 339.12
R1081 VPWR VPWR.t1432 339.12
R1082 VPWR VPWR.t1175 339.12
R1083 VPWR VPWR.t689 339.12
R1084 VPWR VPWR.t2936 339.12
R1085 VPWR.t627 VPWR 339.12
R1086 VPWR VPWR.t1629 339.12
R1087 VPWR.t3182 VPWR.t6769 337.964
R1088 VPWR VPWR.t2271 336.807
R1089 VPWR VPWR.t3734 336.807
R1090 VPWR VPWR.t3066 336.807
R1091 VPWR.t2953 VPWR.t4309 333.776
R1092 VPWR.t7012 VPWR.t1320 333.334
R1093 VPWR.t2285 VPWR.t5393 333.334
R1094 VPWR.t94 VPWR.t3290 329.861
R1095 VPWR.t7059 VPWR.t2160 329.861
R1096 VPWR.t804 VPWR.t7043 329.861
R1097 VPWR.t1469 VPWR.t100 329.861
R1098 VPWR.t2352 VPWR.t2348 326.264
R1099 VPWR.t6031 VPWR.t221 325.231
R1100 VPWR.t6417 VPWR.n378 325.231
R1101 VPWR.t3323 VPWR.t3321 324.325
R1102 VPWR.t3325 VPWR.t3324 324.325
R1103 VPWR.t1437 VPWR.t1436 324.325
R1104 VPWR.t358 VPWR.t359 324.325
R1105 VPWR.t5519 VPWR.t5521 324.325
R1106 VPWR.t3241 VPWR.t3239 324.325
R1107 VPWR.t5970 VPWR.t5969 324.325
R1108 VPWR.t5454 VPWR.t5455 324.325
R1109 VPWR.t6894 VPWR.t4389 324.075
R1110 VPWR.t2337 VPWR.t6722 324.075
R1111 VPWR.t3285 VPWR.t17 324.075
R1112 VPWR.t7098 VPWR.t3146 322.918
R1113 VPWR.t6385 VPWR.t4902 322.918
R1114 VPWR.n1093 VPWR.t27 322.918
R1115 VPWR.t5747 VPWR.t161 322.918
R1116 VPWR.t6412 VPWR.t5752 322.741
R1117 VPWR.t96 VPWR.n935 317.13
R1118 VPWR.t6633 VPWR.t922 317.13
R1119 VPWR.t91 VPWR.t5276 317.13
R1120 VPWR.t1350 VPWR.t163 317.13
R1121 VPWR.t5221 VPWR.t98 317.13
R1122 VPWR.t6823 VPWR.t4269 317.13
R1123 VPWR.t4433 VPWR.t1589 314.815
R1124 VPWR.t1684 VPWR.t3972 314.815
R1125 VPWR.t1167 VPWR.t5157 314.815
R1126 VPWR.t5609 VPWR.t3338 314.815
R1127 VPWR.t849 VPWR 313.658
R1128 VPWR.t5544 VPWR.t2638 312.5
R1129 VPWR.t2419 VPWR.t1156 312.5
R1130 VPWR.t6363 VPWR.t4422 312.5
R1131 VPWR.t3983 VPWR.t2533 312.5
R1132 VPWR.t6901 VPWR.t6099 311.344
R1133 VPWR.t3158 VPWR.t4450 310.185
R1134 VPWR.t835 VPWR.t5085 310.185
R1135 VPWR.t2578 VPWR.t3934 310.185
R1136 VPWR VPWR.t4523 309.029
R1137 VPWR VPWR.t594 309.029
R1138 VPWR VPWR.t1222 309.029
R1139 VPWR VPWR.t470 309.029
R1140 VPWR VPWR.t4890 309.029
R1141 VPWR.t6817 VPWR 308.88
R1142 VPWR VPWR.t52 308.88
R1143 VPWR.t7048 VPWR 308.88
R1144 VPWR.t179 VPWR 308.88
R1145 VPWR.t5462 VPWR.n756 303.241
R1146 VPWR.t1849 VPWR.t877 303.241
R1147 VPWR.t4798 VPWR.t4132 300.926
R1148 VPWR VPWR.n1522 299.228
R1149 VPWR VPWR.t1163 299.228
R1150 VPWR VPWR.n1523 299.228
R1151 VPWR VPWR.t2287 299.228
R1152 VPWR VPWR.t1232 299.228
R1153 VPWR VPWR.t778 299.228
R1154 VPWR VPWR.t4153 299.228
R1155 VPWR VPWR.t1659 299.228
R1156 VPWR VPWR.n1526 299.228
R1157 VPWR VPWR.t5317 299.228
R1158 VPWR VPWR.t1312 299.228
R1159 VPWR.t4580 VPWR 299.228
R1160 VPWR.t1903 VPWR 299.228
R1161 VPWR.t2317 VPWR 299.228
R1162 VPWR.n1571 VPWR 299.228
R1163 VPWR VPWR.t543 299.228
R1164 VPWR VPWR.t1407 299.228
R1165 VPWR VPWR.t2628 299.228
R1166 VPWR VPWR.t1131 299.228
R1167 VPWR VPWR.t2758 299.228
R1168 VPWR VPWR.n1535 299.228
R1169 VPWR VPWR.t1028 299.228
R1170 VPWR VPWR.t5634 299.228
R1171 VPWR.t4242 VPWR 299.228
R1172 VPWR VPWR.t5283 299.228
R1173 VPWR.t4828 VPWR 299.228
R1174 VPWR.t5548 VPWR 299.228
R1175 VPWR VPWR.t5494 299.228
R1176 VPWR.n1508 VPWR 299.228
R1177 VPWR VPWR.t5811 299.228
R1178 VPWR VPWR.t3521 299.228
R1179 VPWR VPWR.t3938 299.228
R1180 VPWR VPWR.t4363 299.228
R1181 VPWR VPWR.t1829 299.228
R1182 VPWR VPWR.t4886 299.228
R1183 VPWR VPWR.t3740 299.228
R1184 VPWR VPWR.t1024 299.228
R1185 VPWR VPWR.t864 299.228
R1186 VPWR VPWR.t3926 299.228
R1187 VPWR.t3383 VPWR 299.228
R1188 VPWR VPWR.t867 299.228
R1189 VPWR VPWR.t5170 299.228
R1190 VPWR.t6322 VPWR 299.228
R1191 VPWR.t5129 VPWR 299.228
R1192 VPWR VPWR.t4788 299.228
R1193 VPWR VPWR.t1775 299.228
R1194 VPWR.t6448 VPWR 299.228
R1195 VPWR.t4535 VPWR 299.228
R1196 VPWR VPWR.t2154 299.228
R1197 VPWR VPWR.t3375 299.228
R1198 VPWR.t3699 VPWR 299.228
R1199 VPWR VPWR.t5650 299.228
R1200 VPWR VPWR.t2423 299.228
R1201 VPWR VPWR.t1091 299.228
R1202 VPWR.t2733 VPWR.t4117 298.611
R1203 VPWR.t1882 VPWR.t6400 298.611
R1204 VPWR.t1105 VPWR 292.825
R1205 VPWR.t5142 VPWR.t6511 290.822
R1206 VPWR.t4688 VPWR.t3022 290.822
R1207 VPWR.t21 VPWR 289.353
R1208 VPWR.t2271 VPWR.t2273 289.353
R1209 VPWR.t1067 VPWR.t1069 289.353
R1210 VPWR.t4831 VPWR.t4833 289.353
R1211 VPWR.t1270 VPWR.t1272 289.353
R1212 VPWR.t2398 VPWR.t2400 289.353
R1213 VPWR.t7018 VPWR.t3060 289.353
R1214 VPWR.t2525 VPWR.t2523 289.353
R1215 VPWR.t3734 VPWR.t3736 289.353
R1216 VPWR.t3072 VPWR.t3070 289.353
R1217 VPWR.t4413 VPWR.t4411 289.353
R1218 VPWR.t5319 VPWR.t5321 289.353
R1219 VPWR.t2914 VPWR.t2916 289.353
R1220 VPWR.t2828 VPWR.t2830 289.353
R1221 VPWR.t1493 VPWR.t1491 289.353
R1222 VPWR.t1639 VPWR.t1637 289.353
R1223 VPWR.t1708 VPWR.t1710 289.353
R1224 VPWR VPWR.t6580 289.353
R1225 VPWR.t310 VPWR.t308 289.353
R1226 VPWR.t1769 VPWR.t1767 289.353
R1227 VPWR.t5825 VPWR.t5827 289.353
R1228 VPWR.t1486 VPWR.t1488 289.353
R1229 VPWR.t3066 VPWR.t3068 289.353
R1230 VPWR.t6305 VPWR.t1651 287.038
R1231 VPWR.t6527 VPWR.t3473 287.038
R1232 VPWR.t5857 VPWR.t4071 287.038
R1233 VPWR.t37 VPWR.t2783 287.038
R1234 VPWR.t5914 VPWR.t3872 287.038
R1235 VPWR.t683 VPWR.t1314 287.038
R1236 VPWR.t5674 VPWR.t687 287.038
R1237 VPWR.t2778 VPWR.t1863 287.038
R1238 VPWR.t2890 VPWR.t5425 287.038
R1239 VPWR.t5701 VPWR.t1331 287.038
R1240 VPWR.t5603 VPWR.t1071 287.038
R1241 VPWR.t1455 VPWR.t5250 287.038
R1242 VPWR.t5949 VPWR.t5246 287.038
R1243 VPWR.t2764 VPWR.t6828 287.038
R1244 VPWR.t1511 VPWR.n198 287.038
R1245 VPWR.t5996 VPWR.t5160 287.038
R1246 VPWR.t5062 VPWR.t4037 282.408
R1247 VPWR.t5014 VPWR.t5018 282.408
R1248 VPWR.t5270 VPWR.t323 282.408
R1249 VPWR.t411 VPWR.t6855 282.408
R1250 VPWR.t6040 VPWR.t6046 282.408
R1251 VPWR.t1430 VPWR.t1426 282.408
R1252 VPWR.t1424 VPWR.t1428 282.408
R1253 VPWR.t399 VPWR.t405 282.408
R1254 VPWR.t4699 VPWR.t2951 282.408
R1255 VPWR.t1688 VPWR 281.25
R1256 VPWR VPWR.t2121 281.25
R1257 VPWR.t752 VPWR 281.25
R1258 VPWR.t4742 VPWR.t1383 280.094
R1259 VPWR.t805 VPWR.t6698 277.779
R1260 VPWR.t6595 VPWR 275.464
R1261 VPWR.t3582 VPWR.t6850 273.149
R1262 VPWR.t6718 VPWR.t1011 273.149
R1263 VPWR.t7030 VPWR 273.149
R1264 VPWR.t2586 VPWR.t6674 270.834
R1265 VPWR.t3481 VPWR.t106 270.834
R1266 VPWR.t6760 VPWR.t6738 270.834
R1267 VPWR.t7111 VPWR.t112 270.834
R1268 VPWR.t6587 VPWR.t6860 270.834
R1269 VPWR.t3020 VPWR.t3829 269.693
R1270 VPWR.t3896 VPWR.t3206 268.519
R1271 VPWR.t332 VPWR.t5975 268.519
R1272 VPWR.t6988 VPWR 267.861
R1273 VPWR VPWR.t3754 267.361
R1274 VPWR.t7096 VPWR 267.361
R1275 VPWR.t6814 VPWR 267.361
R1276 VPWR VPWR.t4473 267.361
R1277 VPWR.t50 VPWR 267.361
R1278 VPWR.t41 VPWR.t2361 266.985
R1279 VPWR.t6954 VPWR.t6606 266.985
R1280 VPWR.t1667 VPWR.t3237 266.204
R1281 VPWR.t3944 VPWR.t5164 266.204
R1282 VPWR VPWR.t4047 265.046
R1283 VPWR.t2238 VPWR.t4093 263.889
R1284 VPWR.t4093 VPWR.t6877 262.731
R1285 VPWR.t707 VPWR.t3919 259.26
R1286 VPWR.t3919 VPWR.t1245 259.26
R1287 VPWR.t1245 VPWR.t1457 259.26
R1288 VPWR.t1457 VPWR.t3313 259.26
R1289 VPWR.t3313 VPWR.t3998 259.26
R1290 VPWR.t3998 VPWR.t1230 259.26
R1291 VPWR.t1230 VPWR.t1153 259.26
R1292 VPWR.t1153 VPWR.t5136 259.26
R1293 VPWR.t5136 VPWR.t6284 259.26
R1294 VPWR.t6284 VPWR.t695 259.26
R1295 VPWR.t695 VPWR.t3366 259.26
R1296 VPWR.t3366 VPWR.t442 259.26
R1297 VPWR.t442 VPWR.t6071 259.26
R1298 VPWR.t6071 VPWR.t1461 259.26
R1299 VPWR.t4470 VPWR.t375 259.26
R1300 VPWR.t375 VPWR.t5179 259.26
R1301 VPWR.t5179 VPWR.t2547 259.26
R1302 VPWR.t2547 VPWR.t5239 259.26
R1303 VPWR.t5239 VPWR.t5794 259.26
R1304 VPWR.t5794 VPWR.t5431 259.26
R1305 VPWR.t5431 VPWR.t1196 259.26
R1306 VPWR.t1196 VPWR.t3701 259.26
R1307 VPWR.t3701 VPWR.t2774 259.26
R1308 VPWR.t2774 VPWR.t5262 259.26
R1309 VPWR.t5262 VPWR.t7077 259.26
R1310 VPWR.t7077 VPWR.t6170 259.26
R1311 VPWR.t6170 VPWR.t4506 259.26
R1312 VPWR.t4506 VPWR.t3208 259.26
R1313 VPWR.t889 VPWR.t887 259.26
R1314 VPWR.t6343 VPWR.t6341 259.26
R1315 VPWR.t6635 VPWR.t1532 259.26
R1316 VPWR.t322 VPWR.t5895 259.26
R1317 VPWR.t3179 VPWR.t4316 259.26
R1318 VPWR.t6518 VPWR.t5929 259.26
R1319 VPWR.t6519 VPWR.t6517 259.26
R1320 VPWR.t4962 VPWR.t4960 259.26
R1321 VPWR.t4964 VPWR.t4958 259.26
R1322 VPWR.t5058 VPWR.t2507 259.26
R1323 VPWR.t6037 VPWR.t2508 259.26
R1324 VPWR.t5817 VPWR 259.26
R1325 VPWR.t2880 VPWR.t5620 259.26
R1326 VPWR.t2181 VPWR.t5624 259.26
R1327 VPWR.t2275 VPWR.t1101 259.26
R1328 VPWR.t934 VPWR.t5352 259.26
R1329 VPWR.t1621 VPWR.t1619 259.26
R1330 VPWR.t2990 VPWR.t4560 259.26
R1331 VPWR.t3584 VPWR.t4278 259.26
R1332 VPWR.t1865 VPWR.t5412 259.26
R1333 VPWR.t6572 VPWR.t6568 259.26
R1334 VPWR.t287 VPWR.t281 259.26
R1335 VPWR.t5254 VPWR.t5116 259.26
R1336 VPWR.t271 VPWR.t267 259.26
R1337 VPWR.t6913 VPWR.t6911 259.26
R1338 VPWR.t6919 VPWR.t6921 259.26
R1339 VPWR.t6962 VPWR.t6917 259.26
R1340 VPWR.t6957 VPWR.t3914 259.26
R1341 VPWR.t5713 VPWR.t3913 259.26
R1342 VPWR.t1399 VPWR.t2778 259.26
R1343 VPWR.t3041 VPWR.t1399 259.26
R1344 VPWR.t2752 VPWR.t3041 259.26
R1345 VPWR.t5611 VPWR.t539 259.26
R1346 VPWR.t1192 VPWR.t1627 259.26
R1347 VPWR.t5525 VPWR.t5694 259.26
R1348 VPWR.t6619 VPWR.t2646 259.26
R1349 VPWR.t6290 VPWR.t204 259.26
R1350 VPWR.t3769 VPWR.t7067 259.26
R1351 VPWR.t7067 VPWR.t4056 259.26
R1352 VPWR.t4069 VPWR.t5205 259.26
R1353 VPWR.t618 VPWR.t999 259.26
R1354 VPWR.t3144 VPWR.t618 259.26
R1355 VPWR.t5939 VPWR.t3087 259.26
R1356 VPWR.t6230 VPWR.t5939 259.26
R1357 VPWR.t738 VPWR.t6230 259.26
R1358 VPWR.t409 VPWR.t738 259.26
R1359 VPWR.t1613 VPWR.t5688 259.26
R1360 VPWR.t5941 VPWR.t1613 259.26
R1361 VPWR.t5406 VPWR.t2263 259.26
R1362 VPWR.t2762 VPWR.t5223 259.26
R1363 VPWR.t991 VPWR.t2762 259.26
R1364 VPWR.t4704 VPWR.t991 259.26
R1365 VPWR.t5229 VPWR.t4838 259.26
R1366 VPWR.t5891 VPWR.t5229 259.26
R1367 VPWR.t7121 VPWR.t5891 259.26
R1368 VPWR.t1480 VPWR.t7121 259.26
R1369 VPWR.t3331 VPWR.t1480 259.26
R1370 VPWR.t5728 VPWR.t3331 259.26
R1371 VPWR.t4456 VPWR.t5728 259.26
R1372 VPWR.t811 VPWR.t4456 259.26
R1373 VPWR.t4634 VPWR.t811 259.26
R1374 VPWR.t4916 VPWR.t4634 259.26
R1375 VPWR.t3026 VPWR.t4916 259.26
R1376 VPWR.t5149 VPWR.t3026 259.26
R1377 VPWR.t385 VPWR.t5149 259.26
R1378 VPWR.t3414 VPWR.t385 259.26
R1379 VPWR.t2475 VPWR.t3414 259.26
R1380 VPWR.t2644 VPWR.t2925 259.26
R1381 VPWR.t4318 VPWR.t2644 259.26
R1382 VPWR.t1415 VPWR.t4318 259.26
R1383 VPWR.t2433 VPWR.t1415 259.26
R1384 VPWR.t5041 VPWR.t2433 259.26
R1385 VPWR.t3718 VPWR.t5041 259.26
R1386 VPWR.t2844 VPWR.t3718 259.26
R1387 VPWR.t2052 VPWR.t2844 259.26
R1388 VPWR.t827 VPWR.t2052 259.26
R1389 VPWR.t2711 VPWR.t827 259.26
R1390 VPWR.t1304 VPWR.t2711 259.26
R1391 VPWR.t2373 VPWR.t1304 259.26
R1392 VPWR.t5382 VPWR.t2373 259.26
R1393 VPWR.t2632 VPWR.t5382 259.26
R1394 VPWR.t1649 VPWR.t3652 259.26
R1395 VPWR.t610 VPWR.t1649 259.26
R1396 VPWR.t3884 VPWR.t610 259.26
R1397 VPWR.t4393 VPWR.t3884 259.26
R1398 VPWR.t5772 VPWR.t4393 259.26
R1399 VPWR.t4924 VPWR.t5772 259.26
R1400 VPWR.t1565 VPWR.t4924 259.26
R1401 VPWR.t2846 VPWR.t1565 259.26
R1402 VPWR.t5068 VPWR.t2846 259.26
R1403 VPWR.t1533 VPWR.t5068 259.26
R1404 VPWR.t5376 VPWR.t1533 259.26
R1405 VPWR.t3705 VPWR.t5376 259.26
R1406 VPWR.t1966 VPWR.t3705 259.26
R1407 VPWR.t5104 VPWR.t1966 259.26
R1408 VPWR.t3397 VPWR.t2377 259.26
R1409 VPWR.t3200 VPWR 259.26
R1410 VPWR.t735 VPWR.t4723 259.26
R1411 VPWR.t3990 VPWR.t5337 259.26
R1412 VPWR.t219 VPWR.t1185 259.26
R1413 VPWR.t1921 VPWR.t1907 259.26
R1414 VPWR.t2462 VPWR.t3081 259.26
R1415 VPWR.t7034 VPWR.t197 259.26
R1416 VPWR.t3801 VPWR.t4823 259.26
R1417 VPWR.t4808 VPWR.t1372 259.26
R1418 VPWR.t5007 VPWR.t4808 259.26
R1419 VPWR.t4578 VPWR.t5007 259.26
R1420 VPWR.t5114 VPWR.t2863 259.26
R1421 VPWR.t5490 VPWR.t2857 259.26
R1422 VPWR.t5295 VPWR.t5287 259.26
R1423 VPWR.t5287 VPWR.t3342 259.26
R1424 VPWR.t3894 VPWR.t772 259.26
R1425 VPWR.t772 VPWR.t306 259.26
R1426 VPWR.t306 VPWR.t5032 259.26
R1427 VPWR.t5032 VPWR.t6147 259.26
R1428 VPWR.t2198 VPWR.t4488 259.26
R1429 VPWR.t2115 VPWR.t2198 259.26
R1430 VPWR.t833 VPWR.t2812 259.26
R1431 VPWR.t711 VPWR.t833 259.26
R1432 VPWR.t377 VPWR.t711 259.26
R1433 VPWR.t4552 VPWR.t377 259.26
R1434 VPWR.t5967 VPWR.t4552 259.26
R1435 VPWR.t5761 VPWR.t5967 259.26
R1436 VPWR.t854 VPWR.t4771 259.26
R1437 VPWR.t768 VPWR.t4175 259.26
R1438 VPWR.t2062 VPWR.t768 259.26
R1439 VPWR.t3654 VPWR.t2062 259.26
R1440 VPWR.t3083 VPWR.t3654 259.26
R1441 VPWR.t4618 VPWR.t1375 259.26
R1442 VPWR.t1375 VPWR.t4439 259.26
R1443 VPWR.t4439 VPWR.t5329 259.26
R1444 VPWR.t5329 VPWR.t3904 259.26
R1445 VPWR.t3904 VPWR.t4165 259.26
R1446 VPWR.t4165 VPWR.t4948 259.26
R1447 VPWR.t4948 VPWR.t4103 259.26
R1448 VPWR.t4103 VPWR.t531 259.26
R1449 VPWR.t6203 VPWR.t1779 259.26
R1450 VPWR.t2054 VPWR.t6203 259.26
R1451 VPWR.t4762 VPWR.t2054 259.26
R1452 VPWR.t6250 VPWR.t4762 259.26
R1453 VPWR.t5829 VPWR.t6250 259.26
R1454 VPWR.t3164 VPWR.t5829 259.26
R1455 VPWR.t6092 VPWR.t3164 259.26
R1456 VPWR.t4912 VPWR.t6092 259.26
R1457 VPWR.t2612 VPWR.t4912 259.26
R1458 VPWR.t3876 VPWR.t2612 259.26
R1459 VPWR.t3874 VPWR.t3876 259.26
R1460 VPWR.t4020 VPWR.t3874 259.26
R1461 VPWR.t5866 VPWR.t4020 259.26
R1462 VPWR.t4638 VPWR.t5866 259.26
R1463 VPWR.t4415 VPWR.t4638 259.26
R1464 VPWR.t3242 VPWR.t629 259.26
R1465 VPWR.t3592 VPWR.t4752 259.26
R1466 VPWR.t2068 VPWR.t3592 259.26
R1467 VPWR.t2242 VPWR.t1842 259.26
R1468 VPWR.t2267 VPWR.t2242 259.26
R1469 VPWR.t4737 VPWR.t2267 259.26
R1470 VPWR.t1017 VPWR.t4737 259.26
R1471 VPWR.t419 VPWR.t1017 259.26
R1472 VPWR.t1991 VPWR.t419 259.26
R1473 VPWR.t1633 VPWR.t1991 259.26
R1474 VPWR.t1095 VPWR.t1633 259.26
R1475 VPWR.t3519 VPWR.t1095 259.26
R1476 VPWR.t3024 VPWR.t3519 259.26
R1477 VPWR.t1983 VPWR.t3329 259.26
R1478 VPWR.t3329 VPWR.t635 259.26
R1479 VPWR.t635 VPWR.t4812 259.26
R1480 VPWR.t4812 VPWR.t395 259.26
R1481 VPWR.t395 VPWR.t5440 259.26
R1482 VPWR.t5440 VPWR.t4774 259.26
R1483 VPWR.t4774 VPWR.t852 259.26
R1484 VPWR.t852 VPWR.t1557 259.26
R1485 VPWR.t1557 VPWR.t5233 259.26
R1486 VPWR.t5233 VPWR.t1811 259.26
R1487 VPWR.t1811 VPWR.t616 259.26
R1488 VPWR.t616 VPWR.t4750 259.26
R1489 VPWR.t4750 VPWR.t4781 259.26
R1490 VPWR.t4781 VPWR.t5227 259.26
R1491 VPWR.t5227 VPWR.t6079 259.26
R1492 VPWR.t3936 VPWR.t1173 259.26
R1493 VPWR.t2037 VPWR.t1877 259.26
R1494 VPWR.t6090 VPWR.t2037 259.26
R1495 VPWR.t6431 VPWR.t6090 259.26
R1496 VPWR.t5745 VPWR.t6431 259.26
R1497 VPWR.t7138 VPWR.t5745 259.26
R1498 VPWR.t5471 VPWR.t7138 259.26
R1499 VPWR.t4026 VPWR.t5471 259.26
R1500 VPWR.t6256 VPWR.t4026 259.26
R1501 VPWR.t5696 VPWR.t6256 259.26
R1502 VPWR.t1302 VPWR.t5696 259.26
R1503 VPWR.t1661 VPWR.t1302 259.26
R1504 VPWR.t1804 VPWR.t1661 259.26
R1505 VPWR.t956 VPWR.t6022 259.26
R1506 VPWR.t3958 VPWR.t956 259.26
R1507 VPWR.t367 VPWR.t3958 259.26
R1508 VPWR.t5457 VPWR.t367 259.26
R1509 VPWR.t3552 VPWR.t5457 259.26
R1510 VPWR.t1869 VPWR.t3552 259.26
R1511 VPWR.t5685 VPWR.t1869 259.26
R1512 VPWR.t5102 VPWR.t5685 259.26
R1513 VPWR.t5477 VPWR.t5102 259.26
R1514 VPWR.t4215 VPWR.t5477 259.26
R1515 VPWR.t6224 VPWR.t4215 259.26
R1516 VPWR.t6266 VPWR.t6224 259.26
R1517 VPWR.t1042 VPWR.t6266 259.26
R1518 VPWR.t466 VPWR.t1042 259.26
R1519 VPWR.t5363 VPWR.t466 259.26
R1520 VPWR.t4555 VPWR.t4744 259.26
R1521 VPWR.t5225 VPWR.t4555 259.26
R1522 VPWR.t6123 VPWR.t5225 259.26
R1523 VPWR.t1541 VPWR.t6123 259.26
R1524 VPWR.t4140 VPWR.t1541 259.26
R1525 VPWR.t4291 VPWR.t4140 259.26
R1526 VPWR.t4778 VPWR.t4291 259.26
R1527 VPWR.t3517 VPWR.t4778 259.26
R1528 VPWR.t4734 VPWR.t3517 259.26
R1529 VPWR.t4922 VPWR.t4734 259.26
R1530 VPWR.t454 VPWR.t4922 259.26
R1531 VPWR.t4349 VPWR.t454 259.26
R1532 VPWR.t2682 VPWR.t4349 259.26
R1533 VPWR.t1819 VPWR.t2682 259.26
R1534 VPWR.t4502 VPWR.t6205 259.26
R1535 VPWR.t5842 VPWR.t4502 259.26
R1536 VPWR.t813 VPWR.t5842 259.26
R1537 VPWR.t3525 VPWR.t813 259.26
R1538 VPWR.t431 VPWR.t3525 259.26
R1539 VPWR.t344 VPWR.t431 259.26
R1540 VPWR.t4401 VPWR.t344 259.26
R1541 VPWR.t6196 VPWR.t4401 259.26
R1542 VPWR.t2789 VPWR.t6196 259.26
R1543 VPWR.t2210 VPWR.t2789 259.26
R1544 VPWR.t3694 VPWR.t2210 259.26
R1545 VPWR.t2371 VPWR.t3694 259.26
R1546 VPWR.t5079 VPWR.t2371 259.26
R1547 VPWR.t2310 VPWR.t5079 259.26
R1548 VPWR.t5016 VPWR 258.103
R1549 VPWR.t6874 VPWR 258.103
R1550 VPWR.t6044 VPWR 258.103
R1551 VPWR.t401 VPWR 258.103
R1552 VPWR.t6935 VPWR.t4978 256.945
R1553 VPWR.t4314 VPWR 256.757
R1554 VPWR.t5117 VPWR 255.787
R1555 VPWR.t462 VPWR 253.472
R1556 VPWR.t6933 VPWR.t4983 252.315
R1557 VPWR.t3360 VPWR.t6933 252.315
R1558 VPWR.t6907 VPWR.t3221 251.157
R1559 VPWR.t1292 VPWR 251.157
R1560 VPWR.t6512 VPWR.t3581 250.054
R1561 VPWR.t433 VPWR.t1932 250
R1562 VPWR.t1625 VPWR.t2979 250
R1563 VPWR.t6101 VPWR.t950 250
R1564 VPWR.t119 VPWR.t181 250
R1565 VPWR.t5460 VPWR.t525 250
R1566 VPWR.t932 VPWR.t2966 250
R1567 VPWR.t1463 VPWR.t3235 250
R1568 VPWR.t6262 VPWR.t6420 250
R1569 VPWR.t4014 VPWR.t4012 250
R1570 VPWR.t5552 VPWR.t1046 250
R1571 VPWR.t6859 VPWR 248.844
R1572 VPWR.t4819 VPWR.t3350 248.844
R1573 VPWR.t1528 VPWR.t1524 245.37
R1574 VPWR VPWR.t6612 245.37
R1575 VPWR.t6769 VPWR.t3482 245.37
R1576 VPWR.t6678 VPWR.t6741 245.37
R1577 VPWR.t2729 VPWR.t4155 245.37
R1578 VPWR.t6840 VPWR.t259 245.37
R1579 VPWR.t6832 VPWR.t263 245.37
R1580 VPWR.t6836 VPWR.t261 245.37
R1581 VPWR.t6834 VPWR.t255 245.37
R1582 VPWR.t6838 VPWR.t249 245.37
R1583 VPWR.t6844 VPWR.t243 245.37
R1584 VPWR.t5127 VPWR.t6004 245.37
R1585 VPWR.t4144 VPWR.t4606 245.37
R1586 VPWR.t6162 VPWR.t508 245.37
R1587 VPWR.t506 VPWR.t5187 245.37
R1588 VPWR.t6821 VPWR.t5665 245.37
R1589 VPWR.t4602 VPWR 244.214
R1590 VPWR.t5408 VPWR 244.214
R1591 VPWR.t6570 VPWR.n714 243.056
R1592 VPWR.t803 VPWR.n822 241.899
R1593 VPWR VPWR.t3666 241.314
R1594 VPWR VPWR.t1200 241.314
R1595 VPWR VPWR.t5386 241.314
R1596 VPWR.t2580 VPWR 241.314
R1597 VPWR.t2306 VPWR 241.314
R1598 VPWR.t2148 VPWR 241.314
R1599 VPWR VPWR.t2590 241.314
R1600 VPWR.t5303 VPWR 241.314
R1601 VPWR.t5872 VPWR 241.314
R1602 VPWR.t4123 VPWR 241.314
R1603 VPWR VPWR.t23 241.314
R1604 VPWR VPWR.t6 241.314
R1605 VPWR.t2770 VPWR 241.314
R1606 VPWR.t88 VPWR 241.314
R1607 VPWR.t1294 VPWR.t727 240.742
R1608 VPWR.t199 VPWR.t2598 240.742
R1609 VPWR.t4084 VPWR.t105 239.583
R1610 VPWR.t4330 VPWR.t4742 238.427
R1611 VPWR.n2874 VPWR.t4383 238.427
R1612 VPWR VPWR.t2571 237.269
R1613 VPWR VPWR.t7064 237.269
R1614 VPWR VPWR.t3882 237.269
R1615 VPWR.t2487 VPWR 237.269
R1616 VPWR.t3888 VPWR 237.269
R1617 VPWR.t4437 VPWR 237.269
R1618 VPWR.t1389 VPWR 237.269
R1619 VPWR VPWR.t2367 237.269
R1620 VPWR VPWR.t3174 237.269
R1621 VPWR.t2204 VPWR 237.269
R1622 VPWR.t5074 VPWR 237.269
R1623 VPWR.t6480 VPWR.t158 236.112
R1624 VPWR.t1258 VPWR.t1158 236.112
R1625 VPWR.t5670 VPWR.t413 236.112
R1626 VPWR.t6478 VPWR.t6867 236.112
R1627 VPWR.t6468 VPWR.t7056 236.112
R1628 VPWR.t6779 VPWR.t151 236.112
R1629 VPWR.t5210 VPWR.t1128 236.112
R1630 VPWR.t2659 VPWR.t2652 236.112
R1631 VPWR.t6736 VPWR.t7066 236.112
R1632 VPWR.t7065 VPWR.t3489 236.112
R1633 VPWR.t1034 VPWR.t203 236.112
R1634 VPWR.t6947 VPWR.t6750 236.112
R1635 VPWR.t3180 VPWR.t6026 236.112
R1636 VPWR.t5925 VPWR.t6522 236.112
R1637 VPWR.t2048 VPWR.t2044 236.112
R1638 VPWR.t6494 VPWR.t6905 236.112
R1639 VPWR.t6476 VPWR.t102 236.112
R1640 VPWR.t3669 VPWR.t3671 236.112
R1641 VPWR.t6410 VPWR.t6848 236.112
R1642 VPWR.t6848 VPWR.t4085 236.112
R1643 VPWR.t2557 VPWR.t4087 236.112
R1644 VPWR.t2555 VPWR.t4091 236.112
R1645 VPWR.t4089 VPWR.t1256 236.112
R1646 VPWR.t6850 VPWR.t6408 236.112
R1647 VPWR.t3468 VPWR.t6975 236.112
R1648 VPWR.t4049 VPWR.t6728 236.112
R1649 VPWR.t6638 VPWR.t4282 236.112
R1650 VPWR.t6871 VPWR.t1214 236.112
R1651 VPWR.t1428 VPWR.t1430 236.112
R1652 VPWR.t523 VPWR.t1324 236.112
R1653 VPWR.t6720 VPWR.t4222 236.112
R1654 VPWR.t3950 VPWR.t643 236.112
R1655 VPWR.t645 VPWR.t4698 236.112
R1656 VPWR.t5305 VPWR.t2447 236.112
R1657 VPWR VPWR.t1322 236.112
R1658 VPWR.t3729 VPWR.t3826 236.112
R1659 VPWR.t6466 VPWR.t6383 236.112
R1660 VPWR.t6472 VPWR.t7006 236.112
R1661 VPWR.t6484 VPWR.t6338 236.112
R1662 VPWR.t6856 VPWR.t3636 236.112
R1663 VPWR.t1873 VPWR.t789 236.112
R1664 VPWR.t336 VPWR.t4835 236.112
R1665 VPWR.t6369 VPWR.t6754 236.112
R1666 VPWR.t181 VPWR.t3308 236.112
R1667 VPWR.t2477 VPWR.t14 236.112
R1668 VPWR.t6429 VPWR.t4690 236.112
R1669 VPWR.t3477 VPWR.t480 236.112
R1670 VPWR.t2350 VPWR.t6529 236.112
R1671 VPWR.t3470 VPWR.t477 236.112
R1672 VPWR.t6985 VPWR.t4557 236.112
R1673 VPWR.t167 VPWR.t6406 236.112
R1674 VPWR.t6464 VPWR.t7027 236.112
R1675 VPWR.t169 VPWR.t6993 236.112
R1676 VPWR.t6739 VPWR.t169 236.112
R1677 VPWR.t6470 VPWR.t6388 236.112
R1678 VPWR.t6396 VPWR.t6663 236.112
R1679 VPWR.t6589 VPWR.t6888 236.112
R1680 VPWR.t2545 VPWR.t5590 236.112
R1681 VPWR.t5592 VPWR.t2539 236.112
R1682 VPWR.t4821 VPWR.t2164 236.112
R1683 VPWR.t1861 VPWR.t7025 236.112
R1684 VPWR.t4159 VPWR.t7018 236.112
R1685 VPWR.t6659 VPWR.t154 236.112
R1686 VPWR.t165 VPWR.t4205 236.112
R1687 VPWR.t4231 VPWR.t4819 236.112
R1688 VPWR.t5539 VPWR.t4472 236.112
R1689 VPWR.t267 VPWR.t1264 236.112
R1690 VPWR.t265 VPWR.t6800 236.112
R1691 VPWR.t6602 VPWR.t2378 236.112
R1692 VPWR.t25 VPWR.t6746 236.112
R1693 VPWR.t193 VPWR.t305 236.112
R1694 VPWR.t3395 VPWR.t6826 236.112
R1695 VPWR.t6426 VPWR.t6955 236.112
R1696 VPWR.t4990 VPWR.t4988 236.112
R1697 VPWR.t6890 VPWR.t5120 236.112
R1698 VPWR.t6583 VPWR.t960 236.112
R1699 VPWR.t4999 VPWR.t4326 236.112
R1700 VPWR.t6731 VPWR.t5997 236.112
R1701 VPWR.t4135 VPWR.t5155 236.112
R1702 VPWR.t6881 VPWR.t2704 236.112
R1703 VPWR.t6395 VPWR.t5446 236.112
R1704 VPWR.t6667 VPWR.t199 236.112
R1705 VPWR.t4684 VPWR.t4699 236.112
R1706 VPWR.t4462 VPWR.t300 236.112
R1707 VPWR.t136 VPWR.t4798 236.112
R1708 VPWR.t6852 VPWR 234.804
R1709 VPWR.t2744 VPWR.t7008 233.797
R1710 VPWR.t6533 VPWR.t2346 233.471
R1711 VPWR VPWR.t1520 232.639
R1712 VPWR.t5384 VPWR.t3097 231.482
R1713 VPWR.t5185 VPWR.t843 231.482
R1714 VPWR.t1314 VPWR.t444 231.482
R1715 VPWR.t1863 VPWR.t3797 231.482
R1716 VPWR.t3206 VPWR.t6460 231.482
R1717 VPWR.t7044 VPWR.t332 231.482
R1718 VPWR.t6038 VPWR.t5603 231.482
R1719 VPWR.n458 VPWR.t3112 231.482
R1720 VPWR.t4095 VPWR.t5609 231.482
R1721 VPWR.t4047 VPWR.t216 231.482
R1722 VPWR.t5782 VPWR.n372 231.482
R1723 VPWR.t2640 VPWR 230.325
R1724 VPWR VPWR.t4251 230.325
R1725 VPWR.t6153 VPWR 230.325
R1726 VPWR.t1694 VPWR 230.325
R1727 VPWR VPWR.t7037 229.167
R1728 VPWR.t3868 VPWR.t2618 229.167
R1729 VPWR.t5047 VPWR.t231 229.167
R1730 VPWR.t3577 VPWR 228.01
R1731 VPWR.t727 VPWR 228.01
R1732 VPWR.t48 VPWR.t2702 228.01
R1733 VPWR.t6829 VPWR.t3911 228.01
R1734 VPWR.t6795 VPWR.t1262 227.424
R1735 VPWR.t2951 VPWR.t6804 227.424
R1736 VPWR.t6392 VPWR.t3724 226.852
R1737 VPWR.t439 VPWR.t4463 226.852
R1738 VPWR.t3217 VPWR.t6366 225.695
R1739 VPWR VPWR.t1109 225.695
R1740 VPWR VPWR.t6564 225.695
R1741 VPWR VPWR.t6556 225.695
R1742 VPWR.t237 VPWR 225.695
R1743 VPWR.t6778 VPWR.n929 224.537
R1744 VPWR.t5437 VPWR.t3020 224.537
R1745 VPWR.t6625 VPWR.t6513 224.077
R1746 VPWR.t6623 VPWR.t6509 224.077
R1747 VPWR.t1214 VPWR.t3148 223.381
R1748 VPWR VPWR.t4689 222.885
R1749 VPWR.t6698 VPWR.t7041 222.222
R1750 VPWR.t6700 VPWR.t6492 222.222
R1751 VPWR.t1958 VPWR.t6505 222.222
R1752 VPWR.t1591 VPWR.t5737 222.222
R1753 VPWR.t776 VPWR.t116 222.222
R1754 VPWR.t3422 VPWR.t6744 222.222
R1755 VPWR.t2737 VPWR.t468 222.222
R1756 VPWR.t2837 VPWR.t2772 221.065
R1757 VPWR.t3622 VPWR.t5596 221.065
R1758 VPWR.t2457 VPWR.t2543 221.065
R1759 VPWR.t1473 VPWR.t3303 221.065
R1760 VPWR.t6713 VPWR.t4796 221.065
R1761 VPWR.t6081 VPWR 219.907
R1762 VPWR.t3658 VPWR.t6677 219.907
R1763 VPWR.t2504 VPWR.t4990 219.907
R1764 VPWR.t2735 VPWR.t1948 218.75
R1765 VPWR.t6735 VPWR.t2573 218.75
R1766 VPWR.t158 VPWR.t5062 217.594
R1767 VPWR.t6900 VPWR.t140 217.594
R1768 VPWR.t3535 VPWR.t6778 217.594
R1769 VPWR.t3533 VPWR.t149 217.594
R1770 VPWR.t5921 VPWR.t3229 217.594
R1771 VPWR.t4006 VPWR.t3228 217.594
R1772 VPWR.t5628 VPWR.t6925 217.594
R1773 VPWR.t1268 VPWR.t5488 217.594
R1774 VPWR.t6802 VPWR.t5848 217.594
R1775 VPWR.n3256 VPWR.t3658 215.279
R1776 VPWR.t1668 VPWR.t1790 215.279
R1777 VPWR.t4510 VPWR.t5909 215.279
R1778 VPWR.t4508 VPWR.t5907 215.279
R1779 VPWR.t2997 VPWR.t6131 215.279
R1780 VPWR.t2999 VPWR.t6129 215.279
R1781 VPWR.t1124 VPWR.t606 215.279
R1782 VPWR.t1126 VPWR.t608 215.279
R1783 VPWR.t1368 VPWR.t968 215.279
R1784 VPWR.t1366 VPWR.t966 215.279
R1785 VPWR.t5133 VPWR.t4651 215.279
R1786 VPWR.t5131 VPWR.t4649 215.279
R1787 VPWR.t4062 VPWR.t3573 215.279
R1788 VPWR.t4060 VPWR.t3571 215.279
R1789 VPWR.t877 VPWR.t1944 215.279
R1790 VPWR.t2869 VPWR.t1729 215.279
R1791 VPWR.t2867 VPWR.t1731 215.279
R1792 VPWR.t6239 VPWR.t3016 214.542
R1793 VPWR.t2481 VPWR.t6636 214.226
R1794 VPWR VPWR.t6037 214.12
R1795 VPWR.t1169 VPWR.t6087 214.12
R1796 VPWR.t790 VPWR.t5212 214.12
R1797 VPWR.t1777 VPWR.t6367 212.964
R1798 VPWR.t797 VPWR.t2029 212.964
R1799 VPWR.t7000 VPWR.t6792 212.964
R1800 VPWR.t12 VPWR.t1021 212.964
R1801 VPWR.t2783 VPWR.t5911 212.964
R1802 VPWR.t440 VPWR.t6806 212.964
R1803 VPWR.t131 VPWR.t5001 212.964
R1804 VPWR.t4795 VPWR.t4800 212.964
R1805 VPWR.t3610 VPWR.t5153 212.964
R1806 VPWR.t4527 VPWR.t165 210.649
R1807 VPWR.t6742 VPWR.t20 209.774
R1808 VPWR.t6752 VPWR.t6503 209.774
R1809 VPWR VPWR.t3805 209.492
R1810 VPWR.t1210 VPWR 209.492
R1811 VPWR VPWR.t1333 209.492
R1812 VPWR.t5523 VPWR 209.492
R1813 VPWR VPWR.t7129 209.492
R1814 VPWR.t2387 VPWR 209.492
R1815 VPWR VPWR.t4702 209.492
R1816 VPWR.t2111 VPWR 209.492
R1817 VPWR VPWR.t1522 209.492
R1818 VPWR.t2671 VPWR 209.492
R1819 VPWR VPWR.t7073 209.492
R1820 VPWR.t2787 VPWR 209.492
R1821 VPWR VPWR.t4419 209.492
R1822 VPWR.t2329 VPWR 209.492
R1823 VPWR VPWR.t2188 209.492
R1824 VPWR.t4972 VPWR 209.492
R1825 VPWR VPWR.t516 209.492
R1826 VPWR.t1733 VPWR 209.492
R1827 VPWR VPWR.t5466 209.492
R1828 VPWR.t2742 VPWR 209.492
R1829 VPWR VPWR.t1623 209.492
R1830 VPWR.t7101 VPWR 209.492
R1831 VPWR VPWR.t1306 209.492
R1832 VPWR.t2785 VPWR 209.492
R1833 VPWR VPWR.t3215 209.492
R1834 VPWR.t3924 VPWR 209.492
R1835 VPWR VPWR.t3603 209.492
R1836 VPWR.t80 VPWR 209.492
R1837 VPWR VPWR.t4217 209.492
R1838 VPWR.t3722 VPWR 209.492
R1839 VPWR VPWR.t3837 209.492
R1840 VPWR.t4346 VPWR 209.492
R1841 VPWR VPWR.n101 209.492
R1842 VPWR VPWR.n99 209.492
R1843 VPWR VPWR.n97 209.492
R1844 VPWR.t4494 VPWR 209.492
R1845 VPWR.n965 VPWR 209.492
R1846 VPWR.n947 VPWR 209.492
R1847 VPWR.n938 VPWR 209.492
R1848 VPWR VPWR.n1038 209.492
R1849 VPWR VPWR.n912 209.492
R1850 VPWR.n3355 VPWR 209.492
R1851 VPWR.n853 VPWR 209.492
R1852 VPWR VPWR.n1276 209.492
R1853 VPWR.t1825 VPWR.t7011 209.492
R1854 VPWR.t2050 VPWR.t5058 209.492
R1855 VPWR.t4523 VPWR 209.492
R1856 VPWR.t5658 VPWR 209.492
R1857 VPWR.n1278 VPWR 209.492
R1858 VPWR.t4468 VPWR 209.492
R1859 VPWR.t4468 VPWR 209.492
R1860 VPWR.t4610 VPWR 209.492
R1861 VPWR VPWR.t5803 209.492
R1862 VPWR VPWR.n819 209.492
R1863 VPWR.n822 VPWR 209.492
R1864 VPWR.t5705 VPWR 209.492
R1865 VPWR.t3192 VPWR 209.492
R1866 VPWR.t2427 VPWR 209.492
R1867 VPWR.t3906 VPWR 209.492
R1868 VPWR.t5515 VPWR 209.492
R1869 VPWR VPWR.t6258 209.492
R1870 VPWR.t4714 VPWR 209.492
R1871 VPWR.t3202 VPWR 209.492
R1872 VPWR.t2793 VPWR 209.492
R1873 VPWR.n143 VPWR 209.492
R1874 VPWR VPWR.n136 209.492
R1875 VPWR.n1175 VPWR 209.492
R1876 VPWR VPWR.n724 209.492
R1877 VPWR VPWR.n1778 209.492
R1878 VPWR.t1950 VPWR 209.492
R1879 VPWR.t2479 VPWR 209.492
R1880 VPWR.t4340 VPWR 209.492
R1881 VPWR VPWR.t3271 209.492
R1882 VPWR VPWR.t5574 209.492
R1883 VPWR.t5099 VPWR 209.492
R1884 VPWR.t5833 VPWR 209.492
R1885 VPWR.n628 VPWR 209.492
R1886 VPWR.t3590 VPWR 209.492
R1887 VPWR.t3495 VPWR 209.492
R1888 VPWR.n1087 VPWR 209.492
R1889 VPWR.t764 VPWR 209.492
R1890 VPWR.t5024 VPWR 209.492
R1891 VPWR.t5800 VPWR 209.492
R1892 VPWR.t3850 VPWR 209.492
R1893 VPWR.t1260 VPWR 209.492
R1894 VPWR.t6077 VPWR 209.492
R1895 VPWR.n1936 VPWR 209.492
R1896 VPWR.t5420 VPWR 209.492
R1897 VPWR.t2019 VPWR 209.492
R1898 VPWR VPWR.t3624 209.492
R1899 VPWR VPWR.t1792 209.492
R1900 VPWR.t562 VPWR 209.492
R1901 VPWR.t4045 VPWR 209.492
R1902 VPWR VPWR.t5162 209.492
R1903 VPWR VPWR.t5768 209.492
R1904 VPWR VPWR.t6179 209.492
R1905 VPWR VPWR.t496 209.492
R1906 VPWR VPWR.t2714 209.492
R1907 VPWR.t427 VPWR 209.492
R1908 VPWR.t3617 VPWR 209.492
R1909 VPWR VPWR.t3317 209.492
R1910 VPWR VPWR.t3190 209.492
R1911 VPWR.t5541 VPWR 209.492
R1912 VPWR.t3626 VPWR 209.492
R1913 VPWR.t4525 VPWR 209.492
R1914 VPWR.t1561 VPWR 209.492
R1915 VPWR.t6201 VPWR 209.492
R1916 VPWR.t3523 VPWR 209.492
R1917 VPWR.t3642 VPWR 209.492
R1918 VPWR.t3550 VPWR 209.492
R1919 VPWR.t2449 VPWR 209.492
R1920 VPWR.t5107 VPWR 209.492
R1921 VPWR.t1247 VPWR 209.492
R1922 VPWR.t5555 VPWR 209.492
R1923 VPWR.t547 VPWR 209.492
R1924 VPWR.n2325 VPWR 209.492
R1925 VPWR.t3393 VPWR 209.492
R1926 VPWR.t4933 VPWR 209.492
R1927 VPWR.t2776 VPWR 209.492
R1928 VPWR.t3391 VPWR 209.492
R1929 VPWR.t1040 VPWR 209.492
R1930 VPWR.t5367 VPWR 209.492
R1931 VPWR VPWR.t3389 209.492
R1932 VPWR VPWR.t3795 209.492
R1933 VPWR.t7131 VPWR 209.492
R1934 VPWR.t2718 VPWR 209.492
R1935 VPWR.t4336 VPWR 209.492
R1936 VPWR.t2312 VPWR 209.492
R1937 VPWR.n2066 VPWR 209.492
R1938 VPWR.t5849 VPWR 209.492
R1939 VPWR.n200 VPWR 209.492
R1940 VPWR.n202 VPWR 209.492
R1941 VPWR.n204 VPWR 209.492
R1942 VPWR.n206 VPWR 209.492
R1943 VPWR VPWR.t3727 209.492
R1944 VPWR VPWR.t6301 209.492
R1945 VPWR.t2136 VPWR 209.492
R1946 VPWR.t2025 VPWR 209.492
R1947 VPWR.t3210 VPWR 209.492
R1948 VPWR.t2375 VPWR 209.492
R1949 VPWR.n535 VPWR 209.492
R1950 VPWR.t6418 VPWR.t5823 209.492
R1951 VPWR.n541 VPWR 209.492
R1952 VPWR VPWR.t5796 209.492
R1953 VPWR VPWR.n176 209.492
R1954 VPWR VPWR.n525 209.492
R1955 VPWR.t6133 VPWR 209.492
R1956 VPWR.t4500 VPWR 209.492
R1957 VPWR VPWR.t885 209.492
R1958 VPWR.n395 VPWR 209.492
R1959 VPWR.t2253 VPWR 209.492
R1960 VPWR.t1575 VPWR 209.492
R1961 VPWR.t5666 VPWR 209.492
R1962 VPWR.t1719 VPWR 209.492
R1963 VPWR VPWR.n374 209.492
R1964 VPWR.t5235 VPWR 209.492
R1965 VPWR VPWR.n267 209.492
R1966 VPWR.n2428 VPWR 209.492
R1967 VPWR VPWR.n262 209.492
R1968 VPWR.n2535 VPWR 209.492
R1969 VPWR.n2537 VPWR 209.492
R1970 VPWR.n2539 VPWR 209.492
R1971 VPWR.n2541 VPWR 209.492
R1972 VPWR.n10 VPWR 209.492
R1973 VPWR.n32 VPWR 209.492
R1974 VPWR.n34 VPWR 209.492
R1975 VPWR.n64 VPWR 209.492
R1976 VPWR.n85 VPWR 209.492
R1977 VPWR.n87 VPWR 209.492
R1978 VPWR.t6333 VPWR.t670 208.333
R1979 VPWR.t2562 VPWR.t6402 208.333
R1980 VPWR.t3631 VPWR.t3373 208.333
R1981 VPWR.t4107 VPWR.t4569 208.333
R1982 VPWR.t6552 VPWR.t4908 208.333
R1983 VPWR.t527 VPWR.t6373 208.333
R1984 VPWR.t6925 VPWR.t3731 208.333
R1985 VPWR.t4383 VPWR.t5565 208.333
R1986 VPWR.t5730 VPWR.t3579 207.177
R1987 VPWR VPWR.t3708 207.177
R1988 VPWR VPWR.t3878 207.177
R1989 VPWR VPWR.t3584 207.177
R1990 VPWR VPWR.t1268 207.177
R1991 VPWR.t1601 VPWR 207.177
R1992 VPWR.t1120 VPWR 207.177
R1993 VPWR VPWR.t1725 207.177
R1994 VPWR VPWR.t3990 207.177
R1995 VPWR.n3255 VPWR.t6966 206.019
R1996 VPWR.t3575 VPWR 204.862
R1997 VPWR.t6578 VPWR 204.633
R1998 VPWR VPWR.t6903 204.633
R1999 VPWR.t1381 VPWR 204.633
R2000 VPWR.t320 VPWR 204.633
R2001 VPWR.t1220 VPWR 204.633
R2002 VPWR.t2291 VPWR 204.633
R2003 VPWR.t2227 VPWR.t2519 203.704
R2004 VPWR.t3279 VPWR.t1942 203.704
R2005 VPWR.t918 VPWR.t4866 203.704
R2006 VPWR.t7103 VPWR.t4479 203.704
R2007 VPWR.t4481 VPWR.t6172 203.704
R2008 VPWR.t902 VPWR.t1079 203.704
R2009 VPWR.t2727 VPWR.t4157 203.704
R2010 VPWR.t3310 VPWR.t6544 203.704
R2011 VPWR.t6981 VPWR.t6548 203.704
R2012 VPWR.t6428 VPWR.t5563 203.704
R2013 VPWR VPWR.t5931 202.703
R2014 VPWR.t5927 VPWR 202.703
R2015 VPWR VPWR.t3559 202.703
R2016 VPWR.t45 VPWR 202.703
R2017 VPWR.t108 VPWR 202.703
R2018 VPWR VPWR.t5831 202.703
R2019 VPWR.t6672 VPWR 202.703
R2020 VPWR.t1737 VPWR 202.703
R2021 VPWR VPWR.t7052 202.703
R2022 VPWR.t6764 VPWR 202.703
R2023 VPWR VPWR.t3355 202.703
R2024 VPWR.t8 VPWR 202.703
R2025 VPWR VPWR.t6748 202.703
R2026 VPWR VPWR.t6690 202.547
R2027 VPWR.t1472 VPWR.t896 202.547
R2028 VPWR.t6711 VPWR.t4791 202.547
R2029 VPWR.n954 VPWR.t6680 201.389
R2030 VPWR.t6867 VPWR.t889 201.389
R2031 VPWR.t4870 VPWR.n1035 201.389
R2032 VPWR.t3474 VPWR.t2359 201.389
R2033 VPWR.t5869 VPWR.t3140 201.389
R2034 VPWR.t817 VPWR.t5092 201.389
R2035 VPWR.t4302 VPWR.t91 201.389
R2036 VPWR.t163 VPWR.t3011 201.389
R2037 VPWR.t98 VPWR.t5763 201.389
R2038 VPWR.t6958 VPWR.t227 201.389
R2039 VPWR.t4849 VPWR.t6823 201.389
R2040 VPWR.t6508 VPWR.t2027 200.238
R2041 VPWR VPWR.t3295 200.232
R2042 VPWR.t4514 VPWR.t5777 199.075
R2043 VPWR.t314 VPWR.t3833 199.075
R2044 VPWR.t4655 VPWR.t6787 199.075
R2045 VPWR.t612 VPWR.t2227 199.075
R2046 VPWR.t3045 VPWR.t3255 199.075
R2047 VPWR.t1796 VPWR.t5569 199.075
R2048 VPWR.t5146 VPWR.t6377 199.075
R2049 VPWR.t3570 VPWR.t5594 197.917
R2050 VPWR.t4237 VPWR.t3305 197.917
R2051 VPWR.t3671 VPWR.t1599 196.76
R2052 VPWR.t2378 VPWR.n624 196.76
R2053 VPWR.t3140 VPWR 195.602
R2054 VPWR.t3142 VPWR 195.602
R2055 VPWR.t6125 VPWR.t7098 195.602
R2056 VPWR.t2174 VPWR.t6385 195.602
R2057 VPWR.t161 VPWR.t3821 195.602
R2058 VPWR.t100 VPWR.t4717 195.602
R2059 VPWR.t6682 VPWR.t1690 194.445
R2060 VPWR.t15 VPWR.t7035 194.445
R2061 VPWR.t2959 VPWR.t3631 194.445
R2062 VPWR.t4569 VPWR.t4105 194.445
R2063 VPWR.t3476 VPWR.t6540 194.445
R2064 VPWR.t6107 VPWR.t3344 194.445
R2065 VPWR VPWR.t6694 193.287
R2066 VPWR.t5632 VPWR.t3729 193.287
R2067 VPWR.t3623 VPWR.t2545 193.287
R2068 VPWR.t3569 VPWR.t2537 193.287
R2069 VPWR VPWR.t279 193.287
R2070 VPWR.t6931 VPWR 193.287
R2071 VPWR.t2559 VPWR.t5231 192.131
R2072 VPWR.t7062 VPWR.n1392 192.131
R2073 VPWR.t2560 VPWR.n115 192.131
R2074 VPWR.n3269 VPWR.t1337 192.131
R2075 VPWR.t6909 VPWR.t4980 192.131
R2076 VPWR.t6611 VPWR.t6819 191.895
R2077 VPWR.t6949 VPWR 191.895
R2078 VPWR.t5257 VPWR 190.972
R2079 VPWR.t6046 VPWR.t411 189.815
R2080 VPWR.t6964 VPWR.t2085 189.815
R2081 VPWR.t3934 VPWR.t6035 189.815
R2082 VPWR.t1595 VPWR 188.657
R2083 VPWR.t942 VPWR 188.657
R2084 VPWR.n920 VPWR.t5921 187.5
R2085 VPWR.t6905 VPWR.t5544 187.5
R2086 VPWR.t6808 VPWR.t5397 187.5
R2087 VPWR.t4079 VPWR.t6369 187.5
R2088 VPWR.t7027 VPWR.t6363 187.5
R2089 VPWR.t1785 VPWR.t6424 187.5
R2090 VPWR.t3899 VPWR.t6601 187.5
R2091 VPWR.n612 VPWR.t265 187.5
R2092 VPWR.t6939 VPWR.t4981 187.5
R2093 VPWR.t3361 VPWR.t6937 187.5
R2094 VPWR.t2533 VPWR.t25 187.5
R2095 VPWR.t1792 VPWR.t193 187.5
R2096 VPWR.t204 VPWR.t977 187.5
R2097 VPWR.t7115 VPWR.t4550 187.5
R2098 VPWR.t4665 VPWR.t1517 187.5
R2099 VPWR.t5046 VPWR.t229 187.5
R2100 VPWR.t2377 VPWR.n535 187.5
R2101 VPWR.t3346 VPWR.t2196 187.5
R2102 VPWR.t4661 VPWR.t4802 187.5
R2103 VPWR.n371 VPWR.t3462 187.5
R2104 VPWR.t2874 VPWR.t3120 187.5
R2105 VPWR VPWR.t1030 186.344
R2106 VPWR.t1881 VPWR.n1400 186.344
R2107 VPWR.t3752 VPWR.t5442 186.344
R2108 VPWR VPWR.t1155 186.344
R2109 VPWR.t6346 VPWR.t958 186.344
R2110 VPWR.t1928 VPWR.t3219 185.936
R2111 VPWR.t3001 VPWR.t6979 185.797
R2112 VPWR.t138 VPWR.t6896 185.185
R2113 VPWR.t4996 VPWR.t43 185.185
R2114 VPWR.t5896 VPWR.t6216 185.185
R2115 VPWR.t2654 VPWR.t3750 185.185
R2116 VPWR.t4937 VPWR.t6335 185.185
R2117 VPWR.t4521 VPWR.t1411 185.185
R2118 VPWR.t5357 VPWR.t6991 185.185
R2119 VPWR.t6554 VPWR.t3311 185.185
R2120 VPWR.t251 VPWR.t122 185.185
R2121 VPWR.t245 VPWR.t6507 185.185
R2122 VPWR.t5827 VPWR.t5782 185.185
R2123 VPWR VPWR.t970 184.029
R2124 VPWR VPWR.t2562 184.029
R2125 VPWR.t6575 VPWR 184.029
R2126 VPWR.t6774 VPWR.t3575 184.029
R2127 VPWR VPWR.t6986 184.029
R2128 VPWR VPWR.t440 184.029
R2129 VPWR.t6029 VPWR 184.029
R2130 VPWR VPWR.t898 184.029
R2131 VPWR.t4320 VPWR.t4324 184.029
R2132 VPWR.t3297 VPWR.t3299 184.029
R2133 VPWR.n935 VPWR.t3291 182.87
R2134 VPWR.t6677 VPWR.t948 182.87
R2135 VPWR.t1665 VPWR.t4876 182.87
R2136 VPWR.n2866 VPWR.t588 182.87
R2137 VPWR.t5276 VPWR.t1328 182.87
R2138 VPWR.t1467 VPWR.t5221 182.87
R2139 VPWR.t5887 VPWR 181.714
R2140 VPWR VPWR.t4496 181.714
R2141 VPWR.t2602 VPWR 181.714
R2142 VPWR.t6531 VPWR.t6613 181.168
R2143 VPWR.t4036 VPWR.t4397 180.556
R2144 VPWR.t6790 VPWR.t3529 180.556
R2145 VPWR.t614 VPWR.t3413 180.556
R2146 VPWR.t5487 VPWR.t5807 180.556
R2147 VPWR.t1519 VPWR.t6305 180.556
R2148 VPWR.t5617 VPWR.t407 180.556
R2149 VPWR.t2261 VPWR.t3285 180.556
R2150 VPWR.t6008 VPWR.t3371 180.556
R2151 VPWR.t4109 VPWR.t6296 180.556
R2152 VPWR.t3264 VPWR.t817 180.556
R2153 VPWR.t172 VPWR.t4207 180.556
R2154 VPWR.t6984 VPWR.t4211 180.556
R2155 VPWR.t6319 VPWR.t2781 180.556
R2156 VPWR.t4837 VPWR.t3130 180.556
R2157 VPWR.t898 VPWR.t6029 180.556
R2158 VPWR.t5250 VPWR.t5011 180.556
R2159 VPWR.t3253 VPWR.t3944 180.556
R2160 VPWR.t2076 VPWR.t1905 180.556
R2161 VPWR.t2597 VPWR.t1923 180.556
R2162 VPWR.t3978 VPWR 179.399
R2163 VPWR VPWR.t1210 179.399
R2164 VPWR VPWR.t697 179.399
R2165 VPWR.t1997 VPWR 179.399
R2166 VPWR VPWR.t5523 179.399
R2167 VPWR VPWR.t2281 179.399
R2168 VPWR.t429 VPWR 179.399
R2169 VPWR VPWR.t2387 179.399
R2170 VPWR VPWR.t1013 179.399
R2171 VPWR.t3286 VPWR 179.399
R2172 VPWR VPWR.t2111 179.399
R2173 VPWR VPWR.t1899 179.399
R2174 VPWR.t1835 VPWR 179.399
R2175 VPWR VPWR.t2671 179.399
R2176 VPWR VPWR.t328 179.399
R2177 VPWR.t1135 VPWR 179.399
R2178 VPWR VPWR.t2787 179.399
R2179 VPWR VPWR.t3540 179.399
R2180 VPWR.t3650 VPWR 179.399
R2181 VPWR VPWR.t2329 179.399
R2182 VPWR VPWR.t68 179.399
R2183 VPWR.t2849 VPWR 179.399
R2184 VPWR VPWR.t4972 179.399
R2185 VPWR VPWR.t1061 179.399
R2186 VPWR.t5369 VPWR 179.399
R2187 VPWR VPWR.t1733 179.399
R2188 VPWR VPWR.t3340 179.399
R2189 VPWR.t5289 VPWR 179.399
R2190 VPWR VPWR.t2742 179.399
R2191 VPWR VPWR.t2109 179.399
R2192 VPWR.t6067 VPWR 179.399
R2193 VPWR VPWR.t7101 179.399
R2194 VPWR VPWR.t4583 179.399
R2195 VPWR.t4785 VPWR 179.399
R2196 VPWR VPWR.t2785 179.399
R2197 VPWR VPWR.t3594 179.399
R2198 VPWR.t4115 VPWR 179.399
R2199 VPWR VPWR.t3924 179.399
R2200 VPWR VPWR.t4883 179.399
R2201 VPWR.t5313 VPWR 179.399
R2202 VPWR VPWR.t80 179.399
R2203 VPWR VPWR.t482 179.399
R2204 VPWR.t3720 VPWR 179.399
R2205 VPWR VPWR.t3722 179.399
R2206 VPWR VPWR.t2610 179.399
R2207 VPWR.t2168 VPWR 179.399
R2208 VPWR VPWR.t4346 179.399
R2209 VPWR VPWR.t1757 179.399
R2210 VPWR.t3074 VPWR 179.399
R2211 VPWR.t2403 VPWR 179.399
R2212 VPWR.t5416 VPWR 179.399
R2213 VPWR.t1916 VPWR 179.399
R2214 VPWR.t1461 VPWR 179.399
R2215 VPWR.t6442 VPWR 179.399
R2216 VPWR.t3208 VPWR 179.399
R2217 VPWR VPWR.t86 179.399
R2218 VPWR VPWR.n955 179.399
R2219 VPWR VPWR.t4399 179.399
R2220 VPWR.t5656 VPWR 179.399
R2221 VPWR VPWR.n1386 179.399
R2222 VPWR VPWR.t4272 179.399
R2223 VPWR VPWR.n1389 179.399
R2224 VPWR VPWR.t633 179.399
R2225 VPWR VPWR.t4177 179.399
R2226 VPWR VPWR.n3354 179.399
R2227 VPWR VPWR.t3449 179.399
R2228 VPWR.t881 VPWR 179.399
R2229 VPWR VPWR.t5355 179.399
R2230 VPWR VPWR.t6024 179.399
R2231 VPWR VPWR.t2050 179.399
R2232 VPWR VPWR.t5056 179.399
R2233 VPWR VPWR.t3456 179.399
R2234 VPWR VPWR.t1149 179.399
R2235 VPWR VPWR.t5214 179.399
R2236 VPWR VPWR.t1936 179.399
R2237 VPWR VPWR.t6260 179.399
R2238 VPWR VPWR.t2419 179.399
R2239 VPWR VPWR.t4234 179.399
R2240 VPWR VPWR.n1229 179.399
R2241 VPWR VPWR.t1875 179.399
R2242 VPWR.t3906 VPWR 179.399
R2243 VPWR.t5352 VPWR 179.399
R2244 VPWR.t715 VPWR 179.399
R2245 VPWR.t5468 VPWR 179.399
R2246 VPWR.t922 VPWR 179.399
R2247 VPWR VPWR.t4567 179.399
R2248 VPWR VPWR.t4079 179.399
R2249 VPWR VPWR.t3683 179.399
R2250 VPWR.t3170 VPWR 179.399
R2251 VPWR.t397 VPWR 179.399
R2252 VPWR.t928 VPWR 179.399
R2253 VPWR.t3357 VPWR 179.399
R2254 VPWR VPWR.t1882 179.399
R2255 VPWR VPWR.t4994 179.399
R2256 VPWR VPWR.t2245 179.399
R2257 VPWR VPWR.t664 179.399
R2258 VPWR VPWR.t2793 179.399
R2259 VPWR VPWR.t3600 179.399
R2260 VPWR VPWR.t354 179.399
R2261 VPWR.t6291 VPWR.t6990 179.399
R2262 VPWR VPWR.t1635 179.399
R2263 VPWR.t4876 VPWR 179.399
R2264 VPWR.n1783 VPWR 179.399
R2265 VPWR.t5070 VPWR 179.399
R2266 VPWR.t4537 VPWR 179.399
R2267 VPWR.t1609 VPWR 179.399
R2268 VPWR.t502 VPWR 179.399
R2269 VPWR.t5404 VPWR 179.399
R2270 VPWR VPWR.t717 179.399
R2271 VPWR VPWR.t4984 179.399
R2272 VPWR.t5380 VPWR 179.399
R2273 VPWR.t3271 VPWR 179.399
R2274 VPWR.t5331 VPWR 179.399
R2275 VPWR VPWR.t5264 179.399
R2276 VPWR VPWR.t5833 179.399
R2277 VPWR VPWR.t1972 179.399
R2278 VPWR VPWR.t5191 179.399
R2279 VPWR.t4236 VPWR.t5586 179.399
R2280 VPWR VPWR.t0 179.399
R2281 VPWR VPWR.t553 179.399
R2282 VPWR VPWR.n1087 179.399
R2283 VPWR VPWR.t1535 179.399
R2284 VPWR VPWR.t62 179.399
R2285 VPWR VPWR.t5291 179.399
R2286 VPWR VPWR.t2752 179.399
R2287 VPWR VPWR.n1088 179.399
R2288 VPWR VPWR.t5110 179.399
R2289 VPWR VPWR.t2497 179.399
R2290 VPWR VPWR.t3675 179.399
R2291 VPWR VPWR.t514 179.399
R2292 VPWR VPWR.t1672 179.399
R2293 VPWR VPWR.t4064 179.399
R2294 VPWR VPWR.t6077 179.399
R2295 VPWR VPWR.t3056 179.399
R2296 VPWR VPWR.t4621 179.399
R2297 VPWR VPWR.t2766 179.399
R2298 VPWR VPWR.t1192 179.399
R2299 VPWR VPWR.t4926 179.399
R2300 VPWR VPWR.t6327 179.399
R2301 VPWR VPWR.t2851 179.399
R2302 VPWR.t2019 VPWR 179.399
R2303 VPWR.t4427 VPWR 179.399
R2304 VPWR.t786 VPWR 179.399
R2305 VPWR.n187 VPWR 179.399
R2306 VPWR.t3542 VPWR 179.399
R2307 VPWR VPWR.t2894 179.399
R2308 VPWR.t977 VPWR 179.399
R2309 VPWR VPWR.t2515 179.399
R2310 VPWR VPWR.n2866 179.399
R2311 VPWR VPWR.t4045 179.399
R2312 VPWR VPWR.t1081 179.399
R2313 VPWR.t3184 VPWR 179.399
R2314 VPWR.t2218 VPWR 179.399
R2315 VPWR.t6179 VPWR 179.399
R2316 VPWR.t1781 VPWR 179.399
R2317 VPWR.t3231 VPWR 179.399
R2318 VPWR.t496 VPWR 179.399
R2319 VPWR.t3928 VPWR 179.399
R2320 VPWR VPWR.t4395 179.399
R2321 VPWR VPWR.t3617 179.399
R2322 VPWR VPWR.t3037 179.399
R2323 VPWR.t5851 VPWR 179.399
R2324 VPWR.t4653 VPWR 179.399
R2325 VPWR VPWR.t3544 179.399
R2326 VPWR VPWR.t1465 179.399
R2327 VPWR VPWR.t2841 179.399
R2328 VPWR VPWR.t1561 179.399
R2329 VPWR VPWR.t3902 179.399
R2330 VPWR VPWR.t6201 179.399
R2331 VPWR VPWR.t2340 179.399
R2332 VPWR VPWR.t3523 179.399
R2333 VPWR VPWR.t5306 179.399
R2334 VPWR VPWR.t3642 179.399
R2335 VPWR VPWR.t2495 179.399
R2336 VPWR VPWR.t3049 179.399
R2337 VPWR VPWR.t6055 179.399
R2338 VPWR VPWR.t2095 179.399
R2339 VPWR.t3712 VPWR 179.399
R2340 VPWR VPWR.t6444 179.399
R2341 VPWR VPWR.t547 179.399
R2342 VPWR VPWR.t346 179.399
R2343 VPWR VPWR.t5077 179.399
R2344 VPWR VPWR.t3799 179.399
R2345 VPWR VPWR.t3393 179.399
R2346 VPWR VPWR.t930 179.399
R2347 VPWR VPWR.t6456 179.399
R2348 VPWR VPWR.t4016 179.399
R2349 VPWR VPWR.t3391 179.399
R2350 VPWR VPWR.t983 179.399
R2351 VPWR.t4056 VPWR 179.399
R2352 VPWR.t4768 VPWR 179.399
R2353 VPWR.n193 VPWR 179.399
R2354 VPWR.t3762 VPWR 179.399
R2355 VPWR.t5311 VPWR 179.399
R2356 VPWR VPWR.t7131 179.399
R2357 VPWR VPWR.t4573 179.399
R2358 VPWR VPWR.t5427 179.399
R2359 VPWR VPWR.t2312 179.399
R2360 VPWR VPWR.t326 179.399
R2361 VPWR VPWR.t1350 179.399
R2362 VPWR VPWR.t4069 179.399
R2363 VPWR VPWR.t5899 179.399
R2364 VPWR VPWR.t3144 179.399
R2365 VPWR VPWR.t409 179.399
R2366 VPWR VPWR.t5941 179.399
R2367 VPWR VPWR.t940 179.399
R2368 VPWR VPWR.t2810 179.399
R2369 VPWR.t5849 VPWR 179.399
R2370 VPWR VPWR.t6155 179.399
R2371 VPWR VPWR.t5406 179.399
R2372 VPWR VPWR.t4704 179.399
R2373 VPWR VPWR.t387 179.399
R2374 VPWR VPWR.t2475 179.399
R2375 VPWR VPWR.t66 179.399
R2376 VPWR VPWR.t520 179.399
R2377 VPWR VPWR.t423 179.399
R2378 VPWR VPWR.t2632 179.399
R2379 VPWR VPWR.t3767 179.399
R2380 VPWR VPWR.t5104 179.399
R2381 VPWR VPWR.t1543 179.399
R2382 VPWR.t3780 VPWR 179.399
R2383 VPWR.t1178 VPWR 179.399
R2384 VPWR VPWR.t3122 179.399
R2385 VPWR VPWR.t5435 179.399
R2386 VPWR VPWR.t3963 179.399
R2387 VPWR VPWR.t2375 179.399
R2388 VPWR VPWR.t1657 179.399
R2389 VPWR.t6035 VPWR 179.399
R2390 VPWR VPWR.t1747 179.399
R2391 VPWR.t5444 VPWR 179.399
R2392 VPWR.t5402 VPWR 179.399
R2393 VPWR.t5326 VPWR 179.399
R2394 VPWR VPWR.n511 179.399
R2395 VPWR VPWR.t5087 179.399
R2396 VPWR VPWR.n2953 179.399
R2397 VPWR VPWR.t2344 179.399
R2398 VPWR.n180 VPWR 179.399
R2399 VPWR.t1831 VPWR 179.399
R2400 VPWR.t5876 VPWR 179.399
R2401 VPWR.t6168 VPWR 179.399
R2402 VPWR VPWR.t2001 179.399
R2403 VPWR VPWR.n2951 179.399
R2404 VPWR.n395 VPWR 179.399
R2405 VPWR VPWR.t4661 179.399
R2406 VPWR.t1181 VPWR 179.399
R2407 VPWR VPWR.t3801 179.399
R2408 VPWR VPWR.t4578 179.399
R2409 VPWR VPWR.t3446 179.399
R2410 VPWR VPWR.t2321 179.399
R2411 VPWR VPWR.t5315 179.399
R2412 VPWR VPWR.t1964 179.399
R2413 VPWR.t6111 VPWR 179.399
R2414 VPWR.t3342 VPWR 179.399
R2415 VPWR VPWR.t3076 179.399
R2416 VPWR.t1432 VPWR 179.399
R2417 VPWR.t1175 VPWR 179.399
R2418 VPWR.t862 VPWR 179.399
R2419 VPWR.t6147 VPWR 179.399
R2420 VPWR VPWR.t2115 179.399
R2421 VPWR VPWR.t1753 179.399
R2422 VPWR VPWR.t5761 179.399
R2423 VPWR VPWR.t1282 179.399
R2424 VPWR VPWR.t854 179.399
R2425 VPWR VPWR.t3083 179.399
R2426 VPWR.t914 VPWR 179.399
R2427 VPWR.t531 VPWR 179.399
R2428 VPWR.t2685 VPWR 179.399
R2429 VPWR.t2945 VPWR 179.399
R2430 VPWR VPWR.t4415 179.399
R2431 VPWR VPWR.t3127 179.399
R2432 VPWR VPWR.t3242 179.399
R2433 VPWR VPWR.t2068 179.399
R2434 VPWR VPWR.t5308 179.399
R2435 VPWR VPWR.t3024 179.399
R2436 VPWR VPWR.t2103 179.399
R2437 VPWR VPWR.t627 179.399
R2438 VPWR.t6079 VPWR 179.399
R2439 VPWR VPWR.t574 179.399
R2440 VPWR.t1173 VPWR 179.399
R2441 VPWR.t3258 VPWR 179.399
R2442 VPWR VPWR.t5972 179.399
R2443 VPWR VPWR.t1804 179.399
R2444 VPWR VPWR.t2972 179.399
R2445 VPWR VPWR.t5363 179.399
R2446 VPWR VPWR.t1145 179.399
R2447 VPWR.t5726 VPWR 179.399
R2448 VPWR.t549 VPWR 179.399
R2449 VPWR VPWR.t1819 179.399
R2450 VPWR VPWR.t662 179.399
R2451 VPWR VPWR.t2310 179.399
R2452 VPWR VPWR.t1507 179.399
R2453 VPWR.t2091 VPWR.t3477 178.242
R2454 VPWR.t6911 VPWR.t1787 178.242
R2455 VPWR.t6828 VPWR.t4576 178.242
R2456 VPWR.t2505 VPWR.t233 178.242
R2457 VPWR VPWR.t6508 177.593
R2458 VPWR.t6065 VPWR.t5020 177.083
R2459 VPWR.t4686 VPWR.t6797 176.4
R2460 VPWR.t4701 VPWR.t6810 176.4
R2461 VPWR.t7031 VPWR.t464 176.4
R2462 VPWR.t5738 VPWR.n729 175.927
R2463 VPWR.t14 VPWR.t4125 175.927
R2464 VPWR.t6258 VPWR.t7111 175.927
R2465 VPWR.t6860 VPWR.t3590 175.927
R2466 VPWR.t5796 VPWR.t3348 175.927
R2467 VPWR.t1031 VPWR.t1927 175.493
R2468 VPWR VPWR.t522 174.769
R2469 VPWR VPWR.t3960 174.769
R2470 VPWR.t1619 VPWR.t175 173.612
R2471 VPWR.t2618 VPWR.t5914 173.612
R2472 VPWR.t6574 VPWR 172.826
R2473 VPWR.t3985 VPWR 172.454
R2474 VPWR.t5422 VPWR 172.454
R2475 VPWR.t5160 VPWR.t1167 172.454
R2476 VPWR.t6404 VPWR.t979 171.633
R2477 VPWR.t1356 VPWR.t137 171.297
R2478 VPWR.t157 VPWR.t2380 171.297
R2479 VPWR.t1111 VPWR.t5660 171.297
R2480 VPWR.t879 VPWR.t6946 171.297
R2481 VPWR.t1478 VPWR.t7040 171.297
R2482 VPWR.t6688 VPWR.t1692 171.297
R2483 VPWR.t1676 VPWR.t104 171.297
R2484 VPWR.t1056 VPWR.t6501 171.297
R2485 VPWR.t7004 VPWR.t5985 171.297
R2486 VPWR.t3880 VPWR.t7020 171.297
R2487 VPWR.t4435 VPWR.t7013 171.297
R2488 VPWR.t5790 VPWR.t6371 171.297
R2489 VPWR.t2650 VPWR.t177 171.297
R2490 VPWR.t142 VPWR.t2957 171.297
R2491 VPWR.t220 VPWR.t5460 171.297
R2492 VPWR.t7029 VPWR.t5089 171.297
R2493 VPWR.t6474 VPWR.t5707 171.297
R2494 VPWR.t6776 VPWR.t932 171.297
R2495 VPWR.t6386 VPWR.t2323 171.297
R2496 VPWR.t39 VPWR.t435 171.297
R2497 VPWR.t460 VPWR.t6399 171.297
R2498 VPWR.t6564 VPWR.t191 171.297
R2499 VPWR.t125 VPWR.t283 171.297
R2500 VPWR.t1913 VPWR.t6375 171.297
R2501 VPWR.t153 VPWR.t3899 171.297
R2502 VPWR.t2932 VPWR.t28 171.297
R2503 VPWR.t6616 VPWR.t186 171.297
R2504 VPWR.t120 VPWR.t1463 171.297
R2505 VPWR.t6460 VPWR.t4171 171.297
R2506 VPWR.t2694 VPWR.t6462 171.297
R2507 VPWR.t7046 VPWR.t5095 171.297
R2508 VPWR.t584 VPWR.t7044 171.297
R2509 VPWR.t6942 VPWR.t1833 171.297
R2510 VPWR.t6655 VPWR.t1330 171.297
R2511 VPWR.t2058 VPWR.t101 171.297
R2512 VPWR.t6157 VPWR.t6598 171.297
R2513 VPWR.t216 VPWR.t1751 171.297
R2514 VPWR.t4565 VPWR.t302 171.297
R2515 VPWR.t3915 VPWR 170.139
R2516 VPWR.t6377 VPWR 170.139
R2517 VPWR.t4680 VPWR.t3830 169.25
R2518 VPWR.t6675 VPWR.t5218 168.982
R2519 VPWR.t2483 VPWR.t6873 168.982
R2520 VPWR.t2257 VPWR.t906 168.982
R2521 VPWR.t4804 VPWR.t3054 168.982
R2522 VPWR VPWR.t1886 167.825
R2523 VPWR.t4694 VPWR.t277 166.865
R2524 VPWR.t31 VPWR.t235 166.865
R2525 VPWR.t4697 VPWR.t289 166.865
R2526 VPWR.t7066 VPWR.t5584 166.667
R2527 VPWR.t6996 VPWR.t6783 166.667
R2528 VPWR.t795 VPWR.t2033 166.667
R2529 VPWR.t2394 VPWR.t7022 166.667
R2530 VPWR.t2125 VPWR.t7010 166.667
R2531 VPWR.t1929 VPWR.n946 165.51
R2532 VPWR.t668 VPWR.n928 165.51
R2533 VPWR.t2638 VPWR.n3358 165.51
R2534 VPWR.t2519 VPWR 165.51
R2535 VPWR.t3101 VPWR.t6626 165.51
R2536 VPWR.t6995 VPWR.t6576 165.51
R2537 VPWR.n749 VPWR.t6297 165.51
R2538 VPWR.t6006 VPWR.n755 165.51
R2539 VPWR.t3265 VPWR.n760 165.51
R2540 VPWR.t4422 VPWR.n156 165.51
R2541 VPWR.t6317 VPWR.n142 165.51
R2542 VPWR.n1782 VPWR.t1665 165.51
R2543 VPWR.n1092 VPWR.t3983 165.51
R2544 VPWR.t5423 VPWR.n1938 165.51
R2545 VPWR.t1847 VPWR.n2879 165.51
R2546 VPWR.t1328 VPWR.n2880 165.51
R2547 VPWR.n2748 VPWR.t5012 165.51
R2548 VPWR.n517 VPWR.t3942 165.51
R2549 VPWR.t2598 VPWR.n394 165.51
R2550 VPWR.n377 VPWR.t437 165.51
R2551 VPWR.t5260 VPWR.t6496 164.352
R2552 VPWR.n1386 VPWR.t5270 164.352
R2553 VPWR.t6498 VPWR.t5496 164.352
R2554 VPWR.t3677 VPWR.t4610 164.352
R2555 VPWR.t5803 VPWR.t3679 164.352
R2556 VPWR.t6651 VPWR.t3970 164.352
R2557 VPWR.t1280 VPWR.t6619 164.352
R2558 VPWR.t6756 VPWR.t5511 164.352
R2559 VPWR.t4466 VPWR.t5183 164.352
R2560 VPWR.n523 VPWR.t184 164.352
R2561 VPWR.t6657 VPWR.t1976 164.352
R2562 VPWR.t2453 VPWR.t6762 164.352
R2563 VPWR.t6862 VPWR 163.195
R2564 VPWR.t4682 VPWR.t3349 163.195
R2565 VPWR.t6977 VPWR.t110 162.037
R2566 VPWR.t6777 VPWR.t7002 162.037
R2567 VPWR.t123 VPWR.t6542 162.037
R2568 VPWR.t56 VPWR.t2694 162.037
R2569 VPWR.t5095 VPWR.t6015 162.037
R2570 VPWR.t6591 VPWR.t2392 162.037
R2571 VPWR.t198 VPWR.t1918 162.037
R2572 VPWR.t6335 VPWR.t7054 160.881
R2573 VPWR.t1216 VPWR.t5718 159.722
R2574 VPWR.t1743 VPWR.t2569 159.722
R2575 VPWR.t4872 VPWR.t7016 159.722
R2576 VPWR.t2150 VPWR.t5809 159.722
R2577 VPWR.t5720 VPWR.t3710 159.722
R2578 VPWR.t6303 VPWR.t5705 159.722
R2579 VPWR.t3890 VPWR.t6063 159.722
R2580 VPWR.t2225 VPWR.t6059 159.722
R2581 VPWR.t2593 VPWR.t6243 159.722
R2582 VPWR.t3307 VPWR.t287 159.722
R2583 VPWR.t1387 VPWR.t5883 159.722
R2584 VPWR.t6252 VPWR.t2369 159.722
R2585 VPWR.t2894 VPWR.t363 159.722
R2586 VPWR.t1503 VPWR.t5248 159.722
R2587 VPWR.t2206 VPWR.t3172 159.722
R2588 VPWR.t2202 VPWR.t1403 159.722
R2589 VPWR.t1603 VPWR.t4529 159.722
R2590 VPWR.t1118 VPWR.t5989 159.722
R2591 VPWR.t1513 VPWR.t2365 159.722
R2592 VPWR.t5072 VPWR.t3154 159.722
R2593 VPWR.t6270 VPWR.t5208 158.565
R2594 VPWR.t5085 VPWR 158.565
R2595 VPWR.t5587 VPWR.t297 158.565
R2596 VPWR VPWR.t6876 157.407
R2597 VPWR.t1130 VPWR 157.407
R2598 VPWR.t6789 VPWR.t671 157.407
R2599 VPWR.n1276 VPWR.t4379 157.407
R2600 VPWR.t3434 VPWR.t1067 157.407
R2601 VPWR.t2066 VPWR.t6381 157.407
R2602 VPWR VPWR.t4794 157.407
R2603 VPWR VPWR.t6883 157.407
R2604 VPWR.t1763 VPWR.t5713 157.407
R2605 VPWR.t1581 VPWR.t764 157.407
R2606 VPWR.t2766 VPWR.t5887 157.407
R2607 VPWR.t3795 VPWR.t5319 157.407
R2608 VPWR.t6155 VPWR.t2914 157.407
R2609 VPWR.t2240 VPWR.t2577 157.407
R2610 VPWR.t4998 VPWR 157.407
R2611 VPWR.t4496 VPWR.t5326 157.407
R2612 VPWR.t3446 VPWR.t310 157.407
R2613 VPWR.t4890 VPWR.t1769 157.407
R2614 VPWR.t1964 VPWR.t1486 157.407
R2615 VPWR.n374 VPWR.t5490 157.407
R2616 VPWR.t5122 VPWR.t6270 156.25
R2617 VPWR VPWR.t3411 156.25
R2618 VPWR.t5911 VPWR 156.25
R2619 VPWR.t5868 VPWR.t973 156.25
R2620 VPWR.t297 VPWR.t2805 156.25
R2621 VPWR VPWR.t1467 156.25
R2622 VPWR.t2898 VPWR 156.25
R2623 VPWR.t3401 VPWR 156.25
R2624 VPWR.t5018 VPWR.t6189 155.094
R2625 VPWR.t5022 VPWR.t2170 155.094
R2626 VPWR.t6048 VPWR.t5395 155.094
R2627 VPWR.t403 VPWR.t3192 155.094
R2628 VPWR.t405 VPWR.t5237 155.094
R2629 VPWR VPWR.t6629 153.935
R2630 VPWR.t1083 VPWR 153.935
R2631 VPWR.t5569 VPWR 153.935
R2632 VPWR.t6178 VPWR.t7094 152.779
R2633 VPWR.t4598 VPWR.t6280 152.779
R2634 VPWR.t4600 VPWR.t6274 152.779
R2635 VPWR.t6692 VPWR.t4183 152.779
R2636 VPWR.t6690 VPWR.t4181 152.779
R2637 VPWR.t6780 VPWR.t2046 152.779
R2638 VPWR.t6381 VPWR.t6857 152.779
R2639 VPWR.t4695 VPWR 152.779
R2640 VPWR.t5020 VPWR 151.62
R2641 VPWR.t6788 VPWR 151.62
R2642 VPWR.n1385 VPWR.t6876 151.62
R2643 VPWR.t7060 VPWR 151.62
R2644 VPWR.t407 VPWR 151.62
R2645 VPWR.t3228 VPWR 151.62
R2646 VPWR.t4004 VPWR 151.62
R2647 VPWR.t4431 VPWR 151.62
R2648 VPWR.t178 VPWR.t2959 151.62
R2649 VPWR.t4105 VPWR.t141 151.62
R2650 VPWR VPWR.t143 151.62
R2651 VPWR.t1320 VPWR 151.62
R2652 VPWR.t269 VPWR 151.62
R2653 VPWR VPWR.t6830 151.62
R2654 VPWR.t939 VPWR 151.62
R2655 VPWR.t2979 VPWR.t6125 150.464
R2656 VPWR.t950 VPWR.t2174 150.464
R2657 VPWR.t3821 VPWR.t1595 150.464
R2658 VPWR.t4717 VPWR.t3716 150.464
R2659 VPWR.t3219 VPWR.t6365 150.011
R2660 VPWR VPWR.t6647 148.988
R2661 VPWR.t3949 VPWR.t4220 148.149
R2662 VPWR.t118 VPWR.t4692 148.149
R2663 VPWR.t3992 VPWR.t3471 148.149
R2664 VPWR.t6566 VPWR.t3840 148.149
R2665 VPWR.t6560 VPWR.t6617 148.149
R2666 VPWR.t6562 VPWR.t5961 148.149
R2667 VPWR.t134 VPWR.t1266 148.149
R2668 VPWR.t183 VPWR.t129 148.149
R2669 VPWR.t4228 VPWR.t803 146.992
R2670 VPWR.n2863 VPWR.t4173 146.992
R2671 VPWR.t586 VPWR.n2865 146.992
R2672 VPWR VPWR.t160 145.833
R2673 VPWR.n923 VPWR.t4962 145.833
R2674 VPWR VPWR.t6387 145.833
R2675 VPWR.t281 VPWR.t2918 145.833
R2676 VPWR.t3303 VPWR.n604 145.833
R2677 VPWR.t2541 VPWR.t6927 145.833
R2678 VPWR.t1788 VPWR.t6923 145.833
R2679 VPWR VPWR.t121 145.833
R2680 VPWR.t6490 VPWR 144.677
R2681 VPWR VPWR.t6480 144.677
R2682 VPWR.t6496 VPWR 144.677
R2683 VPWR VPWR.t6482 144.677
R2684 VPWR VPWR.t6486 144.677
R2685 VPWR.t43 VPWR 144.677
R2686 VPWR.t6879 VPWR 144.677
R2687 VPWR.t970 VPWR.t5122 144.677
R2688 VPWR.t1909 VPWR 144.677
R2689 VPWR.t5815 VPWR 144.677
R2690 VPWR.t6331 VPWR 144.677
R2691 VPWR VPWR.t6498 144.677
R2692 VPWR VPWR.t6861 144.677
R2693 VPWR VPWR.t3677 144.677
R2694 VPWR VPWR.t1958 144.677
R2695 VPWR.t908 VPWR 144.677
R2696 VPWR.t643 VPWR 144.677
R2697 VPWR VPWR.t6466 144.677
R2698 VPWR VPWR.t6472 144.677
R2699 VPWR VPWR.t118 144.677
R2700 VPWR.t477 VPWR 144.677
R2701 VPWR.t6991 VPWR 144.677
R2702 VPWR VPWR.t6488 144.677
R2703 VPWR.t475 VPWR 144.677
R2704 VPWR.t5880 VPWR 144.677
R2705 VPWR.t2166 VPWR 144.677
R2706 VPWR VPWR.t3961 144.677
R2707 VPWR VPWR.t6659 144.677
R2708 VPWR VPWR.t1288 144.677
R2709 VPWR VPWR.t19 144.677
R2710 VPWR VPWR.t2648 144.677
R2711 VPWR VPWR.t1761 144.677
R2712 VPWR.t936 VPWR 144.677
R2713 VPWR VPWR.t6756 144.677
R2714 VPWR VPWR.t4466 144.677
R2715 VPWR.t6649 VPWR 144.677
R2716 VPWR VPWR.t6661 144.677
R2717 VPWR VPWR.t5043 144.677
R2718 VPWR VPWR.t6655 144.677
R2719 VPWR VPWR.t6645 144.677
R2720 VPWR.t6643 VPWR 144.677
R2721 VPWR.t6665 VPWR 144.677
R2722 VPWR VPWR.t4986 144.677
R2723 VPWR VPWR.t6892 144.677
R2724 VPWR VPWR.t6585 144.677
R2725 VPWR VPWR.t2331 144.677
R2726 VPWR.t3930 VPWR.t2004 144.677
R2727 VPWR VPWR.t6620 144.677
R2728 VPWR VPWR.t6657 144.677
R2729 VPWR.t5567 VPWR 144.677
R2730 VPWR VPWR.t4684 144.677
R2731 VPWR.t6762 VPWR 144.677
R2732 VPWR.t6366 VPWR 143.519
R2733 VPWR.t5479 VPWR.t837 143.519
R2734 VPWR.t837 VPWR.t4448 143.519
R2735 VPWR.t4448 VPWR.t2161 143.519
R2736 VPWR.t6577 VPWR.t5140 143.519
R2737 VPWR.t5355 VPWR.t3142 143.519
R2738 VPWR.t4219 VPWR.t7039 143.519
R2739 VPWR.t6504 VPWR.t3825 143.519
R2740 VPWR.t6340 VPWR 143.519
R2741 VPWR.t156 VPWR 143.519
R2742 VPWR.t3081 VPWR.t1921 143.519
R2743 VPWR.t3007 VPWR.t6500 143.028
R2744 VPWR.t3005 VPWR.t16 143.028
R2745 VPWR.t4681 VPWR.t241 143.028
R2746 VPWR.t33 VPWR.t293 143.028
R2747 VPWR.t4689 VPWR.t291 143.028
R2748 VPWR.t5208 VPWR.t897 142.362
R2749 VPWR.t2361 VPWR 141.837
R2750 VPWR.t1109 VPWR.t5662 141.204
R2751 VPWR.t4255 VPWR.t879 141.204
R2752 VPWR.t6320 VPWR.t1676 141.204
R2753 VPWR.t5009 VPWR.n833 141.204
R2754 VPWR.t5507 VPWR.t5790 141.204
R2755 VPWR.t435 VPWR.t4747 141.204
R2756 VPWR.t6220 VPWR.t460 141.204
R2757 VPWR.t2134 VPWR.t2342 141.204
R2758 VPWR.t6248 VPWR.t6157 141.204
R2759 VPWR VPWR.n934 138.889
R2760 VPWR.t6365 VPWR.t5051 138.889
R2761 VPWR.t4 VPWR.t314 138.889
R2762 VPWR VPWR.n827 138.889
R2763 VPWR VPWR.n3261 138.889
R2764 VPWR.t6542 VPWR.t1794 138.889
R2765 VPWR.t4879 VPWR.n953 137.732
R2766 VPWR VPWR.t3789 137.732
R2767 VPWR.t6636 VPWR 137.732
R2768 VPWR.t1128 VPWR.t7014 137.732
R2769 VPWR VPWR.t6042 137.732
R2770 VPWR VPWR.t3635 137.732
R2771 VPWR.t4042 VPWR 137.732
R2772 VPWR VPWR.t1490 137.732
R2773 VPWR.t2878 VPWR 137.732
R2774 VPWR VPWR.t5626 137.732
R2775 VPWR VPWR.t1103 137.732
R2776 VPWR VPWR.t1873 137.732
R2777 VPWR VPWR.t4429 137.732
R2778 VPWR VPWR.t5740 137.732
R2779 VPWR.t3841 VPWR 137.732
R2780 VPWR.t7109 VPWR.t4558 137.732
R2781 VPWR.t6970 VPWR.t6968 137.732
R2782 VPWR.t981 VPWR 137.732
R2783 VPWR VPWR.t6396 137.732
R2784 VPWR VPWR.t4280 137.732
R2785 VPWR.t1867 VPWR 137.732
R2786 VPWR VPWR.t1318 137.732
R2787 VPWR.t972 VPWR 137.732
R2788 VPWR VPWR.t3772 137.732
R2789 VPWR VPWR.t253 137.732
R2790 VPWR.t535 VPWR 137.732
R2791 VPWR VPWR.t541 137.732
R2792 VPWR.t5527 VPWR 137.732
R2793 VPWR.t3349 VPWR 137.732
R2794 VPWR.t729 VPWR 137.732
R2795 VPWR.t6706 VPWR.t3200 137.732
R2796 VPWR.t733 VPWR 137.732
R2797 VPWR VPWR.t5339 137.732
R2798 VPWR VPWR.t1749 137.732
R2799 VPWR.t5112 VPWR 137.732
R2800 VPWR VPWR.t2859 137.732
R2801 VPWR VPWR.t2608 136.575
R2802 VPWR VPWR.t211 136.575
R2803 VPWR VPWR.t4365 136.575
R2804 VPWR.t4226 VPWR.t5998 136.575
R2805 VPWR.t6726 VPWR.t6724 136.575
R2806 VPWR.t3683 VPWR.t3264 136.575
R2807 VPWR.t2357 VPWR.n128 136.575
R2808 VPWR.t1635 VPWR.t6319 136.575
R2809 VPWR VPWR.t2455 136.575
R2810 VPWR.t5438 VPWR.t4992 136.575
R2811 VPWR VPWR.t1946 135.417
R2812 VPWR.t6733 VPWR 135.417
R2813 VPWR VPWR.t1339 135.417
R2814 VPWR VPWR.t5835 135.417
R2815 VPWR.t3371 VPWR.t178 135.417
R2816 VPWR.t141 VPWR.t4109 135.417
R2817 VPWR.t4794 VPWR.t239 135.417
R2818 VPWR.t5001 VPWR 135.417
R2819 VPWR.t6486 VPWR.t7136 134.26
R2820 VPWR.t5485 VPWR.t6535 134.26
R2821 VPWR.t4134 VPWR.t5003 134.26
R2822 VPWR.t845 VPWR.n266 134.26
R2823 VPWR.t2335 VPWR 133.102
R2824 VPWR.t4316 VPWR.t2437 133.102
R2825 VPWR.t1054 VPWR.t2158 133.102
R2826 VPWR.t6615 VPWR 133.102
R2827 VPWR.t334 VPWR 133.102
R2828 VPWR.t3283 VPWR 133.102
R2829 VPWR.t201 VPWR.t6288 133.102
R2830 VPWR VPWR.t2727 133.102
R2831 VPWR.t90 VPWR 133.102
R2832 VPWR.t49 VPWR 133.102
R2833 VPWR.t277 VPWR.t29 132.608
R2834 VPWR.t3910 VPWR.t5868 130.787
R2835 VPWR.t6609 VPWR 130.787
R2836 VPWR.t5157 VPWR.t6715 130.787
R2837 VPWR.t1838 VPWR.t3978 129.631
R2838 VPWR.t4904 VPWR.t1997 129.631
R2839 VPWR.t4385 VPWR.t429 129.631
R2840 VPWR.t4627 VPWR.t3286 129.631
R2841 VPWR.t4492 VPWR.t1835 129.631
R2842 VPWR.t4113 VPWR.t1135 129.631
R2843 VPWR.t2665 VPWR.t3650 129.631
R2844 VPWR.t1745 VPWR.t2849 129.631
R2845 VPWR.t2616 VPWR.t5369 129.631
R2846 VPWR.t3464 VPWR.t5289 129.631
R2847 VPWR.t1783 VPWR.t6067 129.631
R2848 VPWR.t3260 VPWR.t4785 129.631
R2849 VPWR.t2405 VPWR.t4115 129.631
R2850 VPWR.t6075 VPWR.t5313 129.631
R2851 VPWR.t5533 VPWR.t3720 129.631
R2852 VPWR.t5550 VPWR.t2168 129.631
R2853 VPWR.n101 VPWR.t5416 129.631
R2854 VPWR.t4258 VPWR.n100 129.631
R2855 VPWR.n99 VPWR.t707 129.631
R2856 VPWR.t2799 VPWR.n98 129.631
R2857 VPWR.n97 VPWR.t6442 129.631
R2858 VPWR.n3435 VPWR.t754 129.631
R2859 VPWR.n955 VPWR.t6446 129.631
R2860 VPWR.t3014 VPWR.t4494 129.631
R2861 VPWR.t147 VPWR.t3531 129.631
R2862 VPWR.t5716 VPWR.t1216 129.631
R2863 VPWR.t2571 VPWR.t1743 129.631
R2864 VPWR.t7016 VPWR.t4868 129.631
R2865 VPWR.t5809 VPWR.t2152 129.631
R2866 VPWR.t6280 VPWR.t4602 129.631
R2867 VPWR.t6276 VPWR.t4598 129.631
R2868 VPWR.t6274 VPWR.t4604 129.631
R2869 VPWR.t6686 VPWR.t4185 129.631
R2870 VPWR.t4183 VPWR.t6686 129.631
R2871 VPWR.t6684 VPWR.t4187 129.631
R2872 VPWR.t4181 VPWR.t6684 129.631
R2873 VPWR.t2046 VPWR.t6789 129.631
R2874 VPWR.t6855 VPWR.t6669 129.631
R2875 VPWR.t3708 VPWR.t5720 129.631
R2876 VPWR.t7011 VPWR 129.631
R2877 VPWR.t3315 VPWR.t5658 129.631
R2878 VPWR.t5056 VPWR.t2901 129.631
R2879 VPWR.t6877 VPWR 129.631
R2880 VPWR.t114 VPWR 129.631
R2881 VPWR.t705 VPWR.t2427 129.631
R2882 VPWR.t6063 VPWR.t3888 129.631
R2883 VPWR.t6057 VPWR.t2225 129.631
R2884 VPWR.t4192 VPWR.t1234 129.631
R2885 VPWR.t1875 VPWR.t5028 129.631
R2886 VPWR.t4567 VPWR.t5515 129.631
R2887 VPWR.t175 VPWR.t187 129.631
R2888 VPWR.t6812 VPWR 129.631
R2889 VPWR VPWR.t6812 129.631
R2890 VPWR.t4209 VPWR.t167 129.631
R2891 VPWR.t4052 VPWR.t4714 129.631
R2892 VPWR.t2245 VPWR.t2415 129.631
R2893 VPWR.t2614 VPWR.t5498 129.631
R2894 VPWR.t3945 VPWR.t5433 129.631
R2895 VPWR.t1593 VPWR.t1413 129.631
R2896 VPWR.t6458 VPWR.t5775 129.631
R2897 VPWR.t2431 VPWR.t600 129.631
R2898 VPWR.t5531 VPWR.t5281 129.631
R2899 VPWR.t4592 VPWR.t4127 129.631
R2900 VPWR.t664 VPWR.t6210 129.631
R2901 VPWR.t6245 VPWR.t2593 129.631
R2902 VPWR.n724 VPWR.t5404 129.631
R2903 VPWR.t717 VPWR.t1950 129.631
R2904 VPWR.t703 VPWR.t2479 129.631
R2905 VPWR.t2947 VPWR.t5861 129.631
R2906 VPWR.t4954 VPWR.t993 129.631
R2907 VPWR.t4984 VPWR.t4935 129.631
R2908 VPWR.t4888 VPWR.t4441 129.631
R2909 VPWR.t1553 VPWR.t1712 129.631
R2910 VPWR.t570 VPWR.t6268 129.631
R2911 VPWR.t1159 VPWR.t823 129.631
R2912 VPWR.t4097 VPWR.t1385 129.631
R2913 VPWR.t2678 VPWR.t5380 129.631
R2914 VPWR.t5574 VPWR.t448 129.631
R2915 VPWR.t6241 VPWR.t5299 129.631
R2916 VPWR.t6349 VPWR.t3644 129.631
R2917 VPWR.t4391 VPWR.t5636 129.631
R2918 VPWR.t1851 VPWR.t4485 129.631
R2919 VPWR.t2385 VPWR.t330 129.631
R2920 VPWR.t3499 VPWR.t5780 129.631
R2921 VPWR.t4058 VPWR.t5331 129.631
R2922 VPWR.t3996 VPWR.t2531 129.631
R2923 VPWR.t5414 VPWR.t1755 129.631
R2924 VPWR.t1395 VPWR.t721 129.631
R2925 VPWR.t1960 VPWR.t709 129.631
R2926 VPWR.t701 VPWR.t1505 129.631
R2927 VPWR.t3921 VPWR.t1827 129.631
R2928 VPWR.t1605 VPWR.t4943 129.631
R2929 VPWR.t5264 VPWR.t2097 129.631
R2930 VPWR.t1453 VPWR.t1663 129.631
R2931 VPWR.t224 VPWR.t6957 129.631
R2932 VPWR.t129 VPWR.t938 129.631
R2933 VPWR.t760 VPWR.t3495 129.631
R2934 VPWR.n1088 VPWR.t5151 129.631
R2935 VPWR.t3675 VPWR.t5024 129.631
R2936 VPWR.t875 VPWR.t5800 129.631
R2937 VPWR.t514 VPWR.t3387 129.631
R2938 VPWR.t1672 VPWR.t3850 129.631
R2939 VPWR.t1717 VPWR.t1260 129.631
R2940 VPWR.t2535 VPWR.t1674 129.631
R2941 VPWR.t1985 VPWR.t631 129.631
R2942 VPWR.t4064 VPWR.t2089 129.631
R2943 VPWR.t5965 VPWR.n1936 129.631
R2944 VPWR.t5883 VPWR.t1389 129.631
R2945 VPWR.t2367 VPWR.t6252 129.631
R2946 VPWR.n1937 VPWR.t5844 129.631
R2947 VPWR.t2070 VPWR.t5420 129.631
R2948 VPWR.t2851 VPWR.t4645 129.631
R2949 VPWR.t3624 VPWR.t4427 129.631
R2950 VPWR.t5558 VPWR.t2853 129.631
R2951 VPWR.t4739 VPWR.t4956 129.631
R2952 VPWR.n2861 VPWR.t1310 129.631
R2953 VPWR.t1846 VPWR.t2035 129.631
R2954 VPWR.t4195 VPWR.t1879 129.631
R2955 VPWR.t2142 VPWR.t4906 129.631
R2956 VPWR.t604 VPWR.t1447 129.631
R2957 VPWR.t1171 VPWR.t1276 129.631
R2958 VPWR.t1773 VPWR.t4357 129.631
R2959 VPWR.t3515 VPWR.t2756 129.631
R2960 VPWR.t5678 VPWR.t3184 129.631
R2961 VPWR.t723 VPWR.t4310 129.631
R2962 VPWR.t4847 VPWR.t2517 129.631
R2963 VPWR.t4367 VPWR.t2319 129.631
R2964 VPWR.t2429 VPWR.t5699 129.631
R2965 VPWR.t6193 VPWR.t6000 129.631
R2966 VPWR.t756 VPWR.t2009 129.631
R2967 VPWR.t1133 VPWR.t4539 129.631
R2968 VPWR.t4969 VPWR.t2218 129.631
R2969 VPWR.t4018 VPWR.t5821 129.631
R2970 VPWR.t2144 VPWR.t3231 129.631
R2971 VPWR.t2714 VPWR.t5978 129.631
R2972 VPWR.t2269 VPWR.t3225 129.631
R2973 VPWR.t1449 VPWR.t4918 129.631
R2974 VPWR.t1278 VPWR.t458 129.631
R2975 VPWR.t4361 VPWR.t5770 129.631
R2976 VPWR.t3246 VPWR.t4162 129.631
R2977 VPWR.t4031 VPWR.t1844 129.631
R2978 VPWR.t3262 VPWR.t3928 129.631
R2979 VPWR.t1549 VPWR.t494 129.631
R2980 VPWR.t2661 VPWR.t3607 129.631
R2981 VPWR.t6282 VPWR.t5709 129.631
R2982 VPWR.t3546 VPWR.t4238 129.631
R2983 VPWR.t4353 VPWR.t3186 129.631
R2984 VPWR.t681 VPWR.t4545 129.631
R2985 VPWR.t1474 VPWR.t5724 129.631
R2986 VPWR.t4395 VPWR.t6159 129.631
R2987 VPWR.t1645 VPWR.t4189 129.631
R2988 VPWR.t1706 VPWR.t2132 129.631
R2989 VPWR.t1228 VPWR.t1007 129.631
R2990 VPWR.t5036 VPWR.t5840 129.631
R2991 VPWR.t4758 VPWR.t2888 129.631
R2992 VPWR.t2200 VPWR.t1089 129.631
R2993 VPWR.t4766 VPWR.t5851 129.631
R2994 VPWR.t3093 VPWR.t4446 129.631
R2995 VPWR.t3853 VPWR.t3815 129.631
R2996 VPWR.t782 VPWR.t2471 129.631
R2997 VPWR.t3774 VPWR.t2493 129.631
R2998 VPWR.t3364 VPWR.t5452 129.631
R2999 VPWR.t4940 VPWR.t3886 129.631
R3000 VPWR.t944 VPWR.t4814 129.631
R3001 VPWR.t4253 VPWR.t4653 129.631
R3002 VPWR.t5172 VPWR.t1765 129.631
R3003 VPWR.t6150 VPWR.t4297 129.631
R3004 VPWR.t5481 VPWR.t4861 129.631
R3005 VPWR.t2056 VPWR.t4706 129.631
R3006 VPWR.t1421 VPWR.t2212 129.631
R3007 VPWR.t3588 VPWR.t744 129.631
R3008 VPWR.t3213 VPWR.t6109 129.631
R3009 VPWR.t3544 VPWR.t5060 129.631
R3010 VPWR.t4512 VPWR.t4008 129.631
R3011 VPWR.t3596 VPWR.t6088 129.631
R3012 VPWR.t4589 VPWR.t5630 129.631
R3013 VPWR.t4454 VPWR.t4351 129.631
R3014 VPWR.t6208 VPWR.t6218 129.631
R3015 VPWR.t3807 VPWR.t60 129.631
R3016 VPWR.t4024 VPWR.t3725 129.631
R3017 VPWR.t1465 VPWR.t1654 129.631
R3018 VPWR.t4914 VPWR.t3817 129.631
R3019 VPWR.t675 VPWR.t488 129.631
R3020 VPWR.t4874 VPWR.t2626 129.631
R3021 VPWR.t3353 VPWR.t6191 129.631
R3022 VPWR.t6053 VPWR.t4490 129.631
R3023 VPWR.t3168 VPWR.t4614 129.631
R3024 VPWR.t5272 VPWR.t4151 129.631
R3025 VPWR.t2841 VPWR.t1853 129.631
R3026 VPWR.t1670 VPWR.t3031 129.631
R3027 VPWR.t2923 VPWR.t6083 129.631
R3028 VPWR.t5668 VPWR.t1249 129.631
R3029 VPWR.t3379 VPWR.t472 129.631
R3030 VPWR.t829 VPWR.t3451 129.631
R3031 VPWR.t4640 VPWR.t3947 129.631
R3032 VPWR.t3049 VPWR.t2060 129.631
R3033 VPWR.t4856 VPWR.t498 129.631
R3034 VPWR.t492 VPWR.t7140 129.631
R3035 VPWR.t3855 VPWR.t7085 129.631
R3036 VPWR.t1194 VPWR.t391 129.631
R3037 VPWR.t1925 VPWR.t4929 129.631
R3038 VPWR.t2192 VPWR.t5955 129.631
R3039 VPWR.t4543 VPWR.t2229 129.631
R3040 VPWR.t6055 VPWR.t2407 129.631
R3041 VPWR.t2797 VPWR.t1417 129.631
R3042 VPWR.t7123 VPWR.t3176 129.631
R3043 VPWR.t3333 VPWR.t3466 129.631
R3044 VPWR.t4458 VPWR.t4806 129.631
R3045 VPWR.t4636 VPWR.t5359 129.631
R3046 VPWR.t2249 VPWR.t4594 129.631
R3047 VPWR.t2425 VPWR.t3035 129.631
R3048 VPWR.t2095 VPWR.t6085 129.631
R3049 VPWR.t5766 VPWR.t5994 129.631
R3050 VPWR.t1759 VPWR.t3194 129.631
R3051 VPWR.t1678 VPWR.t4920 129.631
R3052 VPWR.t1274 VPWR.t679 129.631
R3053 VPWR.t807 VPWR.t2451 129.631
R3054 VPWR.t4643 VPWR.t5943 129.631
R3055 VPWR.t2017 VPWR.t533 129.631
R3056 VPWR.t3537 VPWR.t3712 129.631
R3057 VPWR.t3782 VPWR.t2473 129.631
R3058 VPWR.t5449 VPWR.t2299 129.631
R3059 VPWR.t5509 VPWR.t5605 129.631
R3060 VPWR.t3673 VPWR.t1183 129.631
R3061 VPWR.t1680 VPWR.t3443 129.631
R3062 VPWR.t72 VPWR.t4504 129.631
R3063 VPWR.t6307 VPWR.t1286 129.631
R3064 VPWR.t6444 VPWR.t1409 129.631
R3065 VPWR.n2324 VPWR.n2318 129.631
R3066 VPWR.t5957 VPWR.t4267 129.631
R3067 VPWR.t4274 VPWR.t1555 129.631
R3068 VPWR.t5759 VPWR.t572 129.631
R3069 VPWR.t2190 VPWR.t2441 129.631
R3070 VPWR.t3714 VPWR.t592 129.631
R3071 VPWR.t2105 VPWR.t2146 129.631
R3072 VPWR.t815 VPWR.t1482 129.631
R3073 VPWR.t4119 VPWR.t4571 129.631
R3074 VPWR.t3799 VPWR.t5301 129.631
R3075 VPWR.t6456 VPWR.t4933 129.631
R3076 VPWR.t6435 VPWR.t2776 129.631
R3077 VPWR.t1815 VPWR.t2074 129.631
R3078 VPWR.t3249 VPWR.t5026 129.631
R3079 VPWR.t4016 VPWR.t660 129.631
R3080 VPWR.t4121 VPWR.t1040 129.631
R3081 VPWR.t1855 VPWR.t1344 129.631
R3082 VPWR.t1888 VPWR.t2411 129.631
R3083 VPWR.t555 VPWR.t2156 129.631
R3084 VPWR.t713 VPWR.t2382 129.631
R3085 VPWR.t5755 VPWR.t869 129.631
R3086 VPWR.t5937 VPWR.t312 129.631
R3087 VPWR.t983 VPWR.t4845 129.631
R3088 VPWR.t369 VPWR.t5293 129.631
R3089 VPWR.t3174 VPWR.t2206 129.631
R3090 VPWR.t1403 VPWR.t2204 129.631
R3091 VPWR.t4529 VPWR.t1601 129.631
R3092 VPWR.t6311 VPWR.n193 129.631
R3093 VPWR.t3389 VPWR.t3762 129.631
R3094 VPWR.t5989 VPWR.t1120 129.631
R3095 VPWR.t7083 VPWR.t2718 129.631
R3096 VPWR.t4663 VPWR.t2172 129.631
R3097 VPWR.t3418 VPWR.t564 129.631
R3098 VPWR.t5903 VPWR.t740 129.631
R3099 VPWR.t2700 VPWR.t6105 129.631
R3100 VPWR.t1884 VPWR.t6017 129.631
R3101 VPWR.t5503 VPWR.t1501 129.631
R3102 VPWR.t4573 VPWR.t6324 129.631
R3103 VPWR.t5959 VPWR.t1059 129.631
R3104 VPWR.t5333 VPWR.t3760 129.631
R3105 VPWR.t770 VPWR.t3953 129.631
R3106 VPWR.t5537 VPWR.t1122 129.631
R3107 VPWR.t3062 VPWR.t1641 129.631
R3108 VPWR.t2832 VPWR.t7069 129.631
R3109 VPWR.t6103 VPWR.t4518 129.631
R3110 VPWR.t5427 VPWR.t602 129.631
R3111 VPWR.n2065 VPWR.t4625 129.631
R3112 VPWR.t5654 VPWR.n2066 129.631
R3113 VPWR.t2810 VPWR.t2709 129.631
R3114 VPWR.t2365 VPWR.t1511 129.631
R3115 VPWR.n199 VPWR.t1451 129.631
R3116 VPWR.t4838 VPWR.n200 129.631
R3117 VPWR.n201 VPWR.t2995 129.631
R3118 VPWR.t520 VPWR.n202 129.631
R3119 VPWR.n203 VPWR.t3656 129.631
R3120 VPWR.t2925 VPWR.n204 129.631
R3121 VPWR.n205 VPWR.t5166 129.631
R3122 VPWR.t3767 VPWR.n206 129.631
R3123 VPWR.n207 VPWR.t5963 129.631
R3124 VPWR.t3727 VPWR.t3780 129.631
R3125 VPWR.t6301 VPWR.t4894 129.631
R3126 VPWR.t4073 VPWR.t2079 129.631
R3127 VPWR.t1001 VPWR.t2908 129.631
R3128 VPWR.t3846 VPWR.t1178 129.631
R3129 VPWR.t2876 VPWR.t4647 129.631
R3130 VPWR.t1370 VPWR.t5561 129.631
R3131 VPWR.t4034 VPWR.t2938 129.631
R3132 VPWR.t6187 VPWR.t3614 129.631
R3133 VPWR.t2214 VPWR.t4710 129.631
R3134 VPWR.t3043 VPWR.t3458 129.631
R3135 VPWR.t4950 VPWR.t5644 129.631
R3136 VPWR.t3122 VPWR.t5953 129.631
R3137 VPWR.t4825 VPWR.t2221 129.631
R3138 VPWR.t5335 VPWR.t1890 129.631
R3139 VPWR.t3509 VPWR.t4332 129.631
R3140 VPWR.t2443 VPWR.t2251 129.631
R3141 VPWR.t2723 VPWR.t4424 129.631
R3142 VPWR.t1647 VPWR.t4179 129.631
R3143 VPWR.t2819 VPWR.t4727 129.631
R3144 VPWR.t5435 VPWR.t1798 129.631
R3145 VPWR.t2674 VPWR.t1715 129.631
R3146 VPWR.t3556 VPWR.t5945 129.631
R3147 VPWR.t2549 VPWR.t4199 129.631
R3148 VPWR.t3917 VPWR.t4900 129.631
R3149 VPWR.t5731 VPWR.t2013 129.631
R3150 VPWR.t1003 VPWR.t5750 129.631
R3151 VPWR.t4596 VPWR.t4632 129.631
R3152 VPWR.t3963 VPWR.t598 129.631
R3153 VPWR.t2577 VPWR.t6033 129.631
R3154 VPWR.t6033 VPWR.t213 129.631
R3155 VPWR.t3301 VPWR.t195 129.631
R3156 VPWR.t3864 VPWR.t4616 129.631
R3157 VPWR.t2720 VPWR.t3009 129.631
R3158 VPWR.t6358 VPWR.t2984 129.631
R3159 VPWR.t84 VPWR.t5681 129.631
R3160 VPWR.t4022 VPWR.t2327 129.631
R3161 VPWR.t2344 VPWR.t2295 129.631
R3162 VPWR.t885 VPWR.t3198 129.631
R3163 VPWR.n370 VPWR.t4403 129.631
R3164 VPWR.t2321 VPWR.t1575 129.631
R3165 VPWR.t5315 VPWR.t5666 129.631
R3166 VPWR.t3620 VPWR.t1719 129.631
R3167 VPWR.t5348 VPWR.t7075 129.631
R3168 VPWR.t3154 VPWR.t5074 129.631
R3169 VPWR.n373 VPWR.t2511 129.631
R3170 VPWR.t5582 VPWR.t5235 129.631
R3171 VPWR.t3776 VPWR.t2814 129.631
R3172 VPWR.t3403 VPWR.t3548 129.631
R3173 VPWR.n3707 VPWR.t4374 129.631
R3174 VPWR.n267 VPWR.t3894 129.631
R3175 VPWR.n2427 VPWR.t839 129.631
R3176 VPWR.t4771 VPWR.n2428 129.631
R3177 VPWR.n2429 VPWR.t4783 129.631
R3178 VPWR.n262 VPWR.t4618 129.631
R3179 VPWR.t2138 VPWR.n261 129.631
R3180 VPWR.t1779 VPWR.n2535 129.631
R3181 VPWR.n2536 VPWR.t1723 129.631
R3182 VPWR.t629 VPWR.n2537 129.631
R3183 VPWR.n2538 VPWR.t2716 129.631
R3184 VPWR.t1842 VPWR.n2539 129.631
R3185 VPWR.n2540 VPWR.t4898 129.631
R3186 VPWR.n2541 VPWR.t1983 129.631
R3187 VPWR.t758 VPWR.n1 129.631
R3188 VPWR.n10 VPWR.t3936 129.631
R3189 VPWR.n31 VPWR.t2093 129.631
R3190 VPWR.t1877 VPWR.n32 129.631
R3191 VPWR.n33 VPWR.t6294 129.631
R3192 VPWR.t6022 VPWR.n34 129.631
R3193 VPWR.n35 VPWR.t518 129.631
R3194 VPWR.n64 VPWR.t5726 129.631
R3195 VPWR.t1099 VPWR.n63 129.631
R3196 VPWR.t4744 VPWR.n85 129.631
R3197 VPWR.n86 VPWR.t5535 129.631
R3198 VPWR.t662 VPWR.n87 129.631
R3199 VPWR.n88 VPWR.t6010 129.631
R3200 VPWR.t1354 VPWR.t6900 128.472
R3201 VPWR.t568 VPWR.t3910 128.472
R3202 VPWR.t5005 VPWR 128.472
R3203 VPWR VPWR.t4797 128.472
R3204 VPWR.t6629 VPWR.t5933 127.316
R3205 VPWR.t4387 VPWR.t4082 127.316
R3206 VPWR.t6975 VPWR.t6537 127.316
R3207 VPWR VPWR.t3398 126.341
R3208 VPWR VPWR.t2335 126.157
R3209 VPWR.t2437 VPWR.t2680 126.157
R3210 VPWR.t6729 VPWR 126.157
R3211 VPWR.t3471 VPWR 126.157
R3212 VPWR.t6292 VPWR 126.157
R3213 VPWR.t3870 VPWR 126.157
R3214 VPWR.t6950 VPWR.t5880 126.157
R3215 VPWR.t6288 VPWR.t569 126.157
R3216 VPWR VPWR.t7112 125.15
R3217 VPWR VPWR.t6709 125.15
R3218 VPWR.t6097 VPWR.t6894 125.001
R3219 VPWR.t6973 VPWR.t2354 125.001
R3220 VPWR.t3484 VPWR.t46 125.001
R3221 VPWR.t7023 VPWR.t2499 125.001
R3222 VPWR.t4203 VPWR.t6470 125.001
R3223 VPWR.t6593 VPWR 125.001
R3224 VPWR.t5672 VPWR.t5539 125.001
R3225 VPWR.t6500 VPWR.t3001 123.957
R3226 VPWR.t16 VPWR.t3007 123.957
R3227 VPWR.t235 VPWR.t4681 123.957
R3228 VPWR.t289 VPWR.t33 123.957
R3229 VPWR.t2283 VPWR 123.844
R3230 VPWR VPWR.t1668 123.844
R3231 VPWR.t6797 VPWR.t3018 123.073
R3232 VPWR.t1360 VPWR.t5260 122.686
R3233 VPWR.t2608 VPWR 122.686
R3234 VPWR VPWR.t3752 122.686
R3235 VPWR VPWR.t2837 122.686
R3236 VPWR.t4359 VPWR 122.686
R3237 VPWR VPWR.t3827 122.686
R3238 VPWR.t1322 VPWR 122.686
R3239 VPWR.t4818 VPWR.n3262 122.686
R3240 VPWR.t4365 VPWR 122.686
R3241 VPWR.t5998 VPWR 122.686
R3242 VPWR VPWR.t6726 122.686
R3243 VPWR VPWR.t6429 122.686
R3244 VPWR.t4421 VPWR.t1993 122.686
R3245 VPWR.t4708 VPWR.t5913 122.686
R3246 VPWR VPWR.t4830 122.686
R3247 VPWR.t7022 VPWR.t2396 122.686
R3248 VPWR.t6243 VPWR.t5408 122.686
R3249 VPWR.t7010 VPWR.t2123 122.686
R3250 VPWR.t303 VPWR 122.686
R3251 VPWR.t958 VPWR 122.686
R3252 VPWR VPWR.t6286 122.686
R3253 VPWR VPWR.t2586 121.528
R3254 VPWR.t1161 VPWR 121.528
R3255 VPWR.t4881 VPWR 121.528
R3256 VPWR.t106 VPWR 121.528
R3257 VPWR.t5718 VPWR 121.528
R3258 VPWR.t1212 VPWR 121.528
R3259 VPWR.t2569 VPWR 121.528
R3260 VPWR.t1741 VPWR 121.528
R3261 VPWR.t3789 VPWR 121.528
R3262 VPWR.t4868 VPWR 121.528
R3263 VPWR VPWR.t5935 121.528
R3264 VPWR.t2237 VPWR 121.528
R3265 VPWR.t6793 VPWR 121.528
R3266 VPWR.t7014 VPWR 121.528
R3267 VPWR.t323 VPWR 121.528
R3268 VPWR VPWR.t2655 121.528
R3269 VPWR VPWR.t4600 121.528
R3270 VPWR VPWR.t6278 121.528
R3271 VPWR.t5039 VPWR 121.528
R3272 VPWR.t2768 VPWR 121.528
R3273 VPWR VPWR.t6702 121.528
R3274 VPWR.t6515 VPWR 121.528
R3275 VPWR.t6517 VPWR 121.528
R3276 VPWR.t7054 VPWR.t6333 121.528
R3277 VPWR VPWR.t614 121.528
R3278 VPWR.t793 VPWR 121.528
R3279 VPWR.t3277 VPWR 121.528
R3280 VPWR VPWR.t1940 121.528
R3281 VPWR.t2273 VPWR 121.528
R3282 VPWR.t5722 VPWR 121.528
R3283 VPWR.t3710 VPWR 121.528
R3284 VPWR.t4381 VPWR 121.528
R3285 VPWR.t920 VPWR 121.528
R3286 VPWR VPWR.t4864 121.528
R3287 VPWR VPWR.t3095 121.528
R3288 VPWR.t3150 VPWR 121.528
R3289 VPWR.t3835 VPWR 121.528
R3290 VPWR VPWR.t1954 121.528
R3291 VPWR.t1426 VPWR 121.528
R3292 VPWR.t225 VPWR.t217 121.528
R3293 VPWR VPWR.t4224 121.528
R3294 VPWR VPWR.t6808 121.528
R3295 VPWR VPWR.t5622 121.528
R3296 VPWR.t2183 VPWR 121.528
R3297 VPWR.t1103 VPWR 121.528
R3298 VPWR.t2277 VPWR 121.528
R3299 VPWR VPWR.t2485 121.528
R3300 VPWR VPWR.t3890 121.528
R3301 VPWR VPWR.t6061 121.528
R3302 VPWR.t2223 VPWR 121.528
R3303 VPWR.t6059 VPWR 121.528
R3304 VPWR VPWR.t6633 121.528
R3305 VPWR.t2746 VPWR 121.528
R3306 VPWR.t4833 VPWR 121.528
R3307 VPWR VPWR.t5846 121.528
R3308 VPWR VPWR.t6732 121.528
R3309 VPWR VPWR.t6525 121.528
R3310 VPWR.t479 VPWR 121.528
R3311 VPWR.t6213 VPWR 121.528
R3312 VPWR.t474 VPWR 121.528
R3313 VPWR.t2954 VPWR 121.528
R3314 VPWR.t4201 VPWR 121.528
R3315 VPWR.t6424 VPWR 121.528
R3316 VPWR VPWR.t3568 121.528
R3317 VPWR.t5118 VPWR 121.528
R3318 VPWR VPWR.t841 121.528
R3319 VPWR.t7105 VPWR 121.528
R3320 VPWR VPWR.t4477 121.528
R3321 VPWR.t4483 VPWR 121.528
R3322 VPWR VPWR.t6174 121.528
R3323 VPWR.t904 VPWR 121.528
R3324 VPWR VPWR.t1077 121.528
R3325 VPWR.t3586 VPWR 121.528
R3326 VPWR VPWR.t5410 121.528
R3327 VPWR VPWR.t2398 121.528
R3328 VPWR.t1686 VPWR 121.528
R3329 VPWR VPWR.t4719 121.528
R3330 VPWR.t3058 VPWR 121.528
R3331 VPWR.t1318 VPWR 121.528
R3332 VPWR.t1316 VPWR 121.528
R3333 VPWR VPWR.t1050 121.528
R3334 VPWR.t1587 VPWR 121.528
R3335 VPWR VPWR.t5254 121.528
R3336 VPWR.t6599 VPWR 121.528
R3337 VPWR VPWR.t6607 121.528
R3338 VPWR.t6373 VPWR 121.528
R3339 VPWR.t3772 VPWR 121.528
R3340 VPWR VPWR.t895 121.528
R3341 VPWR.t257 VPWR 121.528
R3342 VPWR.t247 VPWR 121.528
R3343 VPWR VPWR.t6825 121.528
R3344 VPWR.t189 VPWR 121.528
R3345 VPWR VPWR.t2525 121.528
R3346 VPWR.t3736 VPWR 121.528
R3347 VPWR.t5909 VPWR 121.528
R3348 VPWR VPWR.t4508 121.528
R3349 VPWR.t1859 VPWR 121.528
R3350 VPWR VPWR.t1682 121.528
R3351 VPWR VPWR.t6166 121.528
R3352 VPWR.t5613 VPWR 121.528
R3353 VPWR VPWR.t1387 121.528
R3354 VPWR VPWR.t5885 121.528
R3355 VPWR.t6131 VPWR 121.528
R3356 VPWR VPWR.t2999 121.528
R3357 VPWR.t6254 VPWR 121.528
R3358 VPWR.t2369 VPWR 121.528
R3359 VPWR.t5889 VPWR 121.528
R3360 VPWR VPWR.t3072 121.528
R3361 VPWR VPWR.t5692 121.528
R3362 VPWR VPWR.t2119 121.528
R3363 VPWR.t5571 VPWR 121.528
R3364 VPWR VPWR.t5601 121.528
R3365 VPWR.t4550 VPWR 121.528
R3366 VPWR.t3172 VPWR 121.528
R3367 VPWR.t2208 VPWR 121.528
R3368 VPWR VPWR.t1405 121.528
R3369 VPWR VPWR.t2202 121.528
R3370 VPWR VPWR.t4531 121.528
R3371 VPWR VPWR.t1603 121.528
R3372 VPWR VPWR.t1124 121.528
R3373 VPWR.t608 VPWR 121.528
R3374 VPWR VPWR.t5991 121.528
R3375 VPWR VPWR.t1118 121.528
R3376 VPWR VPWR.t5951 121.528
R3377 VPWR.t6391 VPWR 121.528
R3378 VPWR VPWR.t1368 121.528
R3379 VPWR.t966 VPWR 121.528
R3380 VPWR VPWR.t5133 121.528
R3381 VPWR.t4649 VPWR 121.528
R3382 VPWR VPWR.t4062 121.528
R3383 VPWR.t3571 VPWR 121.528
R3384 VPWR VPWR.t2363 121.528
R3385 VPWR VPWR.t1513 121.528
R3386 VPWR.t1517 VPWR 121.528
R3387 VPWR VPWR.t3397 121.528
R3388 VPWR VPWR.t3351 121.528
R3389 VPWR.t6886 VPWR 121.528
R3390 VPWR VPWR.t3346 121.528
R3391 VPWR VPWR.t6591 121.528
R3392 VPWR.t132 VPWR 121.528
R3393 VPWR VPWR.t4134 121.528
R3394 VPWR VPWR.t6706 121.528
R3395 VPWR.t5997 VPWR 121.528
R3396 VPWR VPWR.t6315 121.528
R3397 VPWR.t2826 VPWR 121.528
R3398 VPWR VPWR.t2828 121.528
R3399 VPWR.t750 VPWR 121.528
R3400 VPWR VPWR.t3114 121.528
R3401 VPWR VPWR.t4498 121.528
R3402 VPWR VPWR.t2869 121.528
R3403 VPWR.t1731 VPWR 121.528
R3404 VPWR VPWR.t1727 121.528
R3405 VPWR VPWR.t4721 121.528
R3406 VPWR.t3988 VPWR 121.528
R3407 VPWR.t3336 VPWR 121.528
R3408 VPWR VPWR.t5607 121.528
R3409 VPWR VPWR.t1708 121.528
R3410 VPWR.t5176 VPWR 121.528
R3411 VPWR.t5665 VPWR 121.528
R3412 VPWR.t2706 VPWR 121.528
R3413 VPWR.t2575 VPWR 121.528
R3414 VPWR VPWR.t7032 121.528
R3415 VPWR.t6390 VPWR 121.528
R3416 VPWR.t4802 VPWR 121.528
R3417 VPWR.t3120 VPWR 121.528
R3418 VPWR VPWR.t5072 121.528
R3419 VPWR VPWR.t3152 121.528
R3420 VPWR.t5784 VPWR 121.528
R3421 VPWR VPWR.t2861 121.528
R3422 VPWR.t5492 VPWR 121.528
R3423 VPWR.t3068 VPWR 121.528
R3424 VPWR.t4322 VPWR 121.528
R3425 VPWR.t1932 VPWR.t3217 120.371
R3426 VPWR.t799 VPWR.t2031 120.371
R3427 VPWR.t7002 VPWR.t6784 120.371
R3428 VPWR.t5144 VPWR.t6777 120.371
R3429 VPWR.t5805 VPWR.t6859 120.371
R3430 VPWR.t6488 VPWR.t3162 120.371
R3431 VPWR.t1794 VPWR.t6570 120.371
R3432 VPWR VPWR.t6720 119.213
R3433 VPWR.t4397 VPWR.t6675 118.056
R3434 VPWR.t5662 VPWR.t1111 118.056
R3435 VPWR.t3416 VPWR.t1625 118.056
R3436 VPWR.t2231 VPWR.t6101 118.056
R3437 VPWR.t906 VPWR.t2261 118.056
R3438 VPWR.t6510 VPWR.t6985 118.056
R3439 VPWR.t2595 VPWR.t6245 118.056
R3440 VPWR.t5565 VPWR.t1846 118.056
R3441 VPWR.t1597 VPWR.t1563 118.056
R3442 VPWR VPWR.t2949 117.859
R3443 VPWR.t6865 VPWR.t1031 116.898
R3444 VPWR.t5584 VPWR.t2654 115.742
R3445 VPWR.t6945 VPWR 115.742
R3446 VPWR VPWR.t6907 115.742
R3447 VPWR.t105 VPWR 115.742
R3448 VPWR.t2031 VPWR.t795 115.742
R3449 VPWR.t6784 VPWR.t799 115.742
R3450 VPWR.t6728 VPWR.t5805 115.742
R3451 VPWR.t7039 VPWR.t3950 115.742
R3452 VPWR.t3825 VPWR.t4219 115.742
R3453 VPWR.t4698 VPWR.t6504 115.742
R3454 VPWR.t4224 VPWR.t5305 115.742
R3455 VPWR.t6372 VPWR 115.742
R3456 VPWR.t3162 VPWR.t37 115.742
R3457 VPWR VPWR.t40 115.742
R3458 VPWR.t4719 VPWR.t3058 115.742
R3459 VPWR.t1050 VPWR.t1587 115.742
R3460 VPWR.t6943 VPWR.t5701 115.742
R3461 VPWR VPWR.t93 115.742
R3462 VPWR.t6315 VPWR.t2826 115.742
R3463 VPWR VPWR.t4075 114.584
R3464 VPWR.t2657 VPWR 114.584
R3465 VPWR VPWR.t5923 114.584
R3466 VPWR VPWR.t5919 114.584
R3467 VPWR VPWR.t6998 114.584
R3468 VPWR VPWR.t5475 114.584
R3469 VPWR.t522 VPWR.t225 114.584
R3470 VPWR.t217 VPWR.t4359 114.584
R3471 VPWR.t6952 VPWR 114.584
R3472 VPWR.t3960 VPWR.t3930 114.584
R3473 VPWR.t6620 VPWR 114.584
R3474 VPWR.t5391 VPWR 114.584
R3475 VPWR VPWR.t5567 114.584
R3476 VPWR.t6641 VPWR 114.584
R3477 VPWR VPWR.t1034 113.427
R3478 VPWR.t4958 VPWR.n923 113.427
R3479 VPWR.t7005 VPWR 113.427
R3480 VPWR.t2918 VPWR.t285 113.427
R3481 VPWR.t5589 VPWR.n604 113.427
R3482 VPWR.t6929 VPWR.n612 113.427
R3483 VPWR.t6923 VPWR.t2541 113.427
R3484 VPWR.t6915 VPWR.t1788 113.427
R3485 VPWR.t2734 VPWR.t6097 111.112
R3486 VPWR.t95 VPWR.t6768 111.112
R3487 VPWR.t1256 VPWR.t612 111.112
R3488 VPWR.t2354 VPWR.t6964 111.112
R3489 VPWR.t46 VPWR.t6973 111.112
R3490 VPWR.t2499 VPWR.t3880 111.112
R3491 VPWR.t7013 VPWR.t7023 111.112
R3492 VPWR.t1021 VPWR.t2477 111.112
R3493 VPWR.t6337 VPWR.t6681 111.112
R3494 VPWR.t3840 VPWR.t6560 111.112
R3495 VPWR.t6617 VPWR.t6562 111.112
R3496 VPWR.t5961 VPWR.t6558 111.112
R3497 VPWR.t29 VPWR.t275 111.112
R3498 VPWR VPWR.t6604 111.112
R3499 VPWR.t1266 VPWR.t6616 111.112
R3500 VPWR.t3942 VPWR.t5176 111.112
R3501 VPWR.t437 VPWR.t4322 111.112
R3502 VPWR.t2680 VPWR.t2439 109.954
R3503 VPWR.t819 VPWR 109.954
R3504 VPWR VPWR.t3868 109.954
R3505 VPWR.t569 VPWR.t6950 109.954
R3506 VPWR.t2021 VPWR 109.954
R3507 VPWR.t6264 VPWR 109.954
R3508 VPWR.t4460 VPWR.t6414 109.954
R3509 VPWR.t1907 VPWR 109.954
R3510 VPWR.t5933 VPWR.t6874 108.796
R3511 VPWR.t4247 VPWR.t4255 108.796
R3512 VPWR.t4087 VPWR.t4387 108.796
R3513 VPWR.t4251 VPWR.t6320 108.796
R3514 VPWR.t6537 VPWR.t6977 108.796
R3515 VPWR.n833 VPWR.t910 108.796
R3516 VPWR.t5342 VPWR.t5507 108.796
R3517 VPWR.t4747 VPWR.t6153 108.796
R3518 VPWR.t5642 VPWR.t6220 108.796
R3519 VPWR.t2342 VPWR.t1694 108.796
R3520 VPWR.t1019 VPWR.t6248 108.796
R3521 VPWR VPWR.t7134 107.639
R3522 VPWR.t2435 VPWR 107.639
R3523 VPWR VPWR.t7060 107.639
R3524 VPWR VPWR.t3598 107.639
R3525 VPWR.t3097 VPWR 107.639
R3526 VPWR VPWR.t6869 107.639
R3527 VPWR VPWR.t3507 107.639
R3528 VPWR.t5620 VPWR 107.639
R3529 VPWR VPWR.t2181 107.639
R3530 VPWR VPWR.t2744 107.639
R3531 VPWR.t774 VPWR 107.639
R3532 VPWR.t6863 VPWR 107.639
R3533 VPWR VPWR.t208 107.639
R3534 VPWR VPWR.t946 107.639
R3535 VPWR.t3568 VPWR.t568 107.639
R3536 VPWR.t2023 VPWR 107.639
R3537 VPWR.t843 VPWR 107.639
R3538 VPWR.t5412 VPWR 107.639
R3539 VPWR VPWR.t273 107.639
R3540 VPWR.t6842 VPWR 107.639
R3541 VPWR.t1585 VPWR 107.639
R3542 VPWR VPWR.t3974 107.639
R3543 VPWR VPWR.t5889 107.639
R3544 VPWR.t5694 VPWR 107.639
R3545 VPWR.t210 VPWR 107.639
R3546 VPWR VPWR.t4792 107.639
R3547 VPWR VPWR.t5159 107.639
R3548 VPWR VPWR.t939 107.639
R3549 VPWR.t4465 VPWR 107.639
R3550 VPWR VPWR.t2824 107.639
R3551 VPWR.t6313 VPWR 107.639
R3552 VPWR.t4498 VPWR 107.639
R3553 VPWR.t4723 VPWR 107.639
R3554 VPWR VPWR.t2600 107.639
R3555 VPWR VPWR.t6596 107.639
R3556 VPWR VPWR.t214 107.639
R3557 VPWR.t4840 VPWR 107.639
R3558 VPWR VPWR.t2502 107.639
R3559 VPWR.t2863 VPWR 107.639
R3560 VPWR VPWR.t6415 107.639
R3561 VPWR.t3531 VPWR.t6790 106.481
R3562 VPWR.t2152 VPWR.t5268 106.481
R3563 VPWR.t4604 VPWR.t6276 106.481
R3564 VPWR.t4185 VPWR.t6682 106.481
R3565 VPWR.t4187 VPWR.t6692 106.481
R3566 VPWR.t6669 VPWR.t3637 106.481
R3567 VPWR VPWR.t4851 106.481
R3568 VPWR VPWR.t6639 106.481
R3569 VPWR.t187 VPWR.t6766 106.481
R3570 VPWR VPWR.t3267 106.481
R3571 VPWR.t3473 VPWR.t6213 106.481
R3572 VPWR.t4207 VPWR.t4209 106.481
R3573 VPWR.t2648 VPWR.t224 106.481
R3574 VPWR.t3771 VPWR.t3301 106.481
R3575 VPWR VPWR.t4464 106.481
R3576 VPWR VPWR.t6379 105.325
R3577 VPWR.t6715 VPWR.t4998 105.325
R3578 VPWR.t7056 VPWR.t3481 104.168
R3579 VPWR.t6738 VPWR.t6736 104.168
R3580 VPWR.t480 VPWR.t3357 104.168
R3581 VPWR.t2158 VPWR.t21 103.01
R3582 VPWR.t7058 VPWR 103.01
R3583 VPWR VPWR.t4816 103.01
R3584 VPWR.t973 VPWR.t5599 103.01
R3585 VPWR.t2164 VPWR.t201 103.01
R3586 VPWR.t2805 VPWR.t237 103.01
R3587 VPWR VPWR.t1911 103.01
R3588 VPWR VPWR.t6960 103.01
R3589 VPWR VPWR.t3273 103.01
R3590 VPWR.t4463 VPWR.t6417 103.01
R3591 VPWR.t5218 VPWR.t1161 101.853
R3592 VPWR.t7136 VPWR.t96 101.853
R3593 VPWR.t3529 VPWR.t6779 101.853
R3594 VPWR.t2348 VPWR.t5485 101.853
R3595 VPWR.t1411 VPWR.t6856 101.853
R3596 VPWR.t4234 VPWR.t2487 101.853
R3597 VPWR.t5846 VPWR.t2257 101.853
R3598 VPWR.t3308 VPWR.t2259 101.853
R3599 VPWR.t206 VPWR.t2066 101.853
R3600 VPWR.t1515 VPWR.t4665 101.853
R3601 VPWR.t5003 VPWR.t5996 101.853
R3602 VPWR.t2702 VPWR.t2900 101.853
R3603 VPWR.t300 VPWR.t2737 101.853
R3604 VPWR.t3460 VPWR.n371 101.853
R3605 VPWR.t3118 VPWR.t2874 101.853
R3606 VPWR VPWR.t6538 101.311
R3607 VPWR.t910 VPWR 100.695
R3608 VPWR.t2966 VPWR.t6678 100.695
R3609 VPWR.t239 VPWR.t5587 100.695
R3610 VPWR VPWR.t2930 100.695
R3611 VPWR.t27 VPWR.t936 100.695
R3612 VPWR.t2027 VPWR.t5144 100.445
R3613 VPWR.t20 VPWR.t3005 100.12
R3614 VPWR.t241 VPWR.t4694 100.12
R3615 VPWR.t293 VPWR.t31 100.12
R3616 VPWR.t291 VPWR.t4697 100.12
R3617 VPWR.t6341 VPWR.t3791 99.5375
R3618 VPWR.t7064 VPWR.t2150 99.5375
R3619 VPWR.t3882 VPWR.t3505 99.5375
R3620 VPWR.t7017 VPWR 99.5375
R3621 VPWR.t6724 VPWR.t4226 99.5375
R3622 VPWR.n756 VPWR.t819 99.5375
R3623 VPWR.n128 VPWR.t2350 99.5375
R3624 VPWR.n1783 VPWR.t2021 99.5375
R3625 VPWR.t283 VPWR.t3307 99.5375
R3626 VPWR.t3848 VPWR.t4527 99.5375
R3627 VPWR.t231 VPWR.t5438 99.5375
R3628 VPWR.t3251 VPWR.t1849 99.5375
R3629 VPWR.t4842 VPWR.t5825 99.5375
R3630 VPWR.t1488 VPWR.t2500 99.5375
R3631 VPWR VPWR.t5138 98.9278
R3632 VPWR.t3016 VPWR 98.9278
R3633 VPWR.t6854 VPWR 98.3801
R3634 VPWR VPWR.t788 98.3801
R3635 VPWR.t6986 VPWR.t7109 98.3801
R3636 VPWR.t4558 VPWR.t6970 98.3801
R3637 VPWR.t6968 VPWR.t4561 98.3801
R3638 VPWR VPWR.t6422 98.3801
R3639 VPWR.t3754 VPWR.t4 97.2227
R3640 VPWR.t6216 VPWR.t5039 97.2227
R3641 VPWR.t6548 VPWR.t123 97.2227
R3642 VPWR.t1331 VPWR.t1847 97.2227
R3643 VPWR.t3018 VPWR.t6716 97.2227
R3644 VPWR.t1262 VPWR.t907 96.9562
R3645 VPWR.t6873 VPWR.t2481 96.1416
R3646 VPWR VPWR.t3839 96.0653
R3647 VPWR VPWR.t6862 96.0653
R3648 VPWR VPWR.t4687 96.0653
R3649 VPWR VPWR.t6546 96.0653
R3650 VPWR VPWR.t5589 96.0653
R3651 VPWR.t1326 VPWR 96.0653
R3652 VPWR VPWR.t6582 96.0653
R3653 VPWR VPWR.t6631 94.9079
R3654 VPWR.n1389 VPWR.t2659 94.9079
R3655 VPWR.t5919 VPWR.n920 94.9079
R3656 VPWR.t2325 VPWR.t6494 94.9079
R3657 VPWR.t1698 VPWR.t6476 94.9079
R3658 VPWR.t5216 VPWR.t6484 94.9079
R3659 VPWR.t3633 VPWR.t6094 94.9079
R3660 VPWR.t6754 VPWR.t4043 94.9079
R3661 VPWR.t1995 VPWR.t6464 94.9079
R3662 VPWR.t6746 VPWR.t2176 94.9079
R3663 VPWR.t305 VPWR.t1280 94.9079
R3664 VPWR.t2646 VPWR.t2634 94.9079
R3665 VPWR.n385 VPWR.t136 94.9079
R3666 VPWR.t6982 VPWR.t6752 93.9328
R3667 VPWR.t897 VPWR.t1130 93.7505
R3668 VPWR.t6576 VPWR.t5730 93.7505
R3669 VPWR.t2652 VPWR.t5815 92.5931
R3670 VPWR.t1288 VPWR.t6599 92.5931
R3671 VPWR.t19 VPWR.t245 92.5931
R3672 VPWR VPWR.t1478 91.4357
R3673 VPWR.t5813 VPWR.t6418 91.4357
R3674 VPWR.t2004 VPWR.t303 91.4357
R3675 VPWR.t3413 VPWR.t4084 90.2783
R3676 VPWR.t3826 VPWR.t4228 89.1209
R3677 VPWR.n742 VPWR.n735 89.1209
R3678 VPWR.n392 VPWR.t7031 88.2007
R3679 VPWR.t5660 VPWR.t1107 87.9635
R3680 VPWR.t1690 VPWR.t6688 87.9635
R3681 VPWR.t7055 VPWR.t6791 87.9635
R3682 VPWR.t4220 VPWR.t908 87.9635
R3683 VPWR.t6501 VPWR.t3949 87.9635
R3684 VPWR.t4692 VPWR.t12 87.9635
R3685 VPWR.t6529 VPWR.t3992 87.9635
R3686 VPWR.t948 VPWR.t2954 87.9635
R3687 VPWR.t5855 VPWR.t6988 87.9635
R3688 VPWR.t191 VPWR.t6566 87.9635
R3689 VPWR.t295 VPWR.t125 87.9635
R3690 VPWR.t6806 VPWR.t134 87.9635
R3691 VPWR.t186 VPWR.t183 87.9635
R3692 VPWR.t6015 VPWR.t56 87.9635
R3693 VPWR.t1751 VPWR.t6395 87.9635
R3694 VPWR.t464 VPWR.t198 86.823
R3695 VPWR VPWR.t5422 86.8061
R3696 VPWR.t1046 VPWR.t7034 86.8061
R3697 VPWR.t137 VPWR.n964 85.6486
R3698 VPWR.n953 VPWR.t157 85.6486
R3699 VPWR.n946 VPWR.t6866 85.6486
R3700 VPWR.n934 VPWR.t95 85.6486
R3701 VPWR.t1532 VPWR.t4872 85.6486
R3702 VPWR.n928 VPWR.t7055 85.6486
R3703 VPWR.t3449 VPWR.t3669 85.6486
R3704 VPWR.n3358 VPWR.t6908 85.6486
R3705 VPWR.t104 VPWR.n114 85.6486
R3706 VPWR.n845 VPWR.t6615 85.6486
R3707 VPWR.t1942 VPWR.t3277 85.6486
R3708 VPWR.t1940 VPWR.t3279 85.6486
R3709 VPWR.t4866 VPWR.t920 85.6486
R3710 VPWR.t4864 VPWR.t918 85.6486
R3711 VPWR.n827 VPWR.t7099 85.6486
R3712 VPWR.n3273 VPWR.t6382 85.6486
R3713 VPWR.n3268 VPWR.t7004 85.6486
R3714 VPWR.t177 VPWR.n749 85.6486
R3715 VPWR.t5092 VPWR.t5462 85.6486
R3716 VPWR.n3261 VPWR.t6337 85.6486
R3717 VPWR.n156 VPWR.t7029 85.6486
R3718 VPWR.n141 VPWR.t39 85.6486
R3719 VPWR.t6399 VPWR.n1782 85.6486
R3720 VPWR.t4479 VPWR.t7105 85.6486
R3721 VPWR.t4477 VPWR.t7103 85.6486
R3722 VPWR.t6172 VPWR.t4483 85.6486
R3723 VPWR.t6174 VPWR.t4481 85.6486
R3724 VPWR.t1079 VPWR.t904 85.6486
R3725 VPWR.t1077 VPWR.t902 85.6486
R3726 VPWR.t28 VPWR.n1092 85.6486
R3727 VPWR.n2879 VPWR.t6942 85.6486
R3728 VPWR.n2880 VPWR.t90 85.6486
R3729 VPWR.t162 VPWR.n2748 85.6486
R3730 VPWR.t101 VPWR.n175 85.6486
R3731 VPWR.t2949 VPWR.n181 85.6486
R3732 VPWR.n2952 VPWR.t49 85.6486
R3733 VPWR.t6414 VPWR.n377 85.6486
R3734 VPWR VPWR.t145 84.4912
R3735 VPWR.t6631 VPWR.n1385 84.4912
R3736 VPWR VPWR.t6758 84.4912
R3737 VPWR.t6704 VPWR 84.4912
R3738 VPWR.t6618 VPWR 84.4912
R3739 VPWR VPWR.t3633 84.4912
R3740 VPWR.t6653 VPWR 84.4912
R3741 VPWR.t1583 VPWR 84.4912
R3742 VPWR.t3932 VPWR 84.4912
R3743 VPWR.t7094 VPWR.t1909 83.3338
R3744 VPWR.t3833 VPWR.t6178 83.3338
R3745 VPWR.t6791 VPWR.t4655 83.3338
R3746 VPWR.t4687 VPWR.t1785 83.3338
R3747 VPWR.t6857 VPWR.t2166 83.3338
R3748 VPWR.t215 VPWR.t7115 83.3338
R3749 VPWR.t6885 VPWR.t6168 83.3338
R3750 VPWR.t7025 VPWR 82.1764
R3751 VPWR.t2170 VPWR.t5014 81.019
R3752 VPWR.t5395 VPWR.t6040 81.019
R3753 VPWR.t1599 VPWR.t6044 81.019
R3754 VPWR.t5237 VPWR.t401 81.019
R3755 VPWR.t6260 VPWR.t399 81.019
R3756 VPWR.t4557 VPWR.n3255 81.019
R3757 VPWR.t1787 VPWR.t6915 81.019
R3758 VPWR.t4117 VPWR 79.8616
R3759 VPWR VPWR.t4258 79.8616
R3760 VPWR VPWR.t2799 79.8616
R3761 VPWR VPWR.t4470 79.8616
R3762 VPWR VPWR.t754 79.8616
R3763 VPWR.t6446 VPWR 79.8616
R3764 VPWR VPWR.t5656 79.8616
R3765 VPWR.t7037 VPWR.n819 79.8616
R3766 VPWR.t5214 VPWR 79.8616
R3767 VPWR.t342 VPWR 79.8616
R3768 VPWR.n1229 VPWR 79.8616
R3769 VPWR VPWR.t934 79.8616
R3770 VPWR VPWR.t715 79.8616
R3771 VPWR VPWR.t5468 79.8616
R3772 VPWR VPWR.t2588 79.8616
R3773 VPWR.t2588 VPWR 79.8616
R3774 VPWR.n1779 VPWR 79.8616
R3775 VPWR VPWR.n1779 79.8616
R3776 VPWR VPWR.t683 79.8616
R3777 VPWR VPWR.t5070 79.8616
R3778 VPWR.t582 VPWR 79.8616
R3779 VPWR.t1535 VPWR 79.8616
R3780 VPWR.t5151 VPWR 79.8616
R3781 VPWR.t5110 VPWR 79.8616
R3782 VPWR.t1627 VPWR 79.8616
R3783 VPWR.t5844 VPWR 79.8616
R3784 VPWR.t6327 VPWR 79.8616
R3785 VPWR VPWR.t1310 79.8616
R3786 VPWR VPWR.n2318 79.8616
R3787 VPWR VPWR.t3769 79.8616
R3788 VPWR VPWR.t4768 79.8616
R3789 VPWR VPWR.t6311 79.8616
R3790 VPWR.t5205 VPWR 79.8616
R3791 VPWR.t5899 VPWR 79.8616
R3792 VPWR.t999 VPWR 79.8616
R3793 VPWR.t3087 VPWR 79.8616
R3794 VPWR.t5688 VPWR 79.8616
R3795 VPWR.t4625 VPWR 79.8616
R3796 VPWR VPWR.n198 79.8616
R3797 VPWR.t2263 VPWR 79.8616
R3798 VPWR.t5223 VPWR 79.8616
R3799 VPWR.t1451 VPWR 79.8616
R3800 VPWR.t2995 VPWR 79.8616
R3801 VPWR.t3656 VPWR 79.8616
R3802 VPWR.t5166 VPWR 79.8616
R3803 VPWR.t3652 VPWR 79.8616
R3804 VPWR.t5963 VPWR 79.8616
R3805 VPWR.t4269 VPWR 79.8616
R3806 VPWR.n525 VPWR 79.8616
R3807 VPWR VPWR.t5444 79.8616
R3808 VPWR VPWR.t5402 79.8616
R3809 VPWR VPWR.n180 79.8616
R3810 VPWR VPWR.t4563 79.8616
R3811 VPWR.n381 VPWR 79.8616
R3812 VPWR VPWR.n381 79.8616
R3813 VPWR VPWR.t1181 79.8616
R3814 VPWR VPWR.t4403 79.8616
R3815 VPWR.t4823 VPWR 79.8616
R3816 VPWR.t1372 VPWR 79.8616
R3817 VPWR.t1057 VPWR 79.8616
R3818 VPWR VPWR.t1057 79.8616
R3819 VPWR.t2511 VPWR 79.8616
R3820 VPWR VPWR.t5295 79.8616
R3821 VPWR VPWR.t4374 79.8616
R3822 VPWR VPWR.t845 79.8616
R3823 VPWR.t4488 VPWR 79.8616
R3824 VPWR.t1753 VPWR 79.8616
R3825 VPWR.t2812 VPWR 79.8616
R3826 VPWR.t839 VPWR 79.8616
R3827 VPWR.t4175 VPWR 79.8616
R3828 VPWR.t4783 VPWR 79.8616
R3829 VPWR VPWR.t2138 79.8616
R3830 VPWR.t1723 VPWR 79.8616
R3831 VPWR.t4752 VPWR 79.8616
R3832 VPWR.t2716 VPWR 79.8616
R3833 VPWR.t4898 VPWR 79.8616
R3834 VPWR VPWR.t758 79.8616
R3835 VPWR VPWR.t3258 79.8616
R3836 VPWR VPWR.t2093 79.8616
R3837 VPWR.t6294 VPWR 79.8616
R3838 VPWR.t518 VPWR 79.8616
R3839 VPWR VPWR.t1099 79.8616
R3840 VPWR.t5535 VPWR 79.8616
R3841 VPWR.t6205 VPWR 79.8616
R3842 VPWR.t6010 VPWR 79.8616
R3843 VPWR.t3628 VPWR.n3268 79.1715
R3844 VPWR.t2622 VPWR.n3273 79.1216
R3845 VPWR.t3091 VPWR.n634 79.1216
R3846 VPWR.t5231 VPWR.t4881 78.7042
R3847 VPWR.t3409 VPWR.t2483 78.7042
R3848 VPWR.t671 VPWR.t6331 78.7042
R3849 VPWR.t3221 VPWR.t2637 78.7042
R3850 VPWR.t1761 VPWR.t1763 78.7042
R3851 VPWR.t2331 VPWR.t2240 78.7042
R3852 VPWR.t4012 VPWR.t219 78.7042
R3853 VPWR.t1923 VPWR.t2076 78.7042
R3854 VPWR.t35 VPWR 77.7984
R3855 VPWR VPWR.t1526 77.5468
R3856 VPWR.t1530 VPWR 77.5468
R3857 VPWR VPWR.t2275 77.5468
R3858 VPWR.t1048 VPWR 77.5468
R3859 VPWR VPWR.t5611 77.5468
R3860 VPWR VPWR.t6002 77.5468
R3861 VPWR.t5125 VPWR 77.5468
R3862 VPWR.t3112 VPWR 77.5468
R3863 VPWR VPWR.t4608 77.5468
R3864 VPWR.t4142 VPWR 77.5468
R3865 VPWR VPWR.t510 77.5468
R3866 VPWR.t6164 VPWR 77.5468
R3867 VPWR VPWR.t5189 77.5468
R3868 VPWR.t504 VPWR 77.5468
R3869 VPWR VPWR.t2602 77.5468
R3870 VPWR.t3424 VPWR 77.5468
R3871 VPWR VPWR.t3460 77.5468
R3872 VPWR.t6846 VPWR 77.4737
R3873 VPWR.n1406 VPWR.t7058 76.3894
R3874 VPWR.t7040 VPWR.t3124 76.3894
R3875 VPWR.t5615 VPWR.t2622 76.3894
R3876 VPWR.t4816 VPWR.t3628 76.3894
R3877 VPWR.n735 VPWR.t3283 76.3894
R3878 VPWR.t7117 VPWR.t220 76.3894
R3879 VPWR.t171 VPWR.t6474 76.3894
R3880 VPWR.t371 VPWR.t6776 76.3894
R3881 VPWR.t1911 VPWR.t3091 76.3894
R3882 VPWR.n632 VPWR.t153 76.3894
R3883 VPWR.t2993 VPWR.t120 76.3894
R3884 VPWR.t363 VPWR.t2892 76.3894
R3885 VPWR.t5252 VPWR.t1503 76.3894
R3886 VPWR.t6804 VPWR.t6954 76.2818
R3887 VPWR.t6819 VPWR.t6949 75.0899
R3888 VPWR.t110 VPWR.t3479 74.0746
R3889 VPWR.t3311 VPWR.t6552 74.0746
R3890 VPWR.t122 VPWR.t257 74.0746
R3891 VPWR.t6507 VPWR.t251 74.0746
R3892 VPWR.t5907 VPWR.t4510 74.0746
R3893 VPWR.t6129 VPWR.t2997 74.0746
R3894 VPWR.t606 VPWR.t1126 74.0746
R3895 VPWR.t968 VPWR.t1366 74.0746
R3896 VPWR.t4651 VPWR.t5131 74.0746
R3897 VPWR.t3573 VPWR.t4060 74.0746
R3898 VPWR.t2392 VPWR.t2578 74.0746
R3899 VPWR.t1729 VPWR.t2867 74.0746
R3900 VPWR.t3830 VPWR.t4688 73.898
R3901 VPWR.t1030 VPWR 72.9172
R3902 VPWR VPWR.t2337 72.9172
R3903 VPWR.t4851 VPWR.t900 72.9172
R3904 VPWR.t6639 VPWR.t352 72.9172
R3905 VPWR.t1324 VPWR.t5193 72.9172
R3906 VPWR VPWR.t2357 72.9172
R3907 VPWR.t1155 VPWR 72.9172
R3908 VPWR VPWR.t1667 72.9172
R3909 VPWR.t7047 VPWR.n2863 72.9172
R3910 VPWR.n2865 VPWR.t6463 72.9172
R3911 VPWR.t6585 VPWR.t4682 72.9172
R3912 VPWR.t7134 VPWR.n938 71.7598
R3913 VPWR.t4272 VPWR.t322 71.7598
R3914 VPWR.n846 VPWR.t3468 71.7598
R3915 VPWR.t5496 VPWR.t7096 71.7598
R3916 VPWR.t3598 VPWR.t5168 71.7598
R3917 VPWR.t3507 VPWR.t3809 71.7598
R3918 VPWR.t5397 VPWR.t6814 71.7598
R3919 VPWR.t1069 VPWR.t4966 71.7598
R3920 VPWR.t5740 VPWR.n729 71.7598
R3921 VPWR.n743 VPWR.t3841 71.7598
R3922 VPWR.t3970 VPWR.t222 71.7598
R3923 VPWR.t112 VPWR.t3492 71.7598
R3924 VPWR.t946 VPWR.n3256 71.7598
R3925 VPWR.t1790 VPWR.t2023 71.7598
R3926 VPWR.t4280 VPWR.n1172 71.7598
R3927 VPWR.n725 VPWR.t4437 71.7598
R3928 VPWR.t4205 VPWR.t5757 71.7598
R3929 VPWR.t5365 VPWR.t6587 71.7598
R3930 VPWR.t5191 VPWR.t207 71.7598
R3931 VPWR.t4981 VPWR.t6935 71.7598
R3932 VPWR.t6921 VPWR.t3361 71.7598
R3933 VPWR.t5511 VPWR.t127 71.7598
R3934 VPWR.t5183 VPWR.t6290 71.7598
R3935 VPWR.t5321 VPWR.t2140 71.7598
R3936 VPWR.t2916 VPWR.t5483 71.7598
R3937 VPWR.t4473 VPWR.t5618 71.7598
R3938 VPWR.t1944 VPWR.t3253 71.7598
R3939 VPWR.t5159 VPWR.n523 71.7598
R3940 VPWR.t2600 VPWR.n512 71.7598
R3941 VPWR.t1976 VPWR.t50 71.7598
R3942 VPWR.t308 VPWR.t7125 71.7598
R3943 VPWR.t1767 VPWR.t1063 71.7598
R3944 VPWR.t6415 VPWR.t2453 71.7598
R3945 VPWR.t3581 VPWR.t6404 71.5142
R3946 VPWR.t979 VPWR.t6846 71.5142
R3947 VPWR VPWR.t4247 70.6024
R3948 VPWR.t6624 VPWR.t3101 70.6024
R3949 VPWR.t6626 VPWR.t6995 70.6024
R3950 VPWR VPWR.t5342 70.6024
R3951 VPWR VPWR.t1019 70.6024
R3952 VPWR.t197 VPWR.t2597 70.6024
R3953 VPWR.t2044 VPWR.t4964 69.4449
R3954 VPWR.t6783 VPWR.t7000 69.4449
R3955 VPWR.t2033 VPWR.t6996 69.4449
R3956 VPWR.t6979 VPWR.t3003 69.4449
R3957 VPWR.t2323 VPWR.t4837 69.4449
R3958 VPWR.t2592 VPWR.t2394 69.4449
R3959 VPWR.t737 VPWR.t2125 69.4449
R3960 VPWR.t5393 VPWR.t1294 69.4449
R3961 VPWR VPWR.t5257 68.2875
R3962 VPWR.t6297 VPWR.t1621 67.1301
R3963 VPWR.n142 VPWR.t6676 67.1301
R3964 VPWR.t4980 VPWR.t6913 67.1301
R3965 VPWR.t3054 VPWR.t4999 67.1301
R3966 VPWR.t6744 VPWR.t3424 67.1301
R3967 VPWR.t6810 VPWR.t4686 66.7466
R3968 VPWR.t6709 VPWR.t4701 66.7466
R3969 VPWR VPWR.t173 65.9727
R3970 VPWR.t1383 VPWR.t7030 65.9727
R3971 VPWR VPWR.t6550 65.9727
R3972 VPWR.t285 VPWR 65.9727
R3973 VPWR VPWR.t6929 65.9727
R3974 VPWR VPWR.t6931 65.9727
R3975 VPWR VPWR.t6962 65.9727
R3976 VPWR VPWR.t5813 65.9727
R3977 VPWR.t6511 VPWR 65.5547
R3978 VPWR.t5138 VPWR 65.5547
R3979 VPWR.t6606 VPWR 65.5547
R3980 VPWR.t151 VPWR.t3533 64.8153
R3981 VPWR.t1692 VPWR.t6696 64.8153
R3982 VPWR.t7035 VPWR.t1056 64.8153
R3983 VPWR.t5985 VPWR.t4521 64.8153
R3984 VPWR.t5707 VPWR.t6739 64.8153
R3985 VPWR.t6607 VPWR.t1913 64.8153
R3986 VPWR.t4171 VPWR.t6649 64.8153
R3987 VPWR.t6661 VPWR.t584 64.8153
R3988 VPWR.t1330 VPWR.t6943 64.8153
R3989 VPWR.t468 VPWR.t4565 64.8153
R3990 VPWR.t4563 VPWR.t4462 64.8153
R3991 VPWR VPWR.t3138 63.6579
R3992 VPWR.t40 VPWR.n136 63.6579
R3993 VPWR.t3237 VPWR.t6398 63.6579
R3994 VPWR.t6546 VPWR 63.6579
R3995 VPWR VPWR.t1326 63.6579
R3996 VPWR.t121 VPWR.n187 63.6579
R3997 VPWR.t5164 VPWR.t6595 63.6579
R3998 VPWR.n755 VPWR.t4111 62.5005
R3999 VPWR.t6601 VPWR.t527 62.5005
R4000 VPWR.t6613 VPWR.t2352 61.979
R4001 VPWR.t6647 VPWR.t6531 61.979
R4002 VPWR.t5586 VPWR.t4237 61.3431
R4003 VPWR VPWR.t1597 61.3431
R4004 VPWR.t2739 VPWR.t4460 61.3431
R4005 VPWR VPWR.t2739 61.3431
R4006 VPWR.t6768 VPWR.t4514 60.1857
R4007 VPWR.t6492 VPWR.t6704 60.1857
R4008 VPWR.t5737 VPWR.t336 60.1857
R4009 VPWR.t4125 VPWR.t119 60.1857
R4010 VPWR.t6681 VPWR.t3045 60.1857
R4011 VPWR VPWR.n1397 59.0283
R4012 VPWR VPWR.t3158 59.0283
R4013 VPWR VPWR.t4435 59.0283
R4014 VPWR VPWR.n742 59.0283
R4015 VPWR.t2930 VPWR 59.0283
R4016 VPWR VPWR.n517 59.0283
R4017 VPWR.t1158 VPWR.n954 57.8709
R4018 VPWR.t2380 VPWR.t2559 57.8709
R4019 VPWR.n929 VPWR.t6788 57.8709
R4020 VPWR.t3138 VPWR.t5869 57.8709
R4021 VPWR.t6024 VPWR.t4381 57.8709
R4022 VPWR.t3095 VPWR.t5384 57.8709
R4023 VPWR.t1954 VPWR.n1278 57.8709
R4024 VPWR.t6383 VPWR.t2417 57.8709
R4025 VPWR.t7006 VPWR.t2795 57.8709
R4026 VPWR.n3262 VPWR.t4004 57.8709
R4027 VPWR.t6525 VPWR.t2091 57.8709
R4028 VPWR.t1993 VPWR.t5857 57.8709
R4029 VPWR.t6388 VPWR.n143 57.8709
R4030 VPWR.t3872 VPWR.t4708 57.8709
R4031 VPWR.t841 VPWR.t5185 57.8709
R4032 VPWR.t444 VPWR.t1316 57.8709
R4033 VPWR.n714 VPWR.t269 57.8709
R4034 VPWR.t154 VPWR.t4667 57.8709
R4035 VPWR.t3797 VPWR.t1859 57.8709
R4036 VPWR.t5601 VPWR.t6038 57.8709
R4037 VPWR.t5951 VPWR.t5311 57.8709
R4038 VPWR.t4576 VPWR.t6391 57.8709
R4039 VPWR.t4992 VPWR.t5437 57.8709
R4040 VPWR.t227 VPWR.t2505 57.8709
R4041 VPWR.n541 VPWR.t6886 57.8709
R4042 VPWR.t3114 VPWR.n458 57.8709
R4043 VPWR.n511 VPWR.t1727 57.8709
R4044 VPWR.t5087 VPWR.t3336 57.8709
R4045 VPWR.t5607 VPWR.t4095 57.8709
R4046 VPWR.n372 VPWR.t5784 57.8709
R4047 VPWR.t6503 VPWR.t6742 57.2115
R4048 VPWR VPWR.t4036 56.7135
R4049 VPWR.t6696 VPWR 56.7135
R4050 VPWR VPWR.t4818 56.7135
R4051 VPWR VPWR.t4421 56.7135
R4052 VPWR.t4560 VPWR.t6291 56.7135
R4053 VPWR.t5913 VPWR 56.7135
R4054 VPWR.t896 VPWR.t4236 56.7135
R4055 VPWR.t7008 VPWR.t2746 55.5561
R4056 VPWR.t4211 VPWR.t172 55.5561
R4057 VPWR.t173 VPWR.t6984 55.5561
R4058 VPWR.t3130 VPWR.t475 55.5561
R4059 VPWR.t2400 VPWR.t1270 55.5561
R4060 VPWR.t6550 VPWR.t3310 55.5561
R4061 VPWR.t6544 VPWR.t6981 55.5561
R4062 VPWR.t2121 VPWR.t4413 55.5561
R4063 VPWR.t2830 VPWR.t1493 55.5561
R4064 VPWR.t1637 VPWR.t752 55.5561
R4065 VPWR VPWR.t3182 54.3986
R4066 VPWR.t6379 VPWR 54.3986
R4067 VPWR.n3354 VPWR.t3411 53.2412
R4068 VPWR.t7099 VPWR.t3416 53.2412
R4069 VPWR.t6382 VPWR.t2231 53.2412
R4070 VPWR.t4148 VPWR.t3265 53.2412
R4071 VPWR.t354 VPWR.t6317 53.2412
R4072 VPWR.t4264 VPWR.t5423 53.2412
R4073 VPWR.t1563 VPWR.t162 53.2412
R4074 VPWR.t2255 VPWR.t2764 53.2412
R4075 VPWR.n2953 VPWR.t2898 53.2412
R4076 VPWR.t7112 VPWR.t5142 52.4439
R4077 VPWR.t4082 VPWR 52.0838
R4078 VPWR VPWR.t6624 52.0838
R4079 VPWR.t3579 VPWR.t6774 52.0838
R4080 VPWR.t4379 VPWR 52.0838
R4081 VPWR.t3878 VPWR 52.0838
R4082 VPWR VPWR.t2592 52.0838
R4083 VPWR VPWR.t737 52.0838
R4084 VPWR.t3060 VPWR 52.0838
R4085 VPWR VPWR.t4433 52.0838
R4086 VPWR.t1589 VPWR 52.0838
R4087 VPWR VPWR.t1048 52.0838
R4088 VPWR.t3972 VPWR 52.0838
R4089 VPWR VPWR.t5949 52.0838
R4090 VPWR.t4324 VPWR.t4695 52.0838
R4091 VPWR.t3299 VPWR.t4320 52.0838
R4092 VPWR.t3295 VPWR.t3297 52.0838
R4093 VPWR.t2824 VPWR 52.0838
R4094 VPWR VPWR.t6313 52.0838
R4095 VPWR.t1725 VPWR 52.0838
R4096 VPWR.t3338 VPWR 52.0838
R4097 VPWR.t3398 VPWR.t6611 51.252
R4098 VPWR.t4389 VPWR.t138 50.9264
R4099 VPWR.t6896 VPWR.t6490 50.9264
R4100 VPWR.t3290 VPWR.t147 50.9264
R4101 VPWR.t5777 VPWR.t4996 50.9264
R4102 VPWR.t3750 VPWR.t5896 50.9264
R4103 VPWR.t6787 VPWR.t4937 50.9264
R4104 VPWR.t1011 VPWR.t4049 50.9264
R4105 VPWR.t3255 VPWR.t5357 50.9264
R4106 VPWR.t3961 VPWR.t6554 50.9264
R4107 VPWR.t4908 VPWR.t6572 50.9264
R4108 VPWR.t3731 VPWR.t6919 50.9264
R4109 VPWR.t2035 VPWR.t6262 50.9264
R4110 VPWR.t213 VPWR.t1469 50.9264
R4111 VPWR.n394 VPWR.n393 50.0597
R4112 VPWR.t3805 VPWR 49.769
R4113 VPWR.t1333 VPWR 49.769
R4114 VPWR.t7129 VPWR 49.769
R4115 VPWR.t4702 VPWR 49.769
R4116 VPWR.t1522 VPWR 49.769
R4117 VPWR.t7073 VPWR 49.769
R4118 VPWR.t4419 VPWR 49.769
R4119 VPWR.t2188 VPWR 49.769
R4120 VPWR.t516 VPWR 49.769
R4121 VPWR.t5466 VPWR 49.769
R4122 VPWR.t1623 VPWR 49.769
R4123 VPWR.t1306 VPWR 49.769
R4124 VPWR.t3215 VPWR 49.769
R4125 VPWR.t3603 VPWR 49.769
R4126 VPWR.t4217 VPWR 49.769
R4127 VPWR.t3837 VPWR 49.769
R4128 VPWR.n100 VPWR 49.769
R4129 VPWR.n98 VPWR 49.769
R4130 VPWR VPWR.t3014 49.769
R4131 VPWR.n1400 VPWR.t3179 49.769
R4132 VPWR VPWR.t2325 49.769
R4133 VPWR VPWR.t1698 49.769
R4134 VPWR VPWR.n846 49.769
R4135 VPWR.t5168 VPWR 49.769
R4136 VPWR.t900 VPWR 49.769
R4137 VPWR.t2507 VPWR.t1825 49.769
R4138 VPWR.t352 VPWR 49.769
R4139 VPWR.t3809 VPWR 49.769
R4140 VPWR.t5442 VPWR.t5817 49.769
R4141 VPWR.t5193 VPWR 49.769
R4142 VPWR VPWR.t342 49.769
R4143 VPWR VPWR.t5216 49.769
R4144 VPWR.t6094 VPWR 49.769
R4145 VPWR VPWR.t705 49.769
R4146 VPWR.t4966 VPWR 49.769
R4147 VPWR VPWR.t4192 49.769
R4148 VPWR.t4043 VPWR 49.769
R4149 VPWR VPWR.n743 49.769
R4150 VPWR.t3492 VPWR 49.769
R4151 VPWR VPWR.t1995 49.769
R4152 VPWR VPWR.t2614 49.769
R4153 VPWR.n1172 VPWR 49.769
R4154 VPWR VPWR.n725 49.769
R4155 VPWR VPWR.t582 49.769
R4156 VPWR.t4441 VPWR 49.769
R4157 VPWR.t5757 VPWR 49.769
R4158 VPWR.t6268 VPWR 49.769
R4159 VPWR.t448 VPWR 49.769
R4160 VPWR VPWR.t3996 49.769
R4161 VPWR VPWR.t5365 49.769
R4162 VPWR VPWR.t1453 49.769
R4163 VPWR VPWR.t760 49.769
R4164 VPWR.t2176 VPWR 49.769
R4165 VPWR VPWR.t1717 49.769
R4166 VPWR VPWR.t5965 49.769
R4167 VPWR VPWR.t2070 49.769
R4168 VPWR.t2634 VPWR 49.769
R4169 VPWR.t6453 VPWR 49.769
R4170 VPWR.t4956 VPWR 49.769
R4171 VPWR VPWR.t6264 49.769
R4172 VPWR VPWR.t562 49.769
R4173 VPWR.t5162 VPWR 49.769
R4174 VPWR.t4310 VPWR 49.769
R4175 VPWR.t1071 VPWR 49.769
R4176 VPWR.t5821 VPWR 49.769
R4177 VPWR.t5978 VPWR 49.769
R4178 VPWR VPWR.t1549 49.769
R4179 VPWR.t3317 VPWR 49.769
R4180 VPWR.t4446 VPWR 49.769
R4181 VPWR VPWR.t5172 49.769
R4182 VPWR VPWR.t4512 49.769
R4183 VPWR VPWR.t4914 49.769
R4184 VPWR VPWR.t3550 49.769
R4185 VPWR VPWR.t4856 49.769
R4186 VPWR VPWR.t2797 49.769
R4187 VPWR.t5994 VPWR 49.769
R4188 VPWR VPWR.t3782 49.769
R4189 VPWR VPWR.n2324 49.769
R4190 VPWR VPWR.t985 49.769
R4191 VPWR VPWR.t5957 49.769
R4192 VPWR VPWR.t4274 49.769
R4193 VPWR VPWR.t6435 49.769
R4194 VPWR VPWR.t1855 49.769
R4195 VPWR.t5293 VPWR 49.769
R4196 VPWR.t2140 VPWR 49.769
R4197 VPWR.t5246 VPWR 49.769
R4198 VPWR VPWR.t7083 49.769
R4199 VPWR VPWR.t5959 49.769
R4200 VPWR VPWR.t5654 49.769
R4201 VPWR.t5483 VPWR 49.769
R4202 VPWR VPWR.n203 49.769
R4203 VPWR VPWR.n205 49.769
R4204 VPWR VPWR.t2876 49.769
R4205 VPWR VPWR.t4825 49.769
R4206 VPWR VPWR.t2674 49.769
R4207 VPWR.t5618 VPWR 49.769
R4208 VPWR.n512 VPWR 49.769
R4209 VPWR.t6580 VPWR.t6346 49.769
R4210 VPWR.t3198 VPWR 49.769
R4211 VPWR VPWR.t2253 49.769
R4212 VPWR VPWR.n385 49.769
R4213 VPWR VPWR.n370 49.769
R4214 VPWR.t7125 VPWR 49.769
R4215 VPWR.t1063 VPWR 49.769
R4216 VPWR VPWR.t5348 49.769
R4217 VPWR VPWR.n373 49.769
R4218 VPWR VPWR.t5582 49.769
R4219 VPWR VPWR.t3403 49.769
R4220 VPWR VPWR.n3707 49.769
R4221 VPWR.n63 VPWR 49.769
R4222 VPWR VPWR.n86 49.769
R4223 VPWR.t3839 VPWR.t776 48.6116
R4224 VPWR.t2396 VPWR.t1861 48.6116
R4225 VPWR.t2123 VPWR.t4159 48.6116
R4226 VPWR.t4988 VPWR.t5046 48.6116
R4227 VPWR.t2196 VPWR.t6609 48.6116
R4228 VPWR.n964 VPWR.t2734 48.4402
R4229 VPWR.n963 VPWR 47.9054
R4230 VPWR.n952 VPWR 47.9054
R4231 VPWR.n1402 VPWR 47.9054
R4232 VPWR.n826 VPWR 47.9054
R4233 VPWR.n3260 VPWR 47.9054
R4234 VPWR.n149 VPWR 47.9054
R4235 VPWR.t3479 VPWR 47.4542
R4236 VPWR.t6716 VPWR 47.4542
R4237 VPWR.t5140 VPWR.t6623 46.9764
R4238 VPWR.t6674 VPWR.t6361 46.2968
R4239 VPWR.t2085 VPWR.t3474 46.2968
R4240 VPWR VPWR.t6468 45.1394
R4241 VPWR.t145 VPWR 45.1394
R4242 VPWR.t4075 VPWR 45.1394
R4243 VPWR VPWR.t2657 45.1394
R4244 VPWR.t3489 VPWR 45.1394
R4245 VPWR.t6758 VPWR 45.1394
R4246 VPWR.t5923 VPWR 45.1394
R4247 VPWR.t6998 VPWR 45.1394
R4248 VPWR.t5475 VPWR 45.1394
R4249 VPWR VPWR.t645 45.1394
R4250 VPWR.t2447 VPWR 45.1394
R4251 VPWR.t789 VPWR.t1169 45.1394
R4252 VPWR.t6087 VPWR.t790 45.1394
R4253 VPWR.t5212 VPWR.t7017 45.1394
R4254 VPWR VPWR.t5391 45.1394
R4255 VPWR.t184 VPWR 45.1394
R4256 VPWR.t5446 VPWR 45.1394
R4257 VPWR.n945 VPWR 44.4063
R4258 VPWR.n933 VPWR 44.4063
R4259 VPWR.n1404 VPWR 44.4063
R4260 VPWR.n844 VPWR 44.4063
R4261 VPWR.n3267 VPWR 44.4063
R4262 VPWR.n741 VPWR 44.4063
R4263 VPWR.t1526 VPWR.t1528 43.982
R4264 VPWR.t1524 VPWR.t1530 43.982
R4265 VPWR.n1392 VPWR.t6733 43.982
R4266 VPWR.n115 VPWR.t2557 43.982
R4267 VPWR.t1651 VPWR.t3748 43.982
R4268 VPWR.t1339 VPWR.n3269 43.982
R4269 VPWR.t4071 VPWR.n151 43.982
R4270 VPWR.t4157 VPWR.t2729 43.982
R4271 VPWR.t5425 VPWR.t3542 43.982
R4272 VPWR.t2064 VPWR.t1455 43.982
R4273 VPWR.t6002 VPWR.t5127 43.982
R4274 VPWR.t6004 VPWR.t5125 43.982
R4275 VPWR.t4608 VPWR.t4144 43.982
R4276 VPWR.t4606 VPWR.t4142 43.982
R4277 VPWR.t510 VPWR.t6162 43.982
R4278 VPWR.t508 VPWR.t6164 43.982
R4279 VPWR.t5189 VPWR.t506 43.982
R4280 VPWR.t5187 VPWR.t504 43.982
R4281 VPWR VPWR.t3409 42.8246
R4282 VPWR.t2637 VPWR 42.8246
R4283 VPWR.t211 VPWR.t5632 42.8246
R4284 VPWR.t2537 VPWR.t3623 42.8246
R4285 VPWR.t5594 VPWR.t3569 42.8246
R4286 VPWR.t2900 VPWR 42.8246
R4287 VPWR VPWR.t171 42.5063
R4288 VPWR.t4960 VPWR.t5925 41.6672
R4289 VPWR.t6861 VPWR.t5487 41.6672
R4290 VPWR.t4222 VPWR.t15 41.6672
R4291 VPWR.t6671 VPWR.t4006 41.6672
R4292 VPWR.t3373 VPWR.t2650 41.6672
R4293 VPWR.t2957 VPWR.t4107 41.6672
R4294 VPWR.t3482 VPWR.t3476 41.6672
R4295 VPWR.t6540 VPWR.t479 41.6672
R4296 VPWR.t3344 VPWR.t4231 41.6672
R4297 VPWR.t6604 VPWR.t6107 41.6672
R4298 VPWR.t6917 VPWR.t5628 41.6672
R4299 VPWR VPWR.t2733 40.5098
R4300 VPWR.t2573 VPWR.t7065 40.5098
R4301 VPWR.t4282 VPWR.t3150 40.5098
R4302 VPWR.t6400 VPWR 40.5098
R4303 VPWR.t2346 VPWR.t41 40.5068
R4304 VPWR.t887 VPWR.t1929 39.3524
R4305 VPWR VPWR.t6081 39.3524
R4306 VPWR.n1397 VPWR 39.3524
R4307 VPWR.n1405 VPWR 39.3524
R4308 VPWR.t4085 VPWR.t881 39.3524
R4309 VPWR VPWR.n150 39.3524
R4310 VPWR.n624 VPWR.t3915 39.3524
R4311 VPWR.n377 VPWR.t4328 38.4207
R4312 VPWR VPWR.t5009 38.1949
R4313 VPWR.t3267 VPWR.t6653 38.1949
R4314 VPWR.t5596 VPWR.t3570 38.1949
R4315 VPWR.t3305 VPWR.t1473 38.1949
R4316 VPWR.t4796 VPWR.t6711 38.1949
R4317 VPWR VPWR.t2134 38.1949
R4318 VPWR VPWR.t4014 38.1949
R4319 VPWR.t6367 VPWR.t1617 37.0375
R4320 VPWR.t2160 VPWR.t5479 37.0375
R4321 VPWR.t2161 VPWR.t804 37.0375
R4322 VPWR.t6505 VPWR.t6618 37.0375
R4323 VPWR.t4155 VPWR.t1583 37.0375
R4324 VPWR.t6420 VPWR.t1796 37.0375
R4325 VPWR.t960 VPWR.t5146 37.0375
R4326 VPWR.t6422 VPWR.t6583 37.0375
R4327 VPWR.t4792 VPWR.t3932 37.0375
R4328 VPWR.t5049 VPWR.t3180 35.8801
R4329 VPWR.t4450 VPWR.t7059 35.8801
R4330 VPWR.t7043 VPWR.t835 35.8801
R4331 VPWR VPWR.t2285 35.8801
R4332 VPWR.t4326 VPWR 35.8801
R4333 VPWR.n1035 VPWR.t6879 34.7227
R4334 VPWR.t6645 VPWR.t4302 34.7227
R4335 VPWR.t3011 VPWR.t6643 34.7227
R4336 VPWR.t5763 VPWR.t6665 34.7227
R4337 VPWR.t4986 VPWR.t6958 34.7227
R4338 VPWR.t6892 VPWR.t4849 34.7227
R4339 VPWR.t1107 VPWR 33.5653
R4340 VPWR VPWR.t5738 33.5653
R4341 VPWR VPWR.t7012 33.5653
R4342 VPWR.t6568 VPWR 33.5653
R4343 VPWR.t6558 VPWR 33.5653
R4344 VPWR.t6556 VPWR 33.5653
R4345 VPWR VPWR.t295 33.5653
R4346 VPWR.t275 VPWR 33.5653
R4347 VPWR.t3350 VPWR 33.5653
R4348 VPWR.t4791 VPWR.t1472 33.5653
R4349 VPWR.t6927 VPWR 33.5653
R4350 VPWR.t5051 VPWR.t433 32.4079
R4351 VPWR.t5563 VPWR.t5571 32.4079
R4352 VPWR.t6955 VPWR.t6428 32.4079
R4353 VPWR VPWR.t6852 32.1817
R4354 VPWR.t6538 VPWR 32.1817
R4355 VPWR VPWR.t3577 31.2505
R4356 VPWR VPWR.t5005 31.2505
R4357 VPWR.t4797 VPWR 31.2505
R4358 VPWR.t5155 VPWR.t6731 31.2505
R4359 VPWR.n1403 VPWR.t1054 31.05
R4360 VPWR.t3829 VPWR.t4680 30.9898
R4361 VPWR.t4399 VPWR.n947 30.0931
R4362 VPWR VPWR.t523 30.0931
R4363 VPWR.t5622 VPWR.t2880 30.0931
R4364 VPWR.t5624 VPWR.t2183 30.0931
R4365 VPWR.t1101 VPWR.t2277 30.0931
R4366 VPWR.t4278 VPWR.t3586 30.0931
R4367 VPWR.t5410 VPWR.t1865 30.0931
R4368 VPWR.t6166 VPWR.t537 30.0931
R4369 VPWR.t539 VPWR.t5613 30.0931
R4370 VPWR.t5692 VPWR.t5525 30.0931
R4371 VPWR.t4721 VPWR.t735 30.0931
R4372 VPWR.t5337 VPWR.t3988 30.0931
R4373 VPWR.n2951 VPWR.t2001 30.0931
R4374 VPWR.t2861 VPWR.t5114 30.0931
R4375 VPWR.t2857 VPWR.t5492 30.0931
R4376 VPWR.t6535 VPWR.n845 29.5926
R4377 VPWR VPWR.t1354 28.9357
R4378 VPWR VPWR.t2640 28.9357
R4379 VPWR VPWR.t3484 28.9357
R4380 VPWR.t6888 VPWR.t35 28.9357
R4381 VPWR.t3716 VPWR 28.9357
R4382 VPWR.t3022 VPWR.t6239 28.606
R4383 VPWR.t4037 VPWR.t4879 27.7783
R4384 VPWR.t670 VPWR.t6780 27.7783
R4385 VPWR.t6402 VPWR.t2555 27.7783
R4386 VPWR.t4334 VPWR.t4431 27.7783
R4387 VPWR.t594 VPWR.t4831 27.7783
R4388 VPWR.t6993 VPWR.t6292 27.7783
R4389 VPWR VPWR.t4821 27.7783
R4390 VPWR.n1175 VPWR.t1688 27.7783
R4391 VPWR.t3070 VPWR.t5323 27.7783
R4392 VPWR.t1905 VPWR.t2462 27.7783
R4393 VPWR.t3291 VPWR 26.6209
R4394 VPWR.t6946 VPWR 26.6209
R4395 VPWR.t1520 VPWR 26.6209
R4396 VPWR.t1156 VPWR 26.6209
R4397 VPWR.t6371 VPWR 26.6209
R4398 VPWR.t6406 VPWR 26.6209
R4399 VPWR.t588 VPWR 26.6209
R4400 VPWR.t5823 VPWR.t6890 26.6209
R4401 VPWR.t6598 VPWR 26.6209
R4402 VPWR.n853 VPWR.t6575 25.4635
R4403 VPWR.t3646 VPWR.t1083 25.4635
R4404 VPWR.t0 VPWR.t849 25.4635
R4405 VPWR.t6582 VPWR.t6881 25.4635
R4406 VPWR VPWR.t5022 24.3061
R4407 VPWR.t413 VPWR.t5016 24.3061
R4408 VPWR VPWR.t6048 24.3061
R4409 VPWR VPWR.t403 24.3061
R4410 VPWR.t6482 VPWR.t1777 23.1486
R4411 VPWR VPWR.t5210 23.1486
R4412 VPWR.t6750 VPWR.t2768 23.1486
R4413 VPWR VPWR.t1881 23.1486
R4414 VPWR.t5929 VPWR.t6515 23.1486
R4415 VPWR.t6522 VPWR.t6519 23.1486
R4416 VPWR.t4091 VPWR.t6854 23.1486
R4417 VPWR.t2029 VPWR.t793 23.1486
R4418 VPWR.t6792 VPWR.t797 23.1486
R4419 VPWR.t788 VPWR.t2238 23.1486
R4420 VPWR.t2508 VPWR.t3835 23.1486
R4421 VPWR.t4111 VPWR.t142 23.1486
R4422 VPWR.t4561 VPWR 23.1486
R4423 VPWR.t1264 VPWR.t247 23.1486
R4424 VPWR.t6800 VPWR.t271 23.1486
R4425 VPWR.t7032 VPWR.t6667 23.1486
R4426 VPWR.t4800 VPWR.t131 23.1486
R4427 VPWR.t5153 VPWR.t4795 23.1486
R4428 VPWR.t4132 VPWR.t3610 23.1486
R4429 VPWR.t3791 VPWR 21.9912
R4430 VPWR VPWR.t6635 21.9912
R4431 VPWR VPWR.t6760 21.9912
R4432 VPWR.t6042 VPWR 21.9912
R4433 VPWR.t3635 VPWR 21.9912
R4434 VPWR VPWR.t4089 21.9912
R4435 VPWR VPWR.t4042 21.9912
R4436 VPWR.t6869 VPWR 21.9912
R4437 VPWR.t3564 VPWR 21.9912
R4438 VPWR VPWR.t1956 21.9912
R4439 VPWR.t3505 VPWR 21.9912
R4440 VPWR.t1490 VPWR 21.9912
R4441 VPWR VPWR.t2878 21.9912
R4442 VPWR.t5626 VPWR 21.9912
R4443 VPWR.t4429 VPWR 21.9912
R4444 VPWR VPWR.t981 21.9912
R4445 VPWR.t2781 VPWR 21.9912
R4446 VPWR VPWR.t1867 21.9912
R4447 VPWR.t1272 VPWR 21.9912
R4448 VPWR VPWR.t972 21.9912
R4449 VPWR.t6883 VPWR.n628 21.9912
R4450 VPWR.t253 VPWR 21.9912
R4451 VPWR VPWR.t1581 21.9912
R4452 VPWR VPWR.t1684 21.9912
R4453 VPWR VPWR.t535 21.9912
R4454 VPWR.t541 VPWR 21.9912
R4455 VPWR VPWR.t5527 21.9912
R4456 VPWR.t4411 VPWR 21.9912
R4457 VPWR VPWR.t729 21.9912
R4458 VPWR.t1491 VPWR 21.9912
R4459 VPWR VPWR.t1639 21.9912
R4460 VPWR VPWR.t733 21.9912
R4461 VPWR.t5339 VPWR 21.9912
R4462 VPWR.t1749 VPWR 21.9912
R4463 VPWR.t3462 VPWR 21.9912
R4464 VPWR VPWR.t4842 21.9912
R4465 VPWR.t2500 VPWR 21.9912
R4466 VPWR VPWR.t5112 21.9912
R4467 VPWR.t2859 VPWR 21.9912
R4468 VPWR.n1441 VPWR.t2336 21.6375
R4469 VPWR.n1426 VPWR.t2159 21.6375
R4470 VPWR.n1001 VPWR.t1032 21.6375
R4471 VPWR.n985 VPWR.t4038 21.6375
R4472 VPWR.n3376 VPWR.t6098 21.6375
R4473 VPWR.n997 VPWR.t1930 21.6375
R4474 VPWR.n1010 VPWR.t3292 21.6375
R4475 VPWR.n1611 VPWR.t669 21.6375
R4476 VPWR.n1415 VPWR.t806 21.6375
R4477 VPWR.n906 VPWR.t1521 21.6375
R4478 VPWR.n3366 VPWR.t2639 21.6375
R4479 VPWR.n3352 VPWR.t3412 21.6375
R4480 VPWR.n892 VPWR.t5486 21.6375
R4481 VPWR.n789 VPWR.t6007 21.6375
R4482 VPWR.n774 VPWR.t3266 21.6375
R4483 VPWR.n3308 VPWR.t1157 21.6375
R4484 VPWR.n3279 VPWR.t5616 21.6375
R4485 VPWR.n3297 VPWR.t4817 21.6375
R4486 VPWR.n800 VPWR.t6298 21.6375
R4487 VPWR.n1687 VPWR.t3284 21.6375
R4488 VPWR.n3214 VPWR.t5912 21.6375
R4489 VPWR.n3197 VPWR.t6293 21.6375
R4490 VPWR.n3183 VPWR.t4423 21.6375
R4491 VPWR.n3206 VPWR.t6318 21.6375
R4492 VPWR.n1790 VPWR.t1666 21.6375
R4493 VPWR.n663 VPWR.t1912 21.6375
R4494 VPWR.n1112 VPWR.t3984 21.6375
R4495 VPWR.n1942 VPWR.t5424 21.6375
R4496 VPWR.n2856 VPWR.t3897 21.6375
R4497 VPWR.n2894 VPWR.t1329 21.6375
R4498 VPWR.n2901 VPWR.t1848 21.6375
R4499 VPWR.n184 VPWR.t5976 21.6375
R4500 VPWR.n2796 VPWR.t5013 21.6375
R4501 VPWR.n1871 VPWR.t3943 21.6375
R4502 VPWR.n3029 VPWR.t1468 21.6375
R4503 VPWR.n409 VPWR.t2078 21.6375
R4504 VPWR.n3017 VPWR.t2899 21.6375
R4505 VPWR.n408 VPWR.t2599 21.6375
R4506 VPWR.n433 VPWR.t438 21.6375
R4507 VPWR.t525 VPWR.t6031 20.8338
R4508 VPWR.t3235 VPWR.t786 20.8338
R4509 VPWR.n378 VPWR.t942 20.8338
R4510 VPWR.n1091 VPWR.t2107 19.7193
R4511 VPWR.n3357 VPWR.t3892 19.7133
R4512 VPWR.n155 VPWR.t2801 19.7133
R4513 VPWR VPWR.t2048 19.6764
R4514 VPWR VPWR.t6303 19.6764
R4515 VPWR.t2259 VPWR 19.6764
R4516 VPWR VPWR.t4203 19.6764
R4517 VPWR VPWR.t5672 19.6764
R4518 VPWR.t3273 VPWR.t4135 19.6764
R4519 VPWR.n394 VPWR.t1113 19.6764
R4520 VPWR.n1397 VPWR.t4911 19.2697
R4521 VPWR.n3273 VPWR.t1023 19.2697
R4522 VPWR.n755 VPWR.t5514 19.2697
R4523 VPWR.n760 VPWR.t2940 19.2697
R4524 VPWR.n141 VPWR.t6073 19.2697
R4525 VPWR.n634 VPWR.t1033 19.2697
R4526 VPWR.n1938 VPWR.t2673 19.2697
R4527 VPWR.n2880 VPWR.t638 19.2697
R4528 VPWR.n2748 VPWR.t2636 19.2697
R4529 VPWR.n175 VPWR.t5470 19.2697
R4530 VPWR.n2952 VPWR.t2708 19.2697
R4531 VPWR.n928 VPWR.t3561 19.268
R4532 VPWR.n114 VPWR.t6215 19.268
R4533 VPWR.n749 VPWR.t3630 19.268
R4534 VPWR.n142 VPWR.t3129 19.268
R4535 VPWR.n1782 VPWR.t5641 19.268
R4536 VPWR.n2879 VPWR.t6310 19.268
R4537 VPWR.n377 VPWR.t5977 19.268
R4538 VPWR.t6513 VPWR.t6574 19.0708
R4539 VPWR.t6509 VPWR.t6625 19.0708
R4540 VPWR.n2865 VPWR.n2864 18.5307
R4541 VPWR.n2863 VPWR.n2862 18.5289
R4542 VPWR.t140 VPWR.t6901 18.519
R4543 VPWR.t149 VPWR.t3535 18.519
R4544 VPWR.t3229 VPWR.t6518 18.519
R4545 VPWR.t6676 VPWR.t6386 18.519
R4546 VPWR.t6663 VPWR.t3870 18.519
R4547 VPWR.t5488 VPWR.t6802 18.519
R4548 VPWR.t4173 VPWR.t3896 18.519
R4549 VPWR.t5975 VPWR.t586 18.519
R4550 VPWR.t6960 VPWR.t6426 18.519
R4551 VPWR.t5120 VPWR 18.519
R4552 VPWR.n945 VPWR.t1423 18.2762
R4553 VPWR.n933 VPWR.t851 18.2762
R4554 VPWR.n1404 VPWR.t5084 18.2762
R4555 VPWR.n844 VPWR.t4039 18.2762
R4556 VPWR.n3267 VPWR.t866 18.2762
R4557 VPWR.n741 VPWR.t5256 18.2762
R4558 VPWR.n1092 VPWR.n1091 18.2373
R4559 VPWR.n3358 VPWR.n3357 18.2334
R4560 VPWR.n156 VPWR.n155 18.2334
R4561 VPWR.n963 VPWR.t1177 18.1997
R4562 VPWR.n952 VPWR.t4296 18.1997
R4563 VPWR.n1402 VPWR.t3157 18.1997
R4564 VPWR.n826 VPWR.t299 18.1997
R4565 VPWR.n3260 VPWR.t2301 18.1997
R4566 VPWR.n149 VPWR.t2574 18.1997
R4567 VPWR.t2359 VPWR.t6533 17.6165
R4568 VPWR.t1948 VPWR.t5670 17.3616
R4569 VPWR.t1946 VPWR.t2735 17.3616
R4570 VPWR VPWR.t7062 17.3616
R4571 VPWR.t203 VPWR.t6735 17.3616
R4572 VPWR VPWR.t2560 17.3616
R4573 VPWR.t1337 VPWR 17.3616
R4574 VPWR.t5590 VPWR.t6589 17.3616
R4575 VPWR VPWR.t94 16.2042
R4576 VPWR.n1038 VPWR.t1105 16.2042
R4577 VPWR.t6694 VPWR.n912 16.2042
R4578 VPWR VPWR.t6340 16.2042
R4579 VPWR.n1778 VPWR.t279 16.2042
R4580 VPWR VPWR.t156 16.2042
R4581 VPWR.t233 VPWR.t2504 16.2042
R4582 VPWR VPWR.t1258 15.0468
R4583 VPWR VPWR.t6478 15.0468
R4584 VPWR.t5268 VPWR 15.0468
R4585 VPWR.t6026 VPWR.t2435 15.0468
R4586 VPWR.t3637 VPWR 15.0468
R4587 VPWR.t3679 VPWR 15.0468
R4588 VPWR.t2772 VPWR.t114 15.0468
R4589 VPWR VPWR.t6982 15.0468
R4590 VPWR.t6766 VPWR 15.0468
R4591 VPWR VPWR.t6651 15.0468
R4592 VPWR.t2543 VPWR.t3622 15.0468
R4593 VPWR.t2539 VPWR.t2457 15.0468
R4594 VPWR.t907 VPWR 15.0468
R4595 VPWR.t895 VPWR.t6713 15.0468
R4596 VPWR.t938 VPWR 15.0468
R4597 VPWR VPWR.t6952 15.0468
R4598 VPWR VPWR.t3771 15.0468
R4599 VPWR.t4464 VPWR.t4465 15.0468
R4600 VPWR VPWR.t6641 15.0468
R4601 VPWR.t1927 VPWR.t1928 14.0933
R4602 VPWR.t160 VPWR 13.8894
R4603 VPWR.t7041 VPWR.t6700 13.8894
R4604 VPWR.t5807 VPWR.t6718 13.8894
R4605 VPWR.t6612 VPWR 13.8894
R4606 VPWR.t7020 VPWR.t1591 13.8894
R4607 VPWR.t116 VPWR.t774 13.8894
R4608 VPWR.t6296 VPWR.t6008 13.8894
R4609 VPWR.t221 VPWR 13.8894
R4610 VPWR.t208 VPWR.t6863 13.8894
R4611 VPWR.t6741 VPWR.t2990 13.8894
R4612 VPWR.t6387 VPWR 13.8894
R4613 VPWR.t273 VPWR.t6840 13.8894
R4614 VPWR.t259 VPWR.t6832 13.8894
R4615 VPWR.t263 VPWR.t6836 13.8894
R4616 VPWR.t261 VPWR.t6834 13.8894
R4617 VPWR.t255 VPWR.t6838 13.8894
R4618 VPWR.t249 VPWR.t6844 13.8894
R4619 VPWR.t243 VPWR.t6842 13.8894
R4620 VPWR.t687 VPWR.t3223 13.8894
R4621 VPWR.t6825 VPWR.t6602 13.8894
R4622 VPWR.t3974 VPWR.t1585 13.8894
R4623 VPWR.t6826 VPWR.t210 13.8894
R4624 VPWR.t93 VPWR 13.8894
R4625 VPWR.t6596 VPWR.t3422 13.8894
R4626 VPWR.t214 VPWR.t6821 13.8894
R4627 VPWR.t2502 VPWR.t4840 13.8894
R4628 VPWR.n2864 VPWR.t3898 13.358
R4629 VPWR.n2862 VPWR.t5974 13.3555
R4630 VPWR.n618 VPWR.t4982 12.8338
R4631 VPWR.n530 VPWR.t5439 12.8338
R4632 VPWR.t3148 VPWR.t6638 12.732
R4633 VPWR.t4309 VPWR 12.732
R4634 VPWR.t6462 VPWR.t7047 12.732
R4635 VPWR.t6463 VPWR.t7046 12.732
R4636 VPWR.n517 VPWR.n516 12.2511
R4637 VPWR.n1025 VPWR.t4138 11.8234
R4638 VPWR.n1031 VPWR.t2922 11.8234
R4639 VPWR.n1066 VPWR.t341 11.8234
R4640 VPWR.n1056 VPWR.t1380 11.8234
R4641 VPWR.n621 VPWR.t3732 11.8234
R4642 VPWR.n528 VPWR.t6240 11.8234
R4643 VPWR.t5116 VPWR.t2953 11.7445
R4644 VPWR.n1447 VPWR.t6737 11.662
R4645 VPWR.n965 VPWR.t1356 11.5746
R4646 VPWR.t205 VPWR.t6947 11.5746
R4647 VPWR.t1886 VPWR.n3355 11.5746
R4648 VPWR.t4835 VPWR.t334 11.5746
R4649 VPWR.t5089 VPWR.t4330 11.5746
R4650 VPWR.t553 VPWR.t2932 11.5746
R4651 VPWR.t1833 VPWR.n2874 11.5746
R4652 VPWR.n176 VPWR.t2058 11.5746
R4653 VPWR.n393 VPWR.t2077 11.1222
R4654 VPWR VPWR.t4804 10.4172
R4655 VPWR.n1099 VPWR.t1269 10.4088
R4656 VPWR.n587 VPWR.t6717 10.4088
R4657 VPWR.n1666 VPWR.t6730 10.3175
R4658 VPWR.n3253 VPWR.t6407 10.3175
R4659 VPWR.n3231 VPWR.t3472 10.238
R4660 VPWR.t5848 VPWR.t6795 9.39569
R4661 VPWR.n1371 VPWR.t3834 9.29022
R4662 VPWR.n130 VPWR.t481 9.29022
R4663 VPWR.n126 VPWR.t6987 9.29022
R4664 VPWR.n2868 VPWR.t6393 9.29022
R4665 VPWR.n2869 VPWR.t5564 9.29022
R4666 VPWR.n543 VPWR.t6380 9.29022
R4667 VPWR.n1406 VPWR.n1403 9.25976
R4668 VPWR.n114 VPWR 9.25976
R4669 VPWR VPWR.n141 9.25976
R4670 VPWR.t6375 VPWR.t5674 9.25976
R4671 VPWR.n634 VPWR.n632 9.25976
R4672 VPWR.t3724 VPWR.t3395 9.25976
R4673 VPWR.t5043 VPWR.t6392 9.25976
R4674 VPWR.n175 VPWR 9.25976
R4675 VPWR VPWR.n2952 9.25976
R4676 VPWR.t2704 VPWR.t2575 9.25976
R4677 VPWR.t302 VPWR.t439 9.25976
R4678 VPWR.t1918 VPWR.t5552 9.25976
R4679 VPWR.t3124 VPWR.n1405 9.14042
R4680 VPWR.n760 VPWR.t7117 9.13976
R4681 VPWR.n150 VPWR.t371 9.13976
R4682 VPWR.n1938 VPWR.t2993 9.13976
R4683 VPWR VPWR.t4315 8.64224
R4684 VPWR VPWR.t6630 8.64224
R4685 VPWR VPWR.t47 8.64224
R4686 VPWR VPWR.t6994 8.64224
R4687 VPWR VPWR.t5570 8.64224
R4688 VPWR VPWR.t6412 8.34377
R4689 VPWR.n987 VPWR.t2554 8.32188
R4690 VPWR.n3330 VPWR.t4090 8.32188
R4691 VPWR.n1679 VPWR.t3309 8.32188
R4692 VPWR.n1802 VPWR.t5119 8.32188
R4693 VPWR.n1103 VPWR.t190 8.32188
R4694 VPWR.n642 VPWR.t4206 8.32188
R4695 VPWR.n668 VPWR.t6608 8.32188
R4696 VPWR.n551 VPWR.t6592 8.32188
R4697 VPWR.n559 VPWR.t3352 8.32188
R4698 VPWR.n2940 VPWR.t6882 8.32188
R4699 VPWR.n1452 VPWR.t6734 8.29207
R4700 VPWR.n692 VPWR.t6603 8.29207
R4701 VPWR.n560 VPWR.t6584 8.29207
R4702 VPWR.n420 VPWR.t5002 8.29207
R4703 VPWR.t6680 VPWR 8.10235
R4704 VPWR VPWR.t1212 8.10235
R4705 VPWR VPWR.t1741 8.10235
R4706 VPWR VPWR.t6343 8.10235
R4707 VPWR VPWR.t4870 8.10235
R4708 VPWR.t5935 VPWR 8.10235
R4709 VPWR VPWR.t2237 8.10235
R4710 VPWR VPWR.t6793 8.10235
R4711 VPWR.t5895 VPWR 8.10235
R4712 VPWR.t2655 VPWR 8.10235
R4713 VPWR.t6278 VPWR 8.10235
R4714 VPWR.t102 VPWR 8.10235
R4715 VPWR VPWR.t3582 8.10235
R4716 VPWR VPWR.t5722 8.10235
R4717 VPWR.t6338 VPWR 8.10235
R4718 VPWR.t3636 VPWR.t7005 8.10235
R4719 VPWR.t2485 VPWR 8.10235
R4720 VPWR.t6061 VPWR 8.10235
R4721 VPWR VPWR.t2223 8.10235
R4722 VPWR.t6732 VPWR 8.10235
R4723 VPWR.t143 VPWR 8.10235
R4724 VPWR VPWR.t3470 8.10235
R4725 VPWR VPWR.t474 8.10235
R4726 VPWR.t2455 VPWR.t5592 8.10235
R4727 VPWR VPWR.t5118 8.10235
R4728 VPWR VPWR.t1686 8.10235
R4729 VPWR.t6830 VPWR 8.10235
R4730 VPWR.t4472 VPWR 8.10235
R4731 VPWR.t3914 VPWR 8.10235
R4732 VPWR.t3913 VPWR 8.10235
R4733 VPWR VPWR.t1292 8.10235
R4734 VPWR VPWR.t189 8.10235
R4735 VPWR.t1682 VPWR 8.10235
R4736 VPWR.t5885 VPWR 8.10235
R4737 VPWR VPWR.t6254 8.10235
R4738 VPWR.t2119 VPWR 8.10235
R4739 VPWR VPWR.t2890 8.10235
R4740 VPWR VPWR.t2208 8.10235
R4741 VPWR.t1405 VPWR 8.10235
R4742 VPWR.t4531 VPWR 8.10235
R4743 VPWR.t5991 VPWR 8.10235
R4744 VPWR.t2363 VPWR 8.10235
R4745 VPWR.t3351 VPWR 8.10235
R4746 VPWR VPWR.t132 8.10235
R4747 VPWR VPWR.t750 8.10235
R4748 VPWR VPWR.t2706 8.10235
R4749 VPWR.t1185 VPWR.t48 8.10235
R4750 VPWR.t6286 VPWR.t6829 8.10235
R4751 VPWR.t3911 VPWR.t6390 8.10235
R4752 VPWR.t3152 VPWR 8.10235
R4753 VPWR.n103 VPWR.t6895 8.0005
R4754 VPWR.n831 VPWR.t6719 8.0005
R4755 VPWR.n739 VPWR.t13 8.0005
R4756 VPWR.n380 VPWR.t301 8.0005
R4757 VPWR.n383 VPWR.t4799 8.0005
R4758 VPWR.n1367 VPWR.t6632 7.9297
R4759 VPWR.n1368 VPWR.t5209 7.9297
R4760 VPWR.n961 VPWR.t6902 7.9297
R4761 VPWR.n706 VPWR.t5588 7.9297
R4762 VPWR.n524 VPWR.t5158 7.9297
R4763 VPWR.n893 VPWR.t6536 7.5363
R4764 VPWR.n877 VPWR.t3469 7.5363
R4765 VPWR.n861 VPWR.t6851 7.5363
R4766 VPWR.n3329 VPWR.t4092 7.5363
R4767 VPWR.n1072 VPWR.t7053 7.51784
R4768 VPWR.n1353 VPWR.t6342 7.51784
R4769 VPWR.n1625 VPWR.t6523 7.51784
R4770 VPWR.n1636 VPWR.t1693 7.51784
R4771 VPWR.n1481 VPWR.t9 7.5061
R4772 VPWR.n1416 VPWR.t6703 7.5061
R4773 VPWR.n810 VPWR.t6753 7.5061
R4774 VPWR.n1752 VPWR.t244 7.5061
R4775 VPWR.n1745 VPWR.t6841 7.5061
R4776 VPWR.n1836 VPWR.t258 7.5061
R4777 VPWR.n3755 VPWR.n61 7.4975
R4778 VPWR.n1803 VPWR.t4822 7.46
R4779 VPWR.n1805 VPWR.t6951 7.46
R4780 VPWR.n680 VPWR.t6884 7.46
R4781 VPWR.n684 VPWR.t3345 7.46
R4782 VPWR.n563 VPWR.t6419 7.46
R4783 VPWR.n567 VPWR.t4683 7.46
R4784 VPWR.n1399 VPWR.t2436 7.40883
R4785 VPWR.n1409 VPWR.t838 7.40883
R4786 VPWR.n937 VPWR.t7135 7.40883
R4787 VPWR.n948 VPWR.t4398 7.40883
R4788 VPWR.n940 VPWR.t3220 7.40883
R4789 VPWR.n931 VPWR.t3532 7.40883
R4790 VPWR.n924 VPWR.t2047 7.40883
R4791 VPWR.n1408 VPWR.t4449 7.40883
R4792 VPWR.n824 VPWR.t6306 7.40883
R4793 VPWR.n110 VPWR.t615 7.40883
R4794 VPWR.n832 VPWR.t5808 7.40883
R4795 VPWR.n751 VPWR.t3372 7.40883
R4796 VPWR.n757 VPWR.t818 7.40883
R4797 VPWR.n123 VPWR.t947 7.40883
R4798 VPWR.n3259 VPWR.t4005 7.40883
R4799 VPWR.n752 VPWR.t4110 7.40883
R4800 VPWR.n737 VPWR.t2262 7.40883
R4801 VPWR.n135 VPWR.t3873 7.40883
R4802 VPWR.n145 VPWR.t4202 7.40883
R4803 VPWR.n152 VPWR.t5858 7.40883
R4804 VPWR.n139 VPWR.t2782 7.40883
R4805 VPWR.n1784 VPWR.t2024 7.40883
R4806 VPWR.n630 VPWR.t5675 7.40883
R4807 VPWR.n1094 VPWR.t1293 7.40883
R4808 VPWR.n186 VPWR.t2891 7.40883
R4809 VPWR.n2851 VPWR.t587 7.40883
R4810 VPWR.n2875 VPWR.t5702 7.40883
R4811 VPWR.n2871 VPWR.t6263 7.40883
R4812 VPWR.n2848 VPWR.t4174 7.40883
R4813 VPWR.n2750 VPWR.t5251 7.40883
R4814 VPWR.n515 VPWR.t3254 7.40883
R4815 VPWR.n545 VPWR.t6034 7.40883
R4816 VPWR.n386 VPWR.t1906 7.40883
R4817 VPWR.n2943 VPWR.t1750 7.40883
R4818 VPWR.n387 VPWR.t1924 7.40883
R4819 VPWR.n379 VPWR.t4566 7.40883
R4820 VPWR.n1374 VPWR.t4076 7.18658
R4821 VPWR.n1380 VPWR.t1910 7.18658
R4822 VPWR.n3349 VPWR.t3638 7.18658
R4823 VPWR.n3233 VPWR.t478 7.18658
R4824 VPWR.n1730 VPWR.t3962 7.18658
R4825 VPWR.n1100 VPWR.t130 7.18658
R4826 VPWR.n1833 VPWR.t1265 7.18658
R4827 VPWR.n566 VPWR.t6586 7.18658
R4828 VPWR.n401 VPWR.t6394 7.18658
R4829 VPWR.n960 VPWR.t5021 7.16717
R4830 VPWR.n106 VPWR.t6043 7.16717
R4831 VPWR.n3270 VPWR.t408 7.16717
R4832 VPWR.n1469 VPWR.t5271 7.01851
R4833 VPWR.n3346 VPWR.t412 7.01851
R4834 VPWR.n3230 VPWR.t3993 7.01851
R4835 VPWR.n1732 VPWR.t4909 7.01851
R4836 VPWR.n1831 VPWR.t6801 7.01851
R4837 VPWR.n1024 VPWR.t5456 7.0005
R4838 VPWR.n1030 VPWR.t3240 7.0005
R4839 VPWR.n1065 VPWR.t1438 7.0005
R4840 VPWR.n1055 VPWR.t3322 7.0005
R4841 VPWR.n614 VPWR.t1789 7.0005
R4842 VPWR.n534 VPWR.t2506 7.0005
R4843 VPWR VPWR.t6871 6.94494
R4844 VPWR.t3827 VPWR 6.94494
R4845 VPWR.t3146 VPWR.t1519 6.94494
R4846 VPWR.t4902 VPWR.t5617 6.94494
R4847 VPWR.t4830 VPWR 6.94494
R4848 VPWR.t4983 VPWR.t6939 6.94494
R4849 VPWR.t6937 VPWR.t3360 6.94494
R4850 VPWR.n1093 VPWR.t3985 6.94494
R4851 VPWR.t5011 VPWR.t5747 6.94494
R4852 VPWR.t229 VPWR.t5047 6.94494
R4853 VPWR.n1078 VPWR.t1740 6.88796
R4854 VPWR.n1040 VPWR.t1527 6.88796
R4855 VPWR.n1044 VPWR.t5717 6.88796
R4856 VPWR.n1048 VPWR.t2572 6.88796
R4857 VPWR.n1356 VPWR.t4873 6.88796
R4858 VPWR.n1362 VPWR.t5934 6.88796
R4859 VPWR.n1365 VPWR.t2482 6.88796
R4860 VPWR.n1465 VPWR.t2151 6.88796
R4861 VPWR.n1352 VPWR.t3792 6.88796
R4862 VPWR.n1053 VPWR.t5663 6.88796
R4863 VPWR.n1049 VPWR.t1744 6.88796
R4864 VPWR.n1045 VPWR.t1217 6.88796
R4865 VPWR.n1043 VPWR.t1531 6.88796
R4866 VPWR.n1273 VPWR.t3280 6.88796
R4867 VPWR.n1270 VPWR.t2272 6.88796
R4868 VPWR.n1270 VPWR.t2912 6.88796
R4869 VPWR.n1266 VPWR.t3709 6.88796
R4870 VPWR.n1342 VPWR.t4380 6.88796
R4871 VPWR.n1339 VPWR.t4867 6.88796
R4872 VPWR.n1336 VPWR.t3098 6.88796
R4873 VPWR.n1310 VPWR.t1957 6.88796
R4874 VPWR.n1304 VPWR.t3506 6.88796
R4875 VPWR.n1303 VPWR.t3879 6.88796
R4876 VPWR.n1332 VPWR.t3149 6.88796
R4877 VPWR.n1338 VPWR.t919 6.88796
R4878 VPWR.n1267 VPWR.t5721 6.88796
R4879 VPWR.n1274 VPWR.t1943 6.88796
R4880 VPWR.n1227 VPWR.t2881 6.88796
R4881 VPWR.n1220 VPWR.t2182 6.88796
R4882 VPWR.n1217 VPWR.t2276 6.88796
R4883 VPWR.n1263 VPWR.t2488 6.88796
R4884 VPWR.n1257 VPWR.t3889 6.88796
R4885 VPWR.n1251 VPWR.t2226 6.88796
R4886 VPWR.n1695 VPWR.t2745 6.88796
R4887 VPWR.n1693 VPWR.t4832 6.88796
R4888 VPWR.n1706 VPWR.t4432 6.88796
R4889 VPWR.n1246 VPWR.t1068 6.88796
R4890 VPWR.n1250 VPWR.t6058 6.88796
R4891 VPWR.n1256 VPWR.t6064 6.88796
R4892 VPWR.n1218 VPWR.t1102 6.88796
R4893 VPWR.n1222 VPWR.t5625 6.88796
R4894 VPWR.n1228 VPWR.t5621 6.88796
R4895 VPWR.n1171 VPWR.t844 6.88796
R4896 VPWR.n1167 VPWR.t4480 6.88796
R4897 VPWR.n1162 VPWR.t4482 6.88796
R4898 VPWR.n1214 VPWR.t903 6.88796
R4899 VPWR.n1209 VPWR.t4279 6.88796
R4900 VPWR.n1207 VPWR.t5413 6.88796
R4901 VPWR.n1201 VPWR.t1271 6.88796
R4902 VPWR.n1716 VPWR.t4434 6.88796
R4903 VPWR.n1720 VPWR.t1049 6.88796
R4904 VPWR.n1717 VPWR.t1590 6.88796
R4905 VPWR.n1711 VPWR.t1315 6.88796
R4906 VPWR.n1179 VPWR.t1321 6.88796
R4907 VPWR.n1182 VPWR.t3061 6.88796
R4908 VPWR.n1184 VPWR.t2124 6.88796
R4909 VPWR.n1188 VPWR.t4158 6.88796
R4910 VPWR.n1192 VPWR.t1689 6.88796
R4911 VPWR.n1196 VPWR.t6244 6.88796
R4912 VPWR.n1198 VPWR.t2397 6.88796
R4913 VPWR.n1202 VPWR.t2401 6.88796
R4914 VPWR.n1206 VPWR.t1866 6.88796
R4915 VPWR.n1208 VPWR.t3585 6.88796
R4916 VPWR.n1159 VPWR.t1080 6.88796
R4917 VPWR.n1163 VPWR.t6173 6.88796
R4918 VPWR.n1166 VPWR.t7104 6.88796
R4919 VPWR.n1086 VPWR.t2524 6.88796
R4920 VPWR.n1086 VPWR.t6177 6.88796
R4921 VPWR.n1083 VPWR.t3735 6.88796
R4922 VPWR.n1083 VPWR.t5905 6.88796
R4923 VPWR.n1081 VPWR.t4511 6.88796
R4924 VPWR.n1146 VPWR.t1864 6.88796
R4925 VPWR.n1139 VPWR.t1582 6.88796
R4926 VPWR.n1135 VPWR.t1685 6.88796
R4927 VPWR.n1125 VPWR.t540 6.88796
R4928 VPWR.n1124 VPWR.t5612 6.88796
R4929 VPWR.n1131 VPWR.t538 6.88796
R4930 VPWR.n1136 VPWR.t3973 6.88796
R4931 VPWR.n1080 VPWR.t5908 6.88796
R4932 VPWR.n1990 VPWR.t5884 6.88796
R4933 VPWR.n1986 VPWR.t2998 6.88796
R4934 VPWR.n1980 VPWR.t2368 6.88796
R4935 VPWR.n1969 VPWR.t3071 6.88796
R4936 VPWR.n1966 VPWR.t5695 6.88796
R4937 VPWR.n1960 VPWR.t4414 6.88796
R4938 VPWR.n1961 VPWR.t2122 6.88796
R4939 VPWR.n1965 VPWR.t5526 6.88796
R4940 VPWR.n1977 VPWR.t5888 6.88796
R4941 VPWR.n1981 VPWR.t6253 6.88796
R4942 VPWR.n1985 VPWR.t6130 6.88796
R4943 VPWR.n1991 VPWR.t1390 6.88796
R4944 VPWR.n2134 VPWR.t5604 6.88796
R4945 VPWR.n2030 VPWR.t3175 6.88796
R4946 VPWR.n2024 VPWR.t1404 6.88796
R4947 VPWR.n2020 VPWR.t4530 6.88796
R4948 VPWR.n2720 VPWR.t607 6.88796
R4949 VPWR.n2726 VPWR.t1121 6.88796
R4950 VPWR.n2729 VPWR.t5950 6.88796
R4951 VPWR.n2725 VPWR.t5990 6.88796
R4952 VPWR.n2721 VPWR.t1127 6.88796
R4953 VPWR.n2716 VPWR.t5320 6.88796
R4954 VPWR.n2019 VPWR.t1602 6.88796
R4955 VPWR.n2023 VPWR.t2205 6.88796
R4956 VPWR.n2029 VPWR.t2207 6.88796
R4957 VPWR.n2079 VPWR.t6003 6.88796
R4958 VPWR.n2073 VPWR.t1367 6.88796
R4959 VPWR.n2069 VPWR.t5132 6.88796
R4960 VPWR.n197 VPWR.t3574 6.88796
R4961 VPWR.n2701 VPWR.t1512 6.88796
R4962 VPWR.n2697 VPWR.t1516 6.88796
R4963 VPWR.n2693 VPWR.t2915 6.88796
R4964 VPWR.n2702 VPWR.t2366 6.88796
R4965 VPWR.n2706 VPWR.t4061 6.88796
R4966 VPWR.n2070 VPWR.t4652 6.88796
R4967 VPWR.n2074 VPWR.t969 6.88796
R4968 VPWR.n2076 VPWR.t5126 6.88796
R4969 VPWR.n461 VPWR.t2825 6.88796
R4970 VPWR.n467 VPWR.t2831 6.88796
R4971 VPWR.n472 VPWR.t1638 6.88796
R4972 VPWR.n476 VPWR.t3113 6.88796
R4973 VPWR.n480 VPWR.t4143 6.88796
R4974 VPWR.n484 VPWR.t6165 6.88796
R4975 VPWR.n488 VPWR.t505 6.88796
R4976 VPWR.n493 VPWR.t1730 6.88796
R4977 VPWR.n508 VPWR.t4724 6.88796
R4978 VPWR.n502 VPWR.t5338 6.88796
R4979 VPWR.n498 VPWR.t5610 6.88796
R4980 VPWR.n1880 VPWR.t1711 6.88796
R4981 VPWR.n1880 VPWR.t2604 6.88796
R4982 VPWR.n1876 VPWR.t2603 6.88796
R4983 VPWR.n1870 VPWR.t5175 6.88796
R4984 VPWR.n1875 VPWR.t3425 6.88796
R4985 VPWR.n499 VPWR.t3339 6.88796
R4986 VPWR.n501 VPWR.t3991 6.88796
R4987 VPWR.n507 VPWR.t736 6.88796
R4988 VPWR.n509 VPWR.t1726 6.88796
R4989 VPWR.n494 VPWR.t2868 6.88796
R4990 VPWR.n491 VPWR.t4497 6.88796
R4991 VPWR.n485 VPWR.t5190 6.88796
R4992 VPWR.n481 VPWR.t511 6.88796
R4993 VPWR.n477 VPWR.t4609 6.88796
R4994 VPWR.n470 VPWR.t753 6.88796
R4995 VPWR.n466 VPWR.t1494 6.88796
R4996 VPWR.n465 VPWR.t6314 6.88796
R4997 VPWR.n1922 VPWR.t3461 6.88796
R4998 VPWR.n1918 VPWR.t311 6.88796
R4999 VPWR.n1915 VPWR.t3119 6.88796
R5000 VPWR.n1907 VPWR.t1770 6.88796
R5001 VPWR.n1899 VPWR.t3155 6.88796
R5002 VPWR.n1894 VPWR.t5828 6.88796
R5003 VPWR.n1887 VPWR.t2501 6.88796
R5004 VPWR.n453 VPWR.t2864 6.88796
R5005 VPWR.n447 VPWR.t2858 6.88796
R5006 VPWR.n443 VPWR.t3067 6.88796
R5007 VPWR.n443 VPWR.t3420 6.88796
R5008 VPWR.n446 VPWR.t5491 6.88796
R5009 VPWR.n452 VPWR.t5115 6.88796
R5010 VPWR.n1885 VPWR.t1487 6.88796
R5011 VPWR.n1892 VPWR.t4843 6.88796
R5012 VPWR.n1893 VPWR.t5783 6.88796
R5013 VPWR.n1900 VPWR.t5075 6.88796
R5014 VPWR.n1671 VPWR.t218 6.88404
R5015 VPWR.n1311 VPWR.t3565 6.88404
R5016 VPWR.n1236 VPWR.t1874 6.88404
R5017 VPWR.n1734 VPWR.t192 6.88404
R5018 VPWR.n1949 VPWR.t194 6.88404
R5019 VPWR.n1849 VPWR.t196 6.88404
R5020 VPWR.n1860 VPWR.t730 6.88404
R5021 VPWR.n111 VPWR.t1257 6.88383
R5022 VPWR.n738 VPWR.t182 6.88383
R5023 VPWR.n1095 VPWR.t728 6.88383
R5024 VPWR.n635 VPWR.t166 6.88383
R5025 VPWR.n1369 VPWR.t6271 6.8755
R5026 VPWR.n740 VPWR.t4693 6.8755
R5027 VPWR.n716 VPWR.t124 6.8755
R5028 VPWR.n607 VPWR.t1327 6.8755
R5029 VPWR.n1096 VPWR.t135 6.8755
R5030 VPWR.n1651 VPWR.t6815 6.83524
R5031 VPWR.n996 VPWR.t890 6.80877
R5032 VPWR.n799 VPWR.t1622 6.80877
R5033 VPWR.n516 VPWR.t3784 6.80352
R5034 VPWR.n950 VPWR.t4880 6.76717
R5035 VPWR.n1781 VPWR.t6858 6.76717
R5036 VPWR.n629 VPWR.t6376 6.76717
R5037 VPWR.n544 VPWR.t2579 6.76717
R5038 VPWR.n540 VPWR.t6423 6.76717
R5039 VPWR.n179 VPWR.t2705 6.76717
R5040 VPWR.n1021 VPWR.t4678 6.7505
R5041 VPWR.n1034 VPWR.t6875 6.7505
R5042 VPWR.n840 VPWR.t2355 6.7505
R5043 VPWR.n147 VPWR.t170 6.7505
R5044 VPWR.n2872 VPWR.t6421 6.7505
R5045 VPWR.n1398 VPWR.t880 6.22272
R5046 VPWR.n1407 VPWR.t5258 6.22272
R5047 VPWR.n939 VPWR.t434 6.22272
R5048 VPWR.n949 VPWR.t2381 6.22272
R5049 VPWR.n962 VPWR.t1357 6.22272
R5050 VPWR.n941 VPWR.t1778 6.22272
R5051 VPWR.n932 VPWR.t4515 6.22272
R5052 VPWR.n926 VPWR.t4656 6.22272
R5053 VPWR.n1410 VPWR.t1479 6.22272
R5054 VPWR.n825 VPWR.t1626 6.22272
R5055 VPWR.n108 VPWR.t1887 6.22272
R5056 VPWR.n109 VPWR.t1677 6.22272
R5057 VPWR.n834 VPWR.t5010 6.22272
R5058 VPWR.n753 VPWR.t2958 6.22272
R5059 VPWR.n758 VPWR.t5461 6.22272
R5060 VPWR.n3257 VPWR.t3046 6.22272
R5061 VPWR.n3271 VPWR.t6102 6.22272
R5062 VPWR.n3263 VPWR.t5986 6.22272
R5063 VPWR.n750 VPWR.t2651 6.22272
R5064 VPWR.n736 VPWR.t5791 6.22272
R5065 VPWR.n137 VPWR.t436 6.22272
R5066 VPWR.n146 VPWR.t933 6.22272
R5067 VPWR.n153 VPWR.t5090 6.22272
R5068 VPWR.n140 VPWR.t2324 6.22272
R5069 VPWR.n1785 VPWR.t461 6.22272
R5070 VPWR.n631 VPWR.t3900 6.22272
R5071 VPWR.n1090 VPWR.t2933 6.22272
R5072 VPWR.n188 VPWR.t1464 6.22272
R5073 VPWR.n2849 VPWR.t2695 6.22272
R5074 VPWR.n2877 VPWR.t2135 6.22272
R5075 VPWR.n2873 VPWR.t1834 6.22272
R5076 VPWR.n2850 VPWR.t5096 6.22272
R5077 VPWR.n2749 VPWR.t1598 6.22272
R5078 VPWR.n514 VPWR.t6158 6.22272
R5079 VPWR.n177 VPWR.t2059 6.22272
R5080 VPWR.n388 VPWR.t5553 6.22272
R5081 VPWR.n2944 VPWR.t4015 6.22272
R5082 VPWR.n389 VPWR.t465 6.22272
R5083 VPWR.n376 VPWR.t2740 6.22272
R5084 VPWR.n1063 VPWR.t7 5.9474
R5085 VPWR.n1062 VPWR.t24 5.9474
R5086 VPWR.n956 VPWR.t6497 5.9474
R5087 VPWR.n835 VPWR.t2353 5.79932
R5088 VPWR.n838 VPWR.t2347 5.79932
R5089 VPWR.n856 VPWR.t6405 5.79932
R5090 VPWR.n118 VPWR.t6411 5.79932
R5091 VPWR.n1430 VPWR.t2438 5.78954
R5092 VPWR.n1017 VPWR.t3536 5.78954
R5093 VPWR.n1620 VPWR.t2045 5.78954
R5094 VPWR.n791 VPWR.t4112 5.78954
R5095 VPWR.n1789 VPWR.t3871 5.78954
R5096 VPWR.n2837 VPWR.t2893 5.78954
R5097 VPWR.n2917 VPWR.t589 5.78954
R5098 VPWR.n2786 VPWR.t5253 5.78954
R5099 VPWR VPWR.t2283 5.78754
R5100 VPWR.t6722 VPWR.t6945 5.78754
R5101 VPWR.t17 VPWR.t6372 5.78754
R5102 VPWR VPWR.t462 5.78754
R5103 VPWR.n1394 VPWR.t3751 5.6005
R5104 VPWR.n623 VPWR.t6963 5.6005
R5105 VPWR.n538 VPWR.t5814 5.6005
R5106 VPWR.n384 VPWR.t4133 5.6005
R5107 VPWR.n1434 VPWR.n1399 5.49789
R5108 VPWR.n1420 VPWR.n1409 5.49789
R5109 VPWR.n1006 VPWR.n937 5.49789
R5110 VPWR.n990 VPWR.n948 5.49789
R5111 VPWR.n1002 VPWR.n940 5.49789
R5112 VPWR.n1014 VPWR.n931 5.49789
R5113 VPWR.n1616 VPWR.n924 5.49789
R5114 VPWR.n1421 VPWR.n1408 5.49789
R5115 VPWR.n1645 VPWR.n824 5.49789
R5116 VPWR.n3333 VPWR.n110 5.49789
R5117 VPWR.n896 VPWR.n832 5.49789
R5118 VPWR.n795 VPWR.n751 5.49789
R5119 VPWR.n780 VPWR.n757 5.49789
R5120 VPWR.n3313 VPWR.n123 5.49789
R5121 VPWR.n3302 VPWR.n3259 5.49789
R5122 VPWR.n794 VPWR.n752 5.49789
R5123 VPWR.n1682 VPWR.n737 5.49789
R5124 VPWR.n3220 VPWR.n135 5.49789
R5125 VPWR.n3202 VPWR.n145 5.49789
R5126 VPWR.n3190 VPWR.n152 5.49789
R5127 VPWR.n3211 VPWR.n139 5.49789
R5128 VPWR.n1796 VPWR.n1784 5.49789
R5129 VPWR.n670 VPWR.n630 5.49789
R5130 VPWR.n1106 VPWR.n1094 5.49789
R5131 VPWR.n2834 VPWR.n186 5.49789
R5132 VPWR.n2852 VPWR.n2851 5.49789
R5133 VPWR.n2900 VPWR.n2875 5.49789
R5134 VPWR.n2907 VPWR.n2871 5.49789
R5135 VPWR.n2855 VPWR.n2848 5.49789
R5136 VPWR.n2789 VPWR.n2750 5.49789
R5137 VPWR.n1865 VPWR.n515 5.49789
R5138 VPWR.n546 VPWR.n545 5.49789
R5139 VPWR.n413 VPWR.n386 5.49789
R5140 VPWR.n2947 VPWR.n2943 5.49789
R5141 VPWR.n412 VPWR.n387 5.49789
R5142 VPWR.n428 VPWR.n379 5.49789
R5143 VPWR.n1437 VPWR.n1398 5.41359
R5144 VPWR.n1423 VPWR.n1407 5.41359
R5145 VPWR.n1003 VPWR.n939 5.41359
R5146 VPWR.n988 VPWR.n949 5.41359
R5147 VPWR.n967 VPWR.n962 5.41359
R5148 VPWR.n1000 VPWR.n941 5.41359
R5149 VPWR.n1011 VPWR.n932 5.41359
R5150 VPWR.n1614 VPWR.n926 5.41359
R5151 VPWR.n1418 VPWR.n1410 5.41359
R5152 VPWR.n909 VPWR.n825 5.41359
R5153 VPWR.n3370 VPWR.n108 5.41359
R5154 VPWR.n3336 VPWR.n109 5.41359
R5155 VPWR.n894 VPWR.n834 5.41359
R5156 VPWR.n792 VPWR.n753 5.41359
R5157 VPWR.n777 VPWR.n758 5.41359
R5158 VPWR.n3310 VPWR.n3257 5.41359
R5159 VPWR.n3282 VPWR.n3271 5.41359
R5160 VPWR.n3300 VPWR.n3263 5.41359
R5161 VPWR.n797 VPWR.n750 5.41359
R5162 VPWR.n1684 VPWR.n736 5.41359
R5163 VPWR.n3216 VPWR.n137 5.41359
R5164 VPWR.n3200 VPWR.n146 5.41359
R5165 VPWR.n3186 VPWR.n153 5.41359
R5166 VPWR.n3208 VPWR.n140 5.41359
R5167 VPWR.n1793 VPWR.n1785 5.41359
R5168 VPWR.n666 VPWR.n631 5.41359
R5169 VPWR.n1109 VPWR.n1090 5.41359
R5170 VPWR.n189 VPWR.n188 5.41359
R5171 VPWR.n2854 VPWR.n2849 5.41359
R5172 VPWR.n2897 VPWR.n2877 5.41359
R5173 VPWR.n2904 VPWR.n2873 5.41359
R5174 VPWR.n2853 VPWR.n2850 5.41359
R5175 VPWR.n2793 VPWR.n2749 5.41359
R5176 VPWR.n1868 VPWR.n514 5.41359
R5177 VPWR.n3025 VPWR.n177 5.41359
R5178 VPWR.n411 VPWR.n388 5.41359
R5179 VPWR.n2945 VPWR.n2944 5.41359
R5180 VPWR.n410 VPWR.n389 5.41359
R5181 VPWR.n430 VPWR.n376 5.41359
R5182 VPWR.n891 VPWR.n835 5.38246
R5183 VPWR.n889 VPWR.n837 5.38246
R5184 VPWR.n888 VPWR.n838 5.38246
R5185 VPWR.n886 VPWR.n839 5.38246
R5186 VPWR.n884 VPWR.n841 5.38246
R5187 VPWR.n881 VPWR.n842 5.38246
R5188 VPWR.n879 VPWR.n843 5.38246
R5189 VPWR.n860 VPWR.n856 5.38246
R5190 VPWR.n858 VPWR.n857 5.38246
R5191 VPWR.n119 VPWR.n118 5.38246
R5192 VPWR.n3322 VPWR.n117 5.38246
R5193 VPWR.n3323 VPWR.n116 5.38246
R5194 VPWR.n3326 VPWR.n113 5.38246
R5195 VPWR.n3328 VPWR.n112 5.38246
R5196 VPWR.n1444 VPWR.n1395 5.36093
R5197 VPWR.n1331 VPWR.n1277 5.36093
R5198 VPWR.n1652 VPWR.n823 5.36093
R5199 VPWR.n1813 VPWR.n701 5.36093
R5200 VPWR.n1839 VPWR.n606 5.36093
R5201 VPWR.n1479 VPWR.n1028 5.35702
R5202 VPWR.n1074 VPWR.n1060 5.35702
R5203 VPWR.n1348 VPWR.n1039 5.35702
R5204 VPWR.n1414 VPWR.n1411 5.35702
R5205 VPWR.n1635 VPWR.n913 5.35702
R5206 VPWR.n1633 VPWR.n915 5.35702
R5207 VPWR.n1631 VPWR.n917 5.35702
R5208 VPWR.n1622 VPWR.n922 5.35702
R5209 VPWR.n1632 VPWR.n916 5.35702
R5210 VPWR.n812 VPWR.n744 5.35702
R5211 VPWR.n1746 VPWR.n713 5.35702
R5212 VPWR.n1748 VPWR.n711 5.35702
R5213 VPWR.n1750 VPWR.n709 5.35702
R5214 VPWR.n1751 VPWR.n708 5.35702
R5215 VPWR.n1749 VPWR.n710 5.35702
R5216 VPWR.n1747 VPWR.n712 5.35702
R5217 VPWR.n1832 VPWR.n610 5.35702
R5218 VPWR.n1834 VPWR.n609 5.35702
R5219 VPWR.n1835 VPWR.n608 5.35702
R5220 VPWR.n1442 VPWR.n1396 5.35271
R5221 VPWR.n1428 VPWR.n1401 5.35271
R5222 VPWR.n999 VPWR.n942 5.35271
R5223 VPWR.n984 VPWR.n951 5.35271
R5224 VPWR.n3378 VPWR.n102 5.35271
R5225 VPWR.n995 VPWR.n944 5.35271
R5226 VPWR.n1008 VPWR.n936 5.35271
R5227 VPWR.n1610 VPWR.n927 5.35271
R5228 VPWR.n1413 VPWR.n1412 5.35271
R5229 VPWR.n904 VPWR.n828 5.35271
R5230 VPWR.n3365 VPWR.n3356 5.35271
R5231 VPWR.n3351 VPWR.n3338 5.35271
R5232 VPWR.n890 VPWR.n836 5.35271
R5233 VPWR.n787 VPWR.n754 5.35271
R5234 VPWR.n772 VPWR.n759 5.35271
R5235 VPWR.n3307 VPWR.n3258 5.35271
R5236 VPWR.n3277 VPWR.n3272 5.35271
R5237 VPWR.n3295 VPWR.n3264 5.35271
R5238 VPWR.n802 VPWR.n747 5.35271
R5239 VPWR.n1689 VPWR.n734 5.35271
R5240 VPWR.n3212 VPWR.n138 5.35271
R5241 VPWR.n3194 VPWR.n148 5.35271
R5242 VPWR.n3182 VPWR.n154 5.35271
R5243 VPWR.n3204 VPWR.n144 5.35271
R5244 VPWR.n1788 VPWR.n1786 5.35271
R5245 VPWR.n661 VPWR.n633 5.35271
R5246 VPWR.n1114 VPWR.n1089 5.35271
R5247 VPWR.n1944 VPWR.n1939 5.35271
R5248 VPWR.n2858 VPWR.n2847 5.35271
R5249 VPWR.n2892 VPWR.n2878 5.35271
R5250 VPWR.n2899 VPWR.n2876 5.35271
R5251 VPWR.n2918 VPWR.n185 5.35271
R5252 VPWR.n2799 VPWR.n2747 5.35271
R5253 VPWR.n1874 VPWR.n513 5.35271
R5254 VPWR.n3031 VPWR.n174 5.35271
R5255 VPWR.n407 VPWR.n390 5.35271
R5256 VPWR.n3015 VPWR.n2954 5.35271
R5257 VPWR.n406 VPWR.n391 5.35271
R5258 VPWR.n435 VPWR.n375 5.35271
R5259 VPWR.n1511 VPWR.n1021 5.34344
R5260 VPWR.n1363 VPWR.n1034 5.34344
R5261 VPWR.n902 VPWR.n829 5.34344
R5262 VPWR.n900 VPWR.n830 5.34344
R5263 VPWR.n885 VPWR.n840 5.34344
R5264 VPWR.n1699 VPWR.n732 5.34344
R5265 VPWR.n1697 VPWR.n733 5.34344
R5266 VPWR.n1199 VPWR.n1173 5.34344
R5267 VPWR.n1183 VPWR.n1177 5.34344
R5268 VPWR.n3196 VPWR.n147 5.34344
R5269 VPWR.n2906 VPWR.n2872 5.34344
R5270 VPWR.n1456 VPWR.n1390 5.32572
R5271 VPWR.n1455 VPWR.n1391 5.32572
R5272 VPWR.n1461 VPWR.n1388 5.32572
R5273 VPWR.n1298 VPWR.n1279 5.32572
R5274 VPWR.n1298 VPWR.n1280 5.32572
R5275 VPWR.n603 VPWR.n602 5.31789
R5276 VPWR.n1850 VPWR.n522 5.31789
R5277 VPWR.n585 VPWR.n526 5.31789
R5278 VPWR.n998 VPWR.n943 5.31697
R5279 VPWR.n801 VPWR.n748 5.31697
R5280 VPWR.n1480 VPWR.n1027 5.31398
R5281 VPWR.n1073 VPWR.n1061 5.31398
R5282 VPWR.n1351 VPWR.n1037 5.31398
R5283 VPWR.n1466 VPWR.n1387 5.31398
R5284 VPWR.n1624 VPWR.n921 5.31398
R5285 VPWR.n1634 VPWR.n914 5.31398
R5286 VPWR.n1358 VPWR.n1036 5.31398
R5287 VPWR.n811 VPWR.n745 5.31398
R5288 VPWR.n809 VPWR.n746 5.31035
R5289 VPWR.n400 VPWR.n396 5.31035
R5290 VPWR.n862 VPWR.n855 5.30903
R5291 VPWR.n864 VPWR.n854 5.30903
R5292 VPWR.n1663 VPWR.n821 5.30615
R5293 VPWR.n1664 VPWR.n820 5.30615
R5294 VPWR.n3227 VPWR.n129 5.30615
R5295 VPWR.n3229 VPWR.n127 5.30615
R5296 VPWR.n3249 VPWR.n3245 5.30615
R5297 VPWR.n3250 VPWR.n3244 5.30615
R5298 VPWR.n1804 VPWR.n1780 5.30615
R5299 VPWR.n682 VPWR.n627 5.30615
R5300 VPWR.n565 VPWR.n537 5.30615
R5301 VPWR.n972 VPWR.n958 5.29976
R5302 VPWR.n3240 VPWR.n125 5.29976
R5303 VPWR.n685 VPWR.n626 5.29976
R5304 VPWR.n1853 VPWR.n520 5.29976
R5305 VPWR.n1487 VPWR.n1023 5.28785
R5306 VPWR.n1484 VPWR.n1025 5.28785
R5307 VPWR.n1032 VPWR.n1031 5.28785
R5308 VPWR.n1067 VPWR.n1066 5.28785
R5309 VPWR.n1057 VPWR.n1056 5.28785
R5310 VPWR.n1627 VPWR.n918 5.28785
R5311 VPWR.n1820 VPWR.n621 5.28785
R5312 VPWR.n582 VPWR.n528 5.28785
R5313 VPWR.n1638 VPWR.n911 5.28659
R5314 VPWR.n1731 VPWR.n723 5.28659
R5315 VPWR.n1733 VPWR.n722 5.28659
R5316 VPWR.n1735 VPWR.n721 5.28659
R5317 VPWR.n1736 VPWR.n720 5.28659
R5318 VPWR.n1738 VPWR.n719 5.28659
R5319 VPWR.n1739 VPWR.n718 5.28659
R5320 VPWR.n1741 VPWR.n717 5.28659
R5321 VPWR.n1743 VPWR.n715 5.28659
R5322 VPWR.n1772 VPWR.n1764 5.28659
R5323 VPWR.n1774 VPWR.n1762 5.28659
R5324 VPWR.n1775 VPWR.n1761 5.28659
R5325 VPWR.n1760 VPWR.n702 5.28659
R5326 VPWR.n1758 VPWR.n703 5.28659
R5327 VPWR.n1757 VPWR.n704 5.28659
R5328 VPWR.n1755 VPWR.n705 5.28659
R5329 VPWR.n1753 VPWR.n707 5.28659
R5330 VPWR.n1819 VPWR.n622 5.28659
R5331 VPWR.n1821 VPWR.n620 5.28659
R5332 VPWR.n1822 VPWR.n619 5.28659
R5333 VPWR.n1824 VPWR.n617 5.28659
R5334 VPWR.n1825 VPWR.n616 5.28659
R5335 VPWR.n1826 VPWR.n615 5.28659
R5336 VPWR.n1828 VPWR.n613 5.28659
R5337 VPWR.n1830 VPWR.n611 5.28659
R5338 VPWR.n1070 VPWR.n1063 5.27991
R5339 VPWR.n1071 VPWR.n1062 5.27991
R5340 VPWR.n977 VPWR.n956 5.27991
R5341 VPWR.n1485 VPWR.n1024 5.25874
R5342 VPWR.n1473 VPWR.n1030 5.25874
R5343 VPWR.n1068 VPWR.n1065 5.25874
R5344 VPWR.n1058 VPWR.n1055 5.25874
R5345 VPWR.n1379 VPWR.n1370 5.25874
R5346 VPWR.n1449 VPWR.n1393 5.25874
R5347 VPWR.n1448 VPWR.n1394 5.25874
R5348 VPWR.n973 VPWR.n957 5.25874
R5349 VPWR.n1377 VPWR.n1372 5.25874
R5350 VPWR.n874 VPWR.n847 5.25874
R5351 VPWR.n873 VPWR.n848 5.25874
R5352 VPWR.n871 VPWR.n850 5.25874
R5353 VPWR.n870 VPWR.n851 5.25874
R5354 VPWR.n868 VPWR.n852 5.25874
R5355 VPWR.n3344 VPWR.n3339 5.25874
R5356 VPWR.n763 VPWR.n761 5.25874
R5357 VPWR.n3289 VPWR.n3265 5.25874
R5358 VPWR.n3241 VPWR.n124 5.25874
R5359 VPWR.n1773 VPWR.n1763 5.25874
R5360 VPWR.n1769 VPWR.n1765 5.25874
R5361 VPWR.n1767 VPWR.n1766 5.25874
R5362 VPWR.n699 VPWR.n698 5.25874
R5363 VPWR.n1814 VPWR.n700 5.25874
R5364 VPWR.n1101 VPWR.n1097 5.25874
R5365 VPWR.n1840 VPWR.n605 5.25874
R5366 VPWR.n1827 VPWR.n614 5.25874
R5367 VPWR.n1823 VPWR.n618 5.25874
R5368 VPWR.n696 VPWR.n623 5.25874
R5369 VPWR.n693 VPWR.n625 5.25874
R5370 VPWR.n2915 VPWR.n2867 5.25874
R5371 VPWR.n2911 VPWR.n2870 5.25874
R5372 VPWR.n1856 VPWR.n518 5.25874
R5373 VPWR.n1854 VPWR.n519 5.25874
R5374 VPWR.n1852 VPWR.n521 5.25874
R5375 VPWR.n583 VPWR.n527 5.25874
R5376 VPWR.n581 VPWR.n529 5.25874
R5377 VPWR.n579 VPWR.n531 5.25874
R5378 VPWR.n578 VPWR.n532 5.25874
R5379 VPWR.n576 VPWR.n533 5.25874
R5380 VPWR.n568 VPWR.n536 5.25874
R5381 VPWR.n564 VPWR.n538 5.25874
R5382 VPWR.n562 VPWR.n539 5.25874
R5383 VPWR.n552 VPWR.n542 5.25874
R5384 VPWR.n575 VPWR.n534 5.25874
R5385 VPWR.n580 VPWR.n530 5.25874
R5386 VPWR.n419 VPWR.n382 5.25874
R5387 VPWR.n417 VPWR.n384 5.25874
R5388 VPWR.n399 VPWR.n397 5.25874
R5389 VPWR.n690 VPWR.t1764 5.15426
R5390 VPWR.n1098 VPWR.t5489 5.15426
R5391 VPWR.n1024 VPWR.t180 5.05606
R5392 VPWR.n1025 VPWR.t5971 5.05606
R5393 VPWR.n1030 VPWR.t7049 5.05606
R5394 VPWR.n1031 VPWR.t5520 5.05606
R5395 VPWR.n1066 VPWR.t360 5.05606
R5396 VPWR.n1065 VPWR.t53 5.05606
R5397 VPWR.n1056 VPWR.t3326 5.05606
R5398 VPWR.n1055 VPWR.t6818 5.05606
R5399 VPWR.n1398 VPWR.t4248 5.05606
R5400 VPWR.n1407 VPWR.t3159 5.05606
R5401 VPWR.n939 VPWR.t1933 5.05606
R5402 VPWR.n949 VPWR.t5232 5.05606
R5403 VPWR.n962 VPWR.t1355 5.05606
R5404 VPWR.n941 VPWR.t1618 5.05606
R5405 VPWR.n932 VPWR.t4997 5.05606
R5406 VPWR.n926 VPWR.t4938 5.05606
R5407 VPWR.n1410 VPWR.t5086 5.05606
R5408 VPWR.n825 VPWR.t2980 5.05606
R5409 VPWR.n108 VPWR.t2641 5.05606
R5410 VPWR.n109 VPWR.t4252 5.05606
R5411 VPWR.n834 VPWR.t911 5.05606
R5412 VPWR.n753 VPWR.t4570 5.05606
R5413 VPWR.n758 VPWR.t526 5.05606
R5414 VPWR.n3257 VPWR.t5358 5.05606
R5415 VPWR.n3271 VPWR.t951 5.05606
R5416 VPWR.n3263 VPWR.t1412 5.05606
R5417 VPWR.n750 VPWR.t3632 5.05606
R5418 VPWR.n736 VPWR.t5343 5.05606
R5419 VPWR.n137 VPWR.t6154 5.05606
R5420 VPWR.n146 VPWR.t2967 5.05606
R5421 VPWR.n153 VPWR.t4743 5.05606
R5422 VPWR.n140 VPWR.t3131 5.05606
R5423 VPWR.n1785 VPWR.t5643 5.05606
R5424 VPWR.n614 VPWR.t2542 5.05606
R5425 VPWR.n618 VPWR.t4979 5.05606
R5426 VPWR.n621 VPWR.t3362 5.05606
R5427 VPWR.n631 VPWR.t528 5.05606
R5428 VPWR.n1090 VPWR.t2931 5.05606
R5429 VPWR.n188 VPWR.t3236 5.05606
R5430 VPWR.n2849 VPWR.t6016 5.05606
R5431 VPWR.n2877 VPWR.t1695 5.05606
R5432 VPWR.n2873 VPWR.t4384 5.05606
R5433 VPWR.n2850 VPWR.t57 5.05606
R5434 VPWR.n2749 VPWR.t1596 5.05606
R5435 VPWR.n514 VPWR.t1020 5.05606
R5436 VPWR.n177 VPWR.t3717 5.05606
R5437 VPWR.n534 VPWR.t6959 5.05606
R5438 VPWR.n530 VPWR.t5048 5.05606
R5439 VPWR.n528 VPWR.t3831 5.05606
R5440 VPWR.n388 VPWR.t1047 5.05606
R5441 VPWR.n2944 VPWR.t4013 5.05606
R5442 VPWR.n389 VPWR.t1919 5.05606
R5443 VPWR.n376 VPWR.t943 5.05606
R5444 VPWR.n1346 VPWR.n1079 4.9415
R5445 VPWR.n1472 VPWR.n1471 4.9415
R5446 VPWR.n1488 VPWR.n817 4.9415
R5447 VPWR.n1640 VPWR.n910 4.9415
R5448 VPWR.n1606 VPWR.n1605 4.9415
R5449 VPWR.n1590 VPWR.n120 4.9415
R5450 VPWR.n3374 VPWR.n104 4.9415
R5451 VPWR.n3443 VPWR.n95 4.9415
R5452 VPWR.n1560 VPWR.n61 4.9415
R5453 VPWR.n1281 VPWR.t1959 4.89499
R5454 VPWR.n1314 VPWR.t5476 4.89499
R5455 VPWR.n1234 VPWR.t5213 4.89499
R5456 VPWR.n1737 VPWR.t5962 4.89499
R5457 VPWR.n1946 VPWR.t2647 4.89499
R5458 VPWR.n599 VPWR.t5392 4.89499
R5459 VPWR.n1857 VPWR.t3933 4.89499
R5460 VPWR.n3816 VPWR.n8 4.8515
R5461 VPWR.n3776 VPWR.n37 4.8515
R5462 VPWR.n807 VPWR.t777 4.79902
R5463 VPWR.n401 VPWR.t4685 4.79802
R5464 VPWR.n970 VPWR.t2736 4.70061
R5465 VPWR.n3242 VPWR.t4562 4.70061
R5466 VPWR.n683 VPWR.t6108 4.70061
R5467 VPWR.n1855 VPWR.t4696 4.70061
R5468 VPWR.t6408 VPWR.t6512 4.69809
R5469 VPWR.n876 VPWR.t6999 4.68691
R5470 VPWR.n1812 VPWR.t5593 4.68691
R5471 VPWR.n574 VPWR.t4987 4.68691
R5472 VPWR.n1662 VPWR.t6721 4.65756
R5473 VPWR.n3226 VPWR.t3483 4.65756
R5474 VPWR.n3248 VPWR.t6401 4.65756
R5475 VPWR.t6702 VPWR.t805 4.63013
R5476 VPWR VPWR.t6593 4.63013
R5477 VPWR.n2326 VPWR.n2325 4.63013
R5478 VPWR.n2955 VPWR.t4500 4.63013
R5479 VPWR.n3685 VPWR.t6111 4.63013
R5480 VPWR.n715 VPWR.t270 4.61026
R5481 VPWR.n707 VPWR.t6831 4.61026
R5482 VPWR.n611 VPWR.t266 4.61026
R5483 VPWR.n866 VPWR.t5141 4.51499
R5484 VPWR.n1776 VPWR.t30 4.51499
R5485 VPWR.n586 VPWR.t3019 4.51499
R5486 VPWR.n3458 VPWR.n3457 4.5005
R5487 VPWR.n3473 VPWR.n3472 4.5005
R5488 VPWR.n3488 VPWR.n3487 4.5005
R5489 VPWR.n3503 VPWR.n3502 4.5005
R5490 VPWR.n3518 VPWR.n3517 4.5005
R5491 VPWR.n3533 VPWR.n3532 4.5005
R5492 VPWR.n3548 VPWR.n3547 4.5005
R5493 VPWR.n3563 VPWR.n3562 4.5005
R5494 VPWR.n3578 VPWR.n3577 4.5005
R5495 VPWR.n3593 VPWR.n3592 4.5005
R5496 VPWR.n3608 VPWR.n3607 4.5005
R5497 VPWR.n3623 VPWR.n3622 4.5005
R5498 VPWR.n3638 VPWR.n3637 4.5005
R5499 VPWR.n3653 VPWR.n3652 4.5005
R5500 VPWR.n3668 VPWR.n3667 4.5005
R5501 VPWR.n3683 VPWR.n3682 4.5005
R5502 VPWR.n1347 VPWR.n1346 4.5005
R5503 VPWR.n1345 VPWR.n1344 4.5005
R5504 VPWR.n1265 VPWR.n1264 4.5005
R5505 VPWR.n1216 VPWR.n1215 4.5005
R5506 VPWR.n1158 VPWR.n1157 4.5005
R5507 VPWR.n2005 VPWR.n2004 4.5005
R5508 VPWR.n2101 VPWR.n2100 4.5005
R5509 VPWR.n296 VPWR.n273 4.5005
R5510 VPWR.n2394 VPWR.n2393 4.5005
R5511 VPWR.n2405 VPWR.n2404 4.5005
R5512 VPWR.n2416 VPWR.n2415 4.5005
R5513 VPWR.n2316 VPWR.n2315 4.5005
R5514 VPWR.n2278 VPWR.n2277 4.5005
R5515 VPWR.n2276 VPWR.n2275 4.5005
R5516 VPWR.n2132 VPWR.n196 4.5005
R5517 VPWR.n1974 VPWR.n195 4.5005
R5518 VPWR.n1126 VPWR.n456 4.5005
R5519 VPWR.n1710 VPWR.n1709 4.5005
R5520 VPWR.n1708 VPWR.n1707 4.5005
R5521 VPWR.n1312 VPWR.n727 4.5005
R5522 VPWR.n1471 VPWR.n1470 4.5005
R5523 VPWR.n2362 VPWR.n264 4.5005
R5524 VPWR.n2383 VPWR.n2382 4.5005
R5525 VPWR.n2343 VPWR.n259 4.5005
R5526 VPWR.n2237 VPWR.n2236 4.5005
R5527 VPWR.n2239 VPWR.n2238 4.5005
R5528 VPWR.n2185 VPWR.n2184 4.5005
R5529 VPWR.n2831 VPWR.n2830 4.5005
R5530 VPWR.n1845 VPWR.n1844 4.5005
R5531 VPWR.n1740 VPWR.n601 4.5005
R5532 VPWR.n1676 VPWR.n1675 4.5005
R5533 VPWR.n1674 VPWR.n1673 4.5005
R5534 VPWR.n1440 VPWR.n817 4.5005
R5535 VPWR.n2829 VPWR.n2828 4.5005
R5536 VPWR.n2710 VPWR.n2709 4.5005
R5537 VPWR.n2054 VPWR.n2053 4.5005
R5538 VPWR.n2797 VPWR.n183 4.5005
R5539 VPWR.n2921 VPWR.n2920 4.5005
R5540 VPWR.n1818 VPWR.n1817 4.5005
R5541 VPWR.n1816 VPWR.n1815 4.5005
R5542 VPWR.n785 VPWR.n697 4.5005
R5543 VPWR.n1642 VPWR.n1641 4.5005
R5544 VPWR.n1640 VPWR.n1639 4.5005
R5545 VPWR.n2645 VPWR.n2644 4.5005
R5546 VPWR.n2669 VPWR.n191 4.5005
R5547 VPWR.n2708 VPWR.n2707 4.5005
R5548 VPWR.n2099 VPWR.n2098 4.5005
R5549 VPWR.n219 VPWR.n3 4.5005
R5550 VPWR.n2763 VPWR.n2762 4.5005
R5551 VPWR.n2891 VPWR.n178 4.5005
R5552 VPWR.n669 VPWR.n133 4.5005
R5553 VPWR.n3222 VPWR.n3221 4.5005
R5554 VPWR.n3224 VPWR.n3223 4.5005
R5555 VPWR.n882 VPWR.n132 4.5005
R5556 VPWR.n1607 VPWR.n1606 4.5005
R5557 VPWR.n3023 VPWR.n3022 4.5005
R5558 VPWR.n577 VPWR.n182 4.5005
R5559 VPWR.n1847 VPWR.n1846 4.5005
R5560 VPWR.n1882 VPWR.n1881 4.5005
R5561 VPWR.n471 VPWR.n359 4.5005
R5562 VPWR.n3107 VPWR.n3106 4.5005
R5563 VPWR.n3109 VPWR.n3108 4.5005
R5564 VPWR.n3195 VPWR.n121 4.5005
R5565 VPWR.n3317 VPWR.n3316 4.5005
R5566 VPWR.n3319 VPWR.n3318 4.5005
R5567 VPWR.n992 VPWR.n120 4.5005
R5568 VPWR.n2990 VPWR.n8 4.5005
R5569 VPWR.n3021 VPWR.n3020 4.5005
R5570 VPWR.n2923 VPWR.n2922 4.5005
R5571 VPWR.n423 VPWR.n190 4.5005
R5572 VPWR.n1884 VPWR.n1883 4.5005
R5573 VPWR.n1925 VPWR.n1924 4.5005
R5574 VPWR.n2971 VPWR.n37 4.5005
R5575 VPWR.n3069 VPWR.n170 4.5005
R5576 VPWR.n3159 VPWR.n3158 4.5005
R5577 VPWR.n3161 VPWR.n3160 4.5005
R5578 VPWR.n3291 VPWR.n105 4.5005
R5579 VPWR.n3373 VPWR.n3372 4.5005
R5580 VPWR.n3375 VPWR.n3374 4.5005
R5581 VPWR.n3776 VPWR.n3775 4.5005
R5582 VPWR.n3817 VPWR.n3816 4.5005
R5583 VPWR.n3837 VPWR.n3836 4.5005
R5584 VPWR.n2643 VPWR.n2642 4.5005
R5585 VPWR.n2602 VPWR.n2601 4.5005
R5586 VPWR.n2501 VPWR.n2500 4.5005
R5587 VPWR.n2457 VPWR.n2456 4.5005
R5588 VPWR.n3715 VPWR.n3714 4.5005
R5589 VPWR.n3443 VPWR.n3442 4.5005
R5590 VPWR.n3717 VPWR.n3716 4.5005
R5591 VPWR.n3778 VPWR.n3777 4.5005
R5592 VPWR.n3815 VPWR.n3814 4.5005
R5593 VPWR.n3839 VPWR.n3838 4.5005
R5594 VPWR.n2575 VPWR.n255 4.5005
R5595 VPWR.n2600 VPWR.n2599 4.5005
R5596 VPWR.n2503 VPWR.n2502 4.5005
R5597 VPWR.n2455 VPWR.n2454 4.5005
R5598 VPWR.n3754 VPWR.n3753 4.5005
R5599 VPWR.n3756 VPWR.n3755 4.5005
R5600 VPWR.n3400 VPWR.n61 4.5005
R5601 VPWR.n1602 VPWR.t1201 4.49963
R5602 VPWR.n1604 VPWR.t1207 4.49963
R5603 VPWR.n1515 VPWR.t3661 4.49963
R5604 VPWR.n1513 VPWR.t3667 4.49963
R5605 VPWR.n1617 VPWR.t6332 4.49963
R5606 VPWR.n1613 VPWR.t6330 4.49963
R5607 VPWR.n1609 VPWR.t146 4.49963
R5608 VPWR.n1013 VPWR.t148 4.49963
R5609 VPWR.n1623 VPWR.t5926 4.49963
R5610 VPWR.n1628 VPWR.t5924 4.49963
R5611 VPWR.n869 VPWR.t2028 4.49963
R5612 VPWR.n875 VPWR.t2030 4.49963
R5613 VPWR.n1575 VPWR.t6904 4.46351
R5614 VPWR.n1576 VPWR.t6898 4.46351
R5615 VPWR.n1595 VPWR.t6628 4.46351
R5616 VPWR.n1596 VPWR.t6579 4.46351
R5617 VPWR.n1425 VPWR.t1055 4.46351
R5618 VPWR.n1427 VPWR.t22 4.46351
R5619 VPWR.n1433 VPWR.t3181 4.46351
R5620 VPWR.n1435 VPWR.t6027 4.46351
R5621 VPWR.n1373 VPWR.t5211 4.46351
R5622 VPWR.n1375 VPWR.t1129 4.46351
R5623 VPWR.n1319 VPWR.t6640 4.46351
R5624 VPWR.n1318 VPWR.t6878 4.46351
R5625 VPWR.n1292 VPWR.t3753 4.46351
R5626 VPWR.n1290 VPWR.t5818 4.46351
R5627 VPWR.n1672 VPWR.t226 4.46351
R5628 VPWR.n1670 VPWR.t4360 4.46351
R5629 VPWR.n1669 VPWR.t7038 4.46351
R5630 VPWR.n1667 VPWR.t3828 4.46351
R5631 VPWR.n1656 VPWR.t6799 4.46351
R5632 VPWR.n1657 VPWR.t1323 4.46351
R5633 VPWR.n1282 VPWR.t1325 4.46351
R5634 VPWR.n1284 VPWR.t524 4.46351
R5635 VPWR.n1285 VPWR.t115 4.46351
R5636 VPWR.n1287 VPWR.t2838 4.46351
R5637 VPWR.n805 VPWR.t4227 4.46351
R5638 VPWR.n803 VPWR.t6727 4.46351
R5639 VPWR.n784 VPWR.t6813 4.46351
R5640 VPWR.n786 VPWR.t3268 4.46351
R5641 VPWR.n788 VPWR.t6430 4.46351
R5642 VPWR.n790 VPWR.t4691 4.46351
R5643 VPWR.n804 VPWR.t6725 4.46351
R5644 VPWR.n806 VPWR.t5999 4.46351
R5645 VPWR.n1768 VPWR.t6590 4.46351
R5646 VPWR.n1770 VPWR.t6889 4.46351
R5647 VPWR.n688 VPWR.t5255 4.46351
R5648 VPWR.n1842 VPWR.t3773 4.46351
R5649 VPWR.n1859 VPWR.t304 4.46351
R5650 VPWR.n1858 VPWR.t3931 4.46351
R5651 VPWR.n590 VPWR.t4136 4.46351
R5652 VPWR.n591 VPWR.t5156 4.46351
R5653 VPWR.n432 VPWR.t4329 4.46351
R5654 VPWR.n431 VPWR.t4461 4.46351
R5655 VPWR.n403 VPWR.t6287 4.46351
R5656 VPWR.n402 VPWR.t3912 4.46351
R5657 VPWR.n2934 VPWR.t6581 4.46351
R5658 VPWR.n2935 VPWR.t959 4.46351
R5659 VPWR.n2924 VPWR.t6820 4.46351
R5660 VPWR.n398 VPWR.t3399 4.46351
R5661 VPWR.n1510 VPWR.t4313 4.45238
R5662 VPWR.n1366 VPWR.t6637 4.45238
R5663 VPWR.n887 VPWR.t42 4.45238
R5664 VPWR.n3193 VPWR.t6989 4.45238
R5665 VPWR.n2905 VPWR.t5566 4.45238
R5666 VPWR.n1843 VPWR.t1263 4.42047
R5667 VPWR.n584 VPWR.t6710 4.42047
R5668 VPWR.n813 VPWR.t6980 4.39118
R5669 VPWR.n2926 VPWR.t2950 4.39018
R5670 VPWR.n1550 VPWR.t2292 4.376
R5671 VPWR.n1554 VPWR.t1221 4.376
R5672 VPWR.n1556 VPWR.t321 4.376
R5673 VPWR.n1559 VPWR.t1382 4.376
R5674 VPWR.n1483 VPWR.t6749 4.36426
R5675 VPWR.n1477 VPWR.t3356 4.36426
R5676 VPWR.n1376 VPWR.t7015 4.36426
R5677 VPWR.n1436 VPWR.t6723 4.36426
R5678 VPWR.n1033 VPWR.t324 4.36426
R5679 VPWR.n1316 VPWR.t2239 4.36426
R5680 VPWR.n1315 VPWR.t6870 4.36426
R5681 VPWR.n1313 VPWR.t3836 4.36426
R5682 VPWR.n818 VPWR.t6506 4.36426
R5683 VPWR.n3348 VPWR.t6670 4.36426
R5684 VPWR.n3371 VPWR.t3222 4.36426
R5685 VPWR.n867 VPWR.t7113 4.36426
R5686 VPWR.n901 VPWR.t5870 4.36426
R5687 VPWR.n1658 VPWR.t4225 4.36426
R5688 VPWR.n1231 VPWR.t6634 4.36426
R5689 VPWR.n1683 VPWR.t18 4.36426
R5690 VPWR.n3234 VPWR.t6214 4.36426
R5691 VPWR.n1130 VPWR.t6167 4.36426
R5692 VPWR.n1848 VPWR.t3302 4.36426
R5693 VPWR.n593 VPWR.t6707 4.36426
R5694 VPWR.n557 VPWR.t6887 4.36426
R5695 VPWR.n572 VPWR.t3400 4.36426
R5696 VPWR.n434 VPWR.t4323 4.36426
R5697 VPWR.n2927 VPWR.t6822 4.36426
R5698 VPWR.n424 VPWR.t4803 4.36426
R5699 VPWR.n3446 VPWR.t1839 4.36035
R5700 VPWR.n3448 VPWR.t1211 4.36035
R5701 VPWR.n3449 VPWR.t1653 4.36035
R5702 VPWR.n3449 VPWR.t485 4.36035
R5703 VPWR.n3444 VPWR.t3429 4.36035
R5704 VPWR.n3444 VPWR.t3649 4.36035
R5705 VPWR.n3456 VPWR.t2886 4.36035
R5706 VPWR.n3456 VPWR.t2903 4.36035
R5707 VPWR.n3455 VPWR.t2823 4.36035
R5708 VPWR.n3455 VPWR.t6198 4.36035
R5709 VPWR.n3454 VPWR.t5178 4.36035
R5710 VPWR.n3454 VPWR.t2643 4.36035
R5711 VPWR.n3453 VPWR.t3270 4.36035
R5712 VPWR.n3453 VPWR.t5067 4.36035
R5713 VPWR.n3452 VPWR.t6052 4.36035
R5714 VPWR.n3452 VPWR.t3824 4.36035
R5715 VPWR.n3451 VPWR.t4858 4.36035
R5716 VPWR.n3451 VPWR.t698 4.36035
R5717 VPWR.n3447 VPWR.t3979 4.36035
R5718 VPWR.n3445 VPWR.t3806 4.36035
R5719 VPWR.n3461 VPWR.t4905 4.36035
R5720 VPWR.n3463 VPWR.t5524 4.36035
R5721 VPWR.n3464 VPWR.t1444 4.36035
R5722 VPWR.n3464 VPWR.t3257 4.36035
R5723 VPWR.n3459 VPWR.t71 4.36035
R5724 VPWR.n3459 VPWR.t3612 4.36035
R5725 VPWR.n3471 VPWR.t2186 4.36035
R5726 VPWR.n3471 VPWR.t4549 4.36035
R5727 VPWR.n3470 VPWR.t3029 4.36035
R5728 VPWR.n3470 VPWR.t3987 4.36035
R5729 VPWR.n3469 VPWR.t5522 4.36035
R5730 VPWR.n3469 VPWR.t4370 4.36035
R5731 VPWR.n3468 VPWR.t3156 4.36035
R5732 VPWR.n3468 VPWR.t963 4.36035
R5733 VPWR.n3467 VPWR.t658 4.36035
R5734 VPWR.n3467 VPWR.t6195 4.36035
R5735 VPWR.n3466 VPWR.t2282 4.36035
R5736 VPWR.n3466 VPWR.t5459 4.36035
R5737 VPWR.n3462 VPWR.t1998 4.36035
R5738 VPWR.n3460 VPWR.t1334 4.36035
R5739 VPWR.n3476 VPWR.t4386 4.36035
R5740 VPWR.n3478 VPWR.t2388 4.36035
R5741 VPWR.n3479 VPWR.t4977 4.36035
R5742 VPWR.n3479 VPWR.t558 4.36035
R5743 VPWR.n3474 VPWR.t4554 4.36035
R5744 VPWR.n3474 VPWR.t1140 4.36035
R5745 VPWR.n3486 VPWR.t6357 4.36035
R5746 VPWR.n3486 VPWR.t3498 4.36035
R5747 VPWR.n3485 VPWR.t5698 4.36035
R5748 VPWR.n3485 VPWR.t1359 4.36035
R5749 VPWR.n3484 VPWR.t621 4.36035
R5750 VPWR.n3484 VPWR.t5676 4.36035
R5751 VPWR.n3483 VPWR.t2402 4.36035
R5752 VPWR.n3483 VPWR.t1398 4.36035
R5753 VPWR.n3482 VPWR.t6229 4.36035
R5754 VPWR.n3482 VPWR.t4418 4.36035
R5755 VPWR.n3481 VPWR.t1014 4.36035
R5756 VPWR.n3481 VPWR.t5344 4.36035
R5757 VPWR.n3477 VPWR.t430 4.36035
R5758 VPWR.n3475 VPWR.t7130 4.36035
R5759 VPWR.n3491 VPWR.t4628 4.36035
R5760 VPWR.n3493 VPWR.t2112 4.36035
R5761 VPWR.n3494 VPWR.t1446 4.36035
R5762 VPWR.n3494 VPWR.t5879 4.36035
R5763 VPWR.n3489 VPWR.t7082 4.36035
R5764 VPWR.n3489 VPWR.t5197 4.36035
R5765 VPWR.n3501 VPWR.t2741 4.36035
R5766 VPWR.n3501 VPWR.t422 4.36035
R5767 VPWR.n3500 VPWR.t3100 4.36035
R5768 VPWR.n3500 VPWR.t3558 4.36035
R5769 VPWR.n3499 VPWR.t3966 4.36035
R5770 VPWR.n3499 VPWR.t4910 4.36035
R5771 VPWR.n3498 VPWR.t3861 4.36035
R5772 VPWR.n3498 VPWR.t2670 4.36035
R5773 VPWR.n3497 VPWR.t426 4.36035
R5774 VPWR.n3497 VPWR.t3491 4.36035
R5775 VPWR.n3496 VPWR.t2821 4.36035
R5776 VPWR.n3496 VPWR.t1900 4.36035
R5777 VPWR.n3492 VPWR.t3287 4.36035
R5778 VPWR.n3490 VPWR.t4703 4.36035
R5779 VPWR.n3506 VPWR.t4493 4.36035
R5780 VPWR.n3508 VPWR.t2672 4.36035
R5781 VPWR.n3509 VPWR.t6152 4.36035
R5782 VPWR.n3509 VPWR.t2008 4.36035
R5783 VPWR.n3504 VPWR.t4780 4.36035
R5784 VPWR.n3504 VPWR.t3090 4.36035
R5785 VPWR.n3516 VPWR.t3820 4.36035
R5786 VPWR.n3516 VPWR.t4030 4.36035
R5787 VPWR.n3515 VPWR.t2316 4.36035
R5788 VPWR.n3515 VPWR.t1299 4.36035
R5789 VPWR.n3514 VPWR.t642 4.36035
R5790 VPWR.n3514 VPWR.t5109 4.36035
R5791 VPWR.n3513 VPWR.t3289 4.36035
R5792 VPWR.n3513 VPWR.t4629 4.36035
R5793 VPWR.n3512 VPWR.t6070 4.36035
R5794 VPWR.n3512 VPWR.t4761 4.36035
R5795 VPWR.n3511 VPWR.t329 4.36035
R5796 VPWR.n3511 VPWR.t3986 4.36035
R5797 VPWR.n3507 VPWR.t1836 4.36035
R5798 VPWR.n3505 VPWR.t1523 4.36035
R5799 VPWR.n3521 VPWR.t4114 4.36035
R5800 VPWR.n3523 VPWR.t2788 4.36035
R5801 VPWR.n3524 VPWR.t2339 4.36035
R5802 VPWR.n3524 VPWR.t3212 4.36035
R5803 VPWR.n3519 VPWR.t4293 4.36035
R5804 VPWR.n3519 VPWR.t3034 4.36035
R5805 VPWR.n3531 VPWR.t7080 4.36035
R5806 VPWR.n3531 VPWR.t5640 4.36035
R5807 VPWR.n3530 VPWR.t6433 4.36035
R5808 VPWR.n3530 VPWR.t4261 4.36035
R5809 VPWR.n3529 VPWR.t559 4.36035
R5810 VPWR.n3529 VPWR.t317 4.36035
R5811 VPWR.n3528 VPWR.t1142 4.36035
R5812 VPWR.n3528 VPWR.t5560 4.36035
R5813 VPWR.n3527 VPWR.t5091 4.36035
R5814 VPWR.n3527 VPWR.t2298 4.36035
R5815 VPWR.n3526 VPWR.t3541 4.36035
R5816 VPWR.n3526 VPWR.t3995 4.36035
R5817 VPWR.n3522 VPWR.t1136 4.36035
R5818 VPWR.n3520 VPWR.t7074 4.36035
R5819 VPWR.n3536 VPWR.t2666 4.36035
R5820 VPWR.n3538 VPWR.t2330 4.36035
R5821 VPWR.n3539 VPWR.t3405 4.36035
R5822 VPWR.n3539 VPWR.t1076 4.36035
R5823 VPWR.n3534 VPWR.t6028 4.36035
R5824 VPWR.n3534 VPWR.t5799 4.36035
R5825 VPWR.n3546 VPWR.t1814 4.36035
R5826 VPWR.n3546 VPWR.t5390 4.36035
R5827 VPWR.n3545 VPWR.t366 4.36035
R5828 VPWR.n3545 VPWR.t3233 4.36035
R5829 VPWR.n3544 VPWR.t2514 4.36035
R5830 VPWR.n3544 VPWR.t4003 4.36035
R5831 VPWR.n3543 VPWR.t2986 4.36035
R5832 VPWR.n3543 VPWR.t2897 4.36035
R5833 VPWR.n3542 VPWR.t1394 4.36035
R5834 VPWR.n3542 VPWR.t2848 4.36035
R5835 VPWR.n3541 VPWR.t69 4.36035
R5836 VPWR.n3541 VPWR.t624 4.36035
R5837 VPWR.n3537 VPWR.t3651 4.36035
R5838 VPWR.n3535 VPWR.t4420 4.36035
R5839 VPWR.n3551 VPWR.t1746 4.36035
R5840 VPWR.n3553 VPWR.t4973 4.36035
R5841 VPWR.n3554 VPWR.t927 4.36035
R5842 VPWR.n3554 VPWR.t2303 4.36035
R5843 VPWR.n3549 VPWR.t7087 4.36035
R5844 VPWR.n3549 VPWR.t5243 4.36035
R5845 VPWR.n3561 VPWR.t2180 4.36035
R5846 VPWR.n3561 VPWR.t4348 4.36035
R5847 VPWR.n3560 VPWR.t3167 4.36035
R5848 VPWR.n3560 VPWR.t4408 4.36035
R5849 VPWR.n3559 VPWR.t5712 4.36035
R5850 VPWR.n3559 VPWR.t6309 4.36035
R5851 VPWR.n3558 VPWR.t2962 4.36035
R5852 VPWR.n3558 VPWR.t6096 4.36035
R5853 VPWR.n3557 VPWR.t2414 4.36035
R5854 VPWR.n3557 VPWR.t5743 4.36035
R5855 VPWR.n3556 VPWR.t4068 4.36035
R5856 VPWR.n3556 VPWR.t1062 4.36035
R5857 VPWR.n3552 VPWR.t2850 4.36035
R5858 VPWR.n3550 VPWR.t2189 4.36035
R5859 VPWR.n3566 VPWR.t2617 4.36035
R5860 VPWR.n3568 VPWR.t1734 4.36035
R5861 VPWR.n3569 VPWR.t6232 4.36035
R5862 VPWR.n3569 VPWR.t2118 4.36035
R5863 VPWR.n3564 VPWR.t3693 4.36035
R5864 VPWR.n3564 VPWR.t1971 4.36035
R5865 VPWR.n3576 VPWR.t874 4.36035
R5866 VPWR.n3576 VPWR.t4588 4.36035
R5867 VPWR.n3575 VPWR.t2302 4.36035
R5868 VPWR.n3575 VPWR.t1568 4.36035
R5869 VPWR.n3574 VPWR.t1086 4.36035
R5870 VPWR.n3574 VPWR.t4246 4.36035
R5871 VPWR.n3573 VPWR.t5371 4.36035
R5872 VPWR.n3573 VPWR.t2040 4.36035
R5873 VPWR.n3572 VPWR.t5733 4.36035
R5874 VPWR.n3572 VPWR.t1242 4.36035
R5875 VPWR.n3571 VPWR.t3341 4.36035
R5876 VPWR.n3571 VPWR.t4194 4.36035
R5877 VPWR.n3567 VPWR.t5370 4.36035
R5878 VPWR.n3565 VPWR.t517 4.36035
R5879 VPWR.n3581 VPWR.t3465 4.36035
R5880 VPWR.n3583 VPWR.t2743 4.36035
R5881 VPWR.n3584 VPWR.t5207 4.36035
R5882 VPWR.n3584 VPWR.t3053 4.36035
R5883 VPWR.n3579 VPWR.t802 4.36035
R5884 VPWR.n3579 VPWR.t3982 4.36035
R5885 VPWR.n3591 VPWR.t5789 4.36035
R5886 VPWR.n3591 VPWR.t3757 4.36035
R5887 VPWR.n3590 VPWR.t4660 4.36035
R5888 VPWR.n3590 VPWR.t3909 4.36035
R5889 VPWR.n3589 VPWR.t1931 4.36035
R5890 VPWR.n3589 VPWR.t694 4.36035
R5891 VPWR.n3588 VPWR.t1291 4.36035
R5892 VPWR.n3588 VPWR.t4317 4.36035
R5893 VPWR.n3587 VPWR.t3863 4.36035
R5894 VPWR.n3587 VPWR.t2217 4.36035
R5895 VPWR.n3586 VPWR.t2110 4.36035
R5896 VPWR.n3586 VPWR.t4773 4.36035
R5897 VPWR.n3582 VPWR.t5290 4.36035
R5898 VPWR.n3580 VPWR.t5467 4.36035
R5899 VPWR.n3596 VPWR.t1784 4.36035
R5900 VPWR.n3598 VPWR.t7102 4.36035
R5901 VPWR.n3599 VPWR.t6212 4.36035
R5902 VPWR.n3599 VPWR.t2234 4.36035
R5903 VPWR.n3594 VPWR.t2866 4.36035
R5904 VPWR.n3594 VPWR.t3923 4.36035
R5905 VPWR.n3606 VPWR.t2391 4.36035
R5906 VPWR.n3606 VPWR.t5053 4.36035
R5907 VPWR.n3605 VPWR.t3048 4.36035
R5908 VPWR.n3605 VPWR.t3078 4.36035
R5909 VPWR.n3604 VPWR.t55 4.36035
R5910 VPWR.n3604 VPWR.t3862 4.36035
R5911 VPWR.n3603 VPWR.t3106 4.36035
R5912 VPWR.n3603 VPWR.t2699 4.36035
R5913 VPWR.n3602 VPWR.t5278 4.36035
R5914 VPWR.n3602 VPWR.t1858 4.36035
R5915 VPWR.n3601 VPWR.t5419 4.36035
R5916 VPWR.n3601 VPWR.t4584 4.36035
R5917 VPWR.n3597 VPWR.t6068 4.36035
R5918 VPWR.n3595 VPWR.t1624 4.36035
R5919 VPWR.n3611 VPWR.t3261 4.36035
R5920 VPWR.n3613 VPWR.t2786 4.36035
R5921 VPWR.n3614 VPWR.t2944 4.36035
R5922 VPWR.n3614 VPWR.t4161 4.36035
R5923 VPWR.n3609 VPWR.t1027 4.36035
R5924 VPWR.n3609 VPWR.t3201 4.36035
R5925 VPWR.n3621 VPWR.t1988 4.36035
R5926 VPWR.n3621 VPWR.t3368 4.36035
R5927 VPWR.n3620 VPWR.t6351 4.36035
R5928 VPWR.n3620 VPWR.t3956 4.36035
R5929 VPWR.n3619 VPWR.t4642 4.36035
R5930 VPWR.n3619 VPWR.t1353 4.36035
R5931 VPWR.n3618 VPWR.t4787 4.36035
R5932 VPWR.n3618 VPWR.t1801 4.36035
R5933 VPWR.n3617 VPWR.t1898 4.36035
R5934 VPWR.n3617 VPWR.t2003 4.36035
R5935 VPWR.n3616 VPWR.t3595 4.36035
R5936 VPWR.n3616 VPWR.t4520 4.36035
R5937 VPWR.n3612 VPWR.t4786 4.36035
R5938 VPWR.n3610 VPWR.t1307 4.36035
R5939 VPWR.n3626 VPWR.t2406 4.36035
R5940 VPWR.n3628 VPWR.t3925 4.36035
R5941 VPWR.n3629 VPWR.t3189 4.36035
R5942 VPWR.n3629 VPWR.t5076 4.36035
R5943 VPWR.n3624 VPWR.t6345 4.36035
R5944 VPWR.n3624 VPWR.t3407 4.36035
R5945 VPWR.n3636 VPWR.t2389 4.36035
R5946 VPWR.n3636 VPWR.t648 4.36035
R5947 VPWR.n3635 VPWR.t4233 4.36035
R5948 VPWR.n3635 VPWR.t2726 4.36035
R5949 VPWR.n3634 VPWR.t4081 4.36035
R5950 VPWR.n3634 VPWR.t4001 4.36035
R5951 VPWR.n3633 VPWR.t1982 4.36035
R5952 VPWR.n3633 VPWR.t3488 4.36035
R5953 VPWR.n3632 VPWR.t2565 4.36035
R5954 VPWR.n3632 VPWR.t4355 4.36035
R5955 VPWR.n3631 VPWR.t4884 4.36035
R5956 VPWR.n3631 VPWR.t5788 4.36035
R5957 VPWR.n3627 VPWR.t4116 4.36035
R5958 VPWR.n3625 VPWR.t3216 4.36035
R5959 VPWR.n3641 VPWR.t6076 4.36035
R5960 VPWR.n3643 VPWR.t81 4.36035
R5961 VPWR.n3644 VPWR.t743 4.36035
R5962 VPWR.n3644 VPWR.t1920 4.36035
R5963 VPWR.n3639 VPWR.t4245 4.36035
R5964 VPWR.n3639 VPWR.t5865 4.36035
R5965 VPWR.n3651 VPWR.t374 4.36035
R5966 VPWR.n3651 VPWR.t4150 4.36035
R5967 VPWR.n3650 VPWR.t5346 4.36035
R5968 VPWR.n3650 VPWR.t6355 4.36035
R5969 VPWR.n3649 VPWR.t4533 4.36035
R5970 VPWR.n3649 VPWR.t792 4.36035
R5971 VPWR.n3648 VPWR.t3 4.36035
R5972 VPWR.n3648 VPWR.t659 4.36035
R5973 VPWR.n3647 VPWR.t6115 4.36035
R5974 VPWR.n3647 VPWR.t6455 4.36035
R5975 VPWR.n3646 VPWR.t4585 4.36035
R5976 VPWR.n3646 VPWR.t483 4.36035
R5977 VPWR.n3642 VPWR.t5314 4.36035
R5978 VPWR.n3640 VPWR.t3604 4.36035
R5979 VPWR.n3656 VPWR.t5534 4.36035
R5980 VPWR.n3658 VPWR.t3723 4.36035
R5981 VPWR.n3659 VPWR.t3445 4.36035
R5982 VPWR.n3659 VPWR.t2583 4.36035
R5983 VPWR.n3654 VPWR.t1189 4.36035
R5984 VPWR.n3654 VPWR.t6019 4.36035
R5985 VPWR.n3666 VPWR.t6816 4.36035
R5986 VPWR.n3666 VPWR.t2755 4.36035
R5987 VPWR.n3665 VPWR.t781 4.36035
R5988 VPWR.n3665 VPWR.t2187 4.36035
R5989 VPWR.n3664 VPWR.t3105 4.36035
R5990 VPWR.n3664 VPWR.t3901 4.36035
R5991 VPWR.n3663 VPWR.t2244 4.36035
R5992 VPWR.n3663 VPWR.t747 4.36035
R5993 VPWR.n3662 VPWR.t3745 4.36035
R5994 VPWR.n3662 VPWR.t4548 4.36035
R5995 VPWR.n3661 VPWR.t2611 4.36035
R5996 VPWR.n3661 VPWR.t3639 4.36035
R5997 VPWR.n3657 VPWR.t3721 4.36035
R5998 VPWR.n3655 VPWR.t4218 4.36035
R5999 VPWR.n3671 VPWR.t5551 4.36035
R6000 VPWR.n3673 VPWR.t4347 4.36035
R6001 VPWR.n3674 VPWR.t1378 4.36035
R6002 VPWR.n3674 VPWR.t3442 4.36035
R6003 VPWR.n3669 VPWR.t5465 4.36035
R6004 VPWR.n3669 VPWR.t6207 4.36035
R6005 VPWR.n3681 VPWR.t4168 4.36035
R6006 VPWR.n3681 VPWR.t5898 4.36035
R6007 VPWR.n3680 VPWR.t4366 4.36035
R6008 VPWR.n3680 VPWR.t3040 4.36035
R6009 VPWR.n3679 VPWR.t384 4.36035
R6010 VPWR.n3679 VPWR.t1915 4.36035
R6011 VPWR.n3678 VPWR.t3453 4.36035
R6012 VPWR.n3678 VPWR.t1363 4.36035
R6013 VPWR.n3677 VPWR.t1460 4.36035
R6014 VPWR.n3677 VPWR.t2907 4.36035
R6015 VPWR.n3676 VPWR.t1758 4.36035
R6016 VPWR.n3676 VPWR.t6021 4.36035
R6017 VPWR.n3672 VPWR.t2169 4.36035
R6018 VPWR.n3670 VPWR.t3838 4.36035
R6019 VPWR.n1541 VPWR.t4243 4.36035
R6020 VPWR.n1540 VPWR.t2835 4.36035
R6021 VPWR.n1539 VPWR.t654 4.36035
R6022 VPWR.n1538 VPWR.t4893 4.36035
R6023 VPWR.n1537 VPWR.t2290 4.36035
R6024 VPWR.n1536 VPWR.t351 4.36035
R6025 VPWR.n1543 VPWR.t5401 4.36035
R6026 VPWR.n1544 VPWR.t6117 4.36035
R6027 VPWR.n1546 VPWR.t5635 4.36035
R6028 VPWR.n1547 VPWR.t859 4.36035
R6029 VPWR.n1548 VPWR.t3766 4.36035
R6030 VPWR.n1549 VPWR.t4343 4.36035
R6031 VPWR.n1551 VPWR.t1029 4.36035
R6032 VPWR.n1552 VPWR.t1705 4.36035
R6033 VPWR.n1555 VPWR.t2759 4.36035
R6034 VPWR.n1557 VPWR.t1132 4.36035
R6035 VPWR.n1558 VPWR.t3941 4.36035
R6036 VPWR.n1561 VPWR.t2629 4.36035
R6037 VPWR.n1564 VPWR.t1408 4.36035
R6038 VPWR.n1565 VPWR.t2446 4.36035
R6039 VPWR.n1567 VPWR.t544 4.36035
R6040 VPWR.n1568 VPWR.t1841 4.36035
R6041 VPWR.n1533 VPWR.t2318 4.36035
R6042 VPWR.n1531 VPWR.t1904 4.36035
R6043 VPWR.n1530 VPWR.t3108 4.36035
R6044 VPWR.n1529 VPWR.t2294 4.36035
R6045 VPWR.n1528 VPWR.t2082 4.36035
R6046 VPWR.n1527 VPWR.t4581 4.36035
R6047 VPWR.n1577 VPWR.t1313 4.36035
R6048 VPWR.n1578 VPWR.t848 4.36035
R6049 VPWR.n1579 VPWR.t5351 4.36035
R6050 VPWR.n1580 VPWR.t546 4.36035
R6051 VPWR.n1581 VPWR.t5318 4.36035
R6052 VPWR.n1584 VPWR.t1660 4.36035
R6053 VPWR.n1585 VPWR.t6200 4.36035
R6054 VPWR.n1587 VPWR.t4154 4.36035
R6055 VPWR.n1588 VPWR.t2585 4.36035
R6056 VPWR.n1589 VPWR.t779 4.36035
R6057 VPWR.n1597 VPWR.t1233 4.36035
R6058 VPWR.n1600 VPWR.t2288 4.36035
R6059 VPWR.n1516 VPWR.t1164 4.36035
R6060 VPWR.n1517 VPWR.t2761 4.36035
R6061 VPWR.n1498 VPWR.t5495 4.36035
R6062 VPWR.n1499 VPWR.t720 4.36035
R6063 VPWR.n1500 VPWR.t5918 4.36035
R6064 VPWR.n1501 VPWR.t5981 4.36035
R6065 VPWR.n1502 VPWR.t3282 4.36035
R6066 VPWR.n1503 VPWR.t4284 4.36035
R6067 VPWR.n1504 VPWR.t623 4.36035
R6068 VPWR.n1505 VPWR.t7128 4.36035
R6069 VPWR.n1497 VPWR.t5549 4.36035
R6070 VPWR.n1496 VPWR.t1953 4.36035
R6071 VPWR.n1495 VPWR.t5298 4.36035
R6072 VPWR.n1494 VPWR.t5430 4.36035
R6073 VPWR.n1493 VPWR.t5530 4.36035
R6074 VPWR.n1492 VPWR.t2969 4.36035
R6075 VPWR.n1491 VPWR.t3065 4.36035
R6076 VPWR.n1490 VPWR.t1152 4.36035
R6077 VPWR.n1476 VPWR.t4829 4.36035
R6078 VPWR.n1076 VPWR.t5284 4.36035
R6079 VPWR.n1354 VPWR.t5657 4.36035
R6080 VPWR.n1417 VPWR.t3125 4.36035
R6081 VPWR.n982 VPWR.t6447 4.36035
R6082 VPWR.n980 VPWR.t4495 4.36035
R6083 VPWR.n3379 VPWR.t4118 4.36035
R6084 VPWR.n3381 VPWR.t6362 4.36035
R6085 VPWR.n3382 VPWR.t3075 4.36035
R6086 VPWR.n3382 VPWR.t7133 4.36035
R6087 VPWR.n3383 VPWR.t2871 4.36035
R6088 VPWR.n3383 VPWR.t2404 4.36035
R6089 VPWR.n3386 VPWR.t4259 4.36035
R6090 VPWR.n3388 VPWR.t3843 4.36035
R6091 VPWR.n3388 VPWR.t79 4.36035
R6092 VPWR.n3389 VPWR.t3502 4.36035
R6093 VPWR.n3389 VPWR.t7081 4.36035
R6094 VPWR.n3390 VPWR.t4426 4.36035
R6095 VPWR.n3390 VPWR.t656 4.36035
R6096 VPWR.n3391 VPWR.t5749 4.36035
R6097 VPWR.n3391 VPWR.t1548 4.36035
R6098 VPWR.n3392 VPWR.t4729 4.36035
R6099 VPWR.n3392 VPWR.t3786 4.36035
R6100 VPWR.n3393 VPWR.t6233 4.36035
R6101 VPWR.n3393 VPWR.t5573 4.36035
R6102 VPWR.n3394 VPWR.t1219 4.36035
R6103 VPWR.n3394 VPWR.t7071 4.36035
R6104 VPWR.n3395 VPWR.t1917 4.36035
R6105 VPWR.n3395 VPWR.t6451 4.36035
R6106 VPWR.n3396 VPWR.t708 4.36035
R6107 VPWR.n3399 VPWR.t1246 4.36035
R6108 VPWR.n3402 VPWR.t3314 4.36035
R6109 VPWR.n3404 VPWR.t1231 4.36035
R6110 VPWR.n3406 VPWR.t5137 4.36035
R6111 VPWR.n3408 VPWR.t696 4.36035
R6112 VPWR.n3410 VPWR.t443 4.36035
R6113 VPWR.n3412 VPWR.t1462 4.36035
R6114 VPWR.n3415 VPWR.t6443 4.36035
R6115 VPWR.n3418 VPWR.t376 4.36035
R6116 VPWR.n3420 VPWR.t2548 4.36035
R6117 VPWR.n3422 VPWR.t5795 4.36035
R6118 VPWR.n3424 VPWR.t1197 4.36035
R6119 VPWR.n3426 VPWR.t2775 4.36035
R6120 VPWR.n3428 VPWR.t7078 4.36035
R6121 VPWR.n3430 VPWR.t4507 4.36035
R6122 VPWR.n3432 VPWR.t755 4.36035
R6123 VPWR.n3433 VPWR.t3431 4.36035
R6124 VPWR.n3433 VPWR.t5765 4.36035
R6125 VPWR.n96 VPWR.t4286 4.36035
R6126 VPWR.n96 VPWR.t4968 4.36035
R6127 VPWR.n3441 VPWR.t3743 4.36035
R6128 VPWR.n3441 VPWR.t5101 4.36035
R6129 VPWR.n3440 VPWR.t1608 4.36035
R6130 VPWR.n3440 VPWR.t6439 4.36035
R6131 VPWR.n3439 VPWR.t2664 4.36035
R6132 VPWR.n3439 VPWR.t5418 4.36035
R6133 VPWR.n3438 VPWR.t2000 4.36035
R6134 VPWR.n3438 VPWR.t4620 4.36035
R6135 VPWR.n3437 VPWR.t3957 4.36035
R6136 VPWR.n3437 VPWR.t2016 4.36035
R6137 VPWR.n3436 VPWR.t5513 4.36035
R6138 VPWR.n3436 VPWR.t87 4.36035
R6139 VPWR.n3431 VPWR.t3209 4.36035
R6140 VPWR.n3429 VPWR.t6171 4.36035
R6141 VPWR.n3427 VPWR.t5263 4.36035
R6142 VPWR.n3425 VPWR.t3702 4.36035
R6143 VPWR.n3423 VPWR.t5432 4.36035
R6144 VPWR.n3421 VPWR.t5240 4.36035
R6145 VPWR.n3419 VPWR.t5180 4.36035
R6146 VPWR.n3417 VPWR.t4471 4.36035
R6147 VPWR.n3413 VPWR.t2800 4.36035
R6148 VPWR.n3411 VPWR.t6072 4.36035
R6149 VPWR.n3409 VPWR.t3367 4.36035
R6150 VPWR.n3407 VPWR.t6285 4.36035
R6151 VPWR.n3405 VPWR.t1154 4.36035
R6152 VPWR.n3403 VPWR.t3999 4.36035
R6153 VPWR.n3401 VPWR.t1458 4.36035
R6154 VPWR.n3398 VPWR.t3920 4.36035
R6155 VPWR.n3384 VPWR.t5417 4.36035
R6156 VPWR.n974 VPWR.t2171 4.36035
R6157 VPWR.n976 VPWR.t6190 4.36035
R6158 VPWR.n978 VPWR.t5261 4.36035
R6159 VPWR.n979 VPWR.t3015 4.36035
R6160 VPWR.n1438 VPWR.t4256 4.36035
R6161 VPWR.n1464 VPWR.t4273 4.36035
R6162 VPWR.n1343 VPWR.t6025 4.36035
R6163 VPWR.n1323 VPWR.t3316 4.36035
R6164 VPWR.n1321 VPWR.t5057 4.36035
R6165 VPWR.n1302 VPWR.t3457 4.36035
R6166 VPWR.n1302 VPWR.t3698 4.36035
R6167 VPWR.n1301 VPWR.t5598 4.36035
R6168 VPWR.n1301 VPWR.t2522 4.36035
R6169 VPWR.n1300 VPWR.t1150 4.36035
R6170 VPWR.n1300 VPWR.t3764 4.36035
R6171 VPWR.n1283 VPWR.t5194 4.36035
R6172 VPWR.n1654 VPWR.t4229 4.36035
R6173 VPWR.n1653 VPWR.t5633 4.36035
R6174 VPWR.n3335 VPWR.t6321 4.36035
R6175 VPWR.n3337 VPWR.t2751 4.36035
R6176 VPWR.n3350 VPWR.t1699 4.36035
R6177 VPWR.n3363 VPWR.t634 4.36035
R6178 VPWR.n3363 VPWR.t2178 4.36035
R6179 VPWR.n3362 VPWR.t5916 4.36035
R6180 VPWR.n3362 VPWR.t2873 4.36035
R6181 VPWR.n3361 VPWR.t4755 4.36035
R6182 VPWR.n3361 VPWR.t2621 4.36035
R6183 VPWR.n3360 VPWR.t4630 4.36035
R6184 VPWR.n3360 VPWR.t1166 4.36035
R6185 VPWR.n3359 VPWR.t5774 4.36035
R6186 VPWR.n3359 VPWR.t4178 4.36035
R6187 VPWR.n3364 VPWR.t2326 4.36035
R6188 VPWR.n3367 VPWR.t5545 4.36035
R6189 VPWR.n3368 VPWR.t3893 4.36035
R6190 VPWR.n3341 VPWR.t3450 4.36035
R6191 VPWR.n3343 VPWR.t1600 4.36035
R6192 VPWR.n3345 VPWR.t5396 4.36035
R6193 VPWR.n3325 VPWR.t4388 4.36035
R6194 VPWR.n3321 VPWR.t882 4.36035
R6195 VPWR.n3320 VPWR.t5753 4.36035
R6196 VPWR.n899 VPWR.t5356 4.36035
R6197 VPWR.n903 VPWR.t5169 4.36035
R6198 VPWR.n905 VPWR.t5497 4.36035
R6199 VPWR.n908 VPWR.t3417 4.36035
R6200 VPWR.n1643 VPWR.t6126 4.36035
R6201 VPWR.n1644 VPWR.t3147 4.36035
R6202 VPWR.n1646 VPWR.t3749 4.36035
R6203 VPWR.n1648 VPWR.t5706 4.36035
R6204 VPWR.n1650 VPWR.t5398 4.36035
R6205 VPWR.n1289 VPWR.t5804 4.36035
R6206 VPWR.n1291 VPWR.t5443 4.36035
R6207 VPWR.n1293 VPWR.t4611 4.36035
R6208 VPWR.n1296 VPWR.t4469 4.36035
R6209 VPWR.n1307 VPWR.t3810 4.36035
R6210 VPWR.n1320 VPWR.t353 4.36035
R6211 VPWR.n1322 VPWR.t2902 4.36035
R6212 VPWR.n1324 VPWR.t5659 4.36035
R6213 VPWR.n1326 VPWR.t4524 4.36035
R6214 VPWR.n1328 VPWR.t2051 4.36035
R6215 VPWR.n1329 VPWR.t1826 4.36035
R6216 VPWR.n1330 VPWR.t901 4.36035
R6217 VPWR.n1335 VPWR.t5385 4.36035
R6218 VPWR.n1259 VPWR.t2428 4.36035
R6219 VPWR.n1249 VPWR.t4967 4.36035
R6220 VPWR.n1247 VPWR.t3435 4.36035
R6221 VPWR.n1244 VPWR.t4193 4.36035
R6222 VPWR.n1242 VPWR.t1876 4.36035
R6223 VPWR.n1238 VPWR.t5353 4.36035
R6224 VPWR.n1233 VPWR.t5469 4.36035
R6225 VPWR.n728 VPWR.t4335 4.36035
R6226 VPWR.n1694 VPWR.t595 4.36035
R6227 VPWR.n1692 VPWR.t5516 4.36035
R6228 VPWR.n1690 VPWR.t4044 4.36035
R6229 VPWR.n1688 VPWR.t4080 4.36035
R6230 VPWR.n1685 VPWR.t5508 4.36035
R6231 VPWR.n768 VPWR.t491 4.36035
R6232 VPWR.n768 VPWR.t6149 4.36035
R6233 VPWR.n767 VPWR.t2684 4.36035
R6234 VPWR.n767 VPWR.t398 4.36035
R6235 VPWR.n766 VPWR.t1574 4.36035
R6236 VPWR.n766 VPWR.t6247 4.36035
R6237 VPWR.n765 VPWR.t929 4.36035
R6238 VPWR.n765 VPWR.t2304 4.36035
R6239 VPWR.n3238 VPWR.t3647 4.36035
R6240 VPWR.n3247 VPWR.t1883 4.36035
R6241 VPWR.n3246 VPWR.t362 4.36035
R6242 VPWR.n3246 VPWR.t3335 4.36035
R6243 VPWR.n122 VPWR.t4995 4.36035
R6244 VPWR.n122 VPWR.t5779 4.36035
R6245 VPWR.n3298 VPWR.t3629 4.36035
R6246 VPWR.n3296 VPWR.t2796 4.36035
R6247 VPWR.n3294 VPWR.t343 4.36035
R6248 VPWR.n3275 VPWR.t3514 4.36035
R6249 VPWR.n3275 VPWR.t2467 4.36035
R6250 VPWR.n3274 VPWR.t5680 4.36035
R6251 VPWR.n3274 VPWR.t1937 4.36035
R6252 VPWR.n3276 VPWR.t5215 4.36035
R6253 VPWR.n3278 VPWR.t2418 4.36035
R6254 VPWR.n3280 VPWR.t2623 4.36035
R6255 VPWR.n3281 VPWR.t2232 4.36035
R6256 VPWR.n3283 VPWR.t2175 4.36035
R6257 VPWR.n3284 VPWR.t4903 4.36035
R6258 VPWR.n3288 VPWR.t6261 4.36035
R6259 VPWR.n3290 VPWR.t5238 4.36035
R6260 VPWR.n3293 VPWR.t3193 4.36035
R6261 VPWR.n3305 VPWR.t6095 4.36035
R6262 VPWR.n3306 VPWR.t5217 4.36035
R6263 VPWR.n3309 VPWR.t2420 4.36035
R6264 VPWR.n3236 VPWR.t3493 4.36035
R6265 VPWR.n3235 VPWR.t6259 4.36035
R6266 VPWR.n762 VPWR.t3358 4.36035
R6267 VPWR.n764 VPWR.t2092 4.36035
R6268 VPWR.n769 VPWR.t3171 4.36035
R6269 VPWR.n773 VPWR.t3971 4.36035
R6270 VPWR.n775 VPWR.t4149 4.36035
R6271 VPWR.n776 VPWR.t7118 4.36035
R6272 VPWR.n778 VPWR.t6032 4.36035
R6273 VPWR.n779 VPWR.t3684 4.36035
R6274 VPWR.n781 VPWR.t5093 4.36035
R6275 VPWR.n1691 VPWR.t4568 4.36035
R6276 VPWR.n1230 VPWR.t923 4.36035
R6277 VPWR.n1232 VPWR.t2589 4.36035
R6278 VPWR.n1237 VPWR.t716 4.36035
R6279 VPWR.n1239 VPWR.t935 4.36035
R6280 VPWR.n1241 VPWR.t3907 4.36035
R6281 VPWR.n1243 VPWR.t5029 4.36035
R6282 VPWR.n1245 VPWR.t1235 4.36035
R6283 VPWR.n1258 VPWR.t706 4.36035
R6284 VPWR.n1262 VPWR.t4235 4.36035
R6285 VPWR.n1178 VPWR.t684 4.36035
R6286 VPWR.n1712 VPWR.t445 4.36035
R6287 VPWR.n1722 VPWR.t5097 4.36035
R6288 VPWR.n1722 VPWR.t4538 4.36035
R6289 VPWR.n1723 VPWR.t1610 4.36035
R6290 VPWR.n1723 VPWR.t2920 4.36035
R6291 VPWR.n1724 VPWR.t1144 4.36035
R6292 VPWR.n1724 VPWR.t2163 4.36035
R6293 VPWR.n1725 VPWR.t1442 4.36035
R6294 VPWR.n1725 VPWR.t3256 4.36035
R6295 VPWR.n1726 VPWR.t6128 4.36035
R6296 VPWR.n1726 VPWR.t503 4.36035
R6297 VPWR.n1759 VPWR.t2919 4.36035
R6298 VPWR.n1797 VPWR.t1791 4.36035
R6299 VPWR.n1795 VPWR.t3238 4.36035
R6300 VPWR.n1794 VPWR.t6221 4.36035
R6301 VPWR.n1792 VPWR.t1538 4.36035
R6302 VPWR.n1791 VPWR.t4877 4.36035
R6303 VPWR.n3210 VPWR.t1636 4.36035
R6304 VPWR.n3207 VPWR.t355 4.36035
R6305 VPWR.n3179 VPWR.t4053 4.36035
R6306 VPWR.n3177 VPWR.t2246 4.36035
R6307 VPWR.n3174 VPWR.t5499 4.36035
R6308 VPWR.n3172 VPWR.t5434 4.36035
R6309 VPWR.n3170 VPWR.t1414 4.36035
R6310 VPWR.n3168 VPWR.t5776 4.36035
R6311 VPWR.n3166 VPWR.t601 4.36035
R6312 VPWR.n3164 VPWR.t5282 4.36035
R6313 VPWR.n3162 VPWR.t4128 4.36035
R6314 VPWR.n168 VPWR.t6211 4.36035
R6315 VPWR.n166 VPWR.t2794 4.36035
R6316 VPWR.n164 VPWR.t5988 4.36035
R6317 VPWR.n164 VPWR.t2128 4.36035
R6318 VPWR.n163 VPWR.t6440 4.36035
R6319 VPWR.n163 VPWR.t1477 4.36035
R6320 VPWR.n162 VPWR.t6354 4.36035
R6321 VPWR.n162 VPWR.t5902 4.36035
R6322 VPWR.n161 VPWR.t1238 4.36035
R6323 VPWR.n161 VPWR.t2687 4.36035
R6324 VPWR.n160 VPWR.t3370 4.36035
R6325 VPWR.n160 VPWR.t3616 4.36035
R6326 VPWR.n159 VPWR.t2992 4.36035
R6327 VPWR.n159 VPWR.t4974 4.36035
R6328 VPWR.n158 VPWR.t5124 4.36035
R6329 VPWR.n158 VPWR.t667 4.36035
R6330 VPWR.n157 VPWR.t7089 4.36035
R6331 VPWR.n157 VPWR.t3601 4.36035
R6332 VPWR.n167 VPWR.t665 4.36035
R6333 VPWR.n169 VPWR.t4593 4.36035
R6334 VPWR.n3163 VPWR.t5532 4.36035
R6335 VPWR.n3165 VPWR.t2432 4.36035
R6336 VPWR.n3167 VPWR.t6459 4.36035
R6337 VPWR.n3169 VPWR.t1594 4.36035
R6338 VPWR.n3171 VPWR.t3946 4.36035
R6339 VPWR.n3173 VPWR.t2615 4.36035
R6340 VPWR.n3176 VPWR.t3203 4.36035
R6341 VPWR.n3178 VPWR.t2416 4.36035
R6342 VPWR.n3180 VPWR.t4715 4.36035
R6343 VPWR.n3181 VPWR.t1996 4.36035
R6344 VPWR.n3184 VPWR.t6364 4.36035
R6345 VPWR.n3185 VPWR.t2802 4.36035
R6346 VPWR.n3187 VPWR.t4331 4.36035
R6347 VPWR.n3188 VPWR.t1384 4.36035
R6348 VPWR.n3189 VPWR.t1994 4.36035
R6349 VPWR.n3199 VPWR.t372 4.36035
R6350 VPWR.n3215 VPWR.t4041 4.36035
R6351 VPWR.n3217 VPWR.t4748 4.36035
R6352 VPWR.n3219 VPWR.t4709 4.36035
R6353 VPWR.n1787 VPWR.t2619 4.36035
R6354 VPWR.n1809 VPWR.t1786 4.36035
R6355 VPWR.n1727 VPWR.t5405 4.36035
R6356 VPWR.n1721 VPWR.t5071 4.36035
R6357 VPWR.n1170 VPWR.t5186 4.36035
R6358 VPWR.n1154 VPWR.t761 4.36035
R6359 VPWR.n1153 VPWR.t1536 4.36035
R6360 VPWR.n1152 VPWR.t63 4.36035
R6361 VPWR.n1152 VPWR.t4971 4.36035
R6362 VPWR.n1151 VPWR.t4844 4.36035
R6363 VPWR.n1151 VPWR.t4410 4.36035
R6364 VPWR.n1150 VPWR.t1037 4.36035
R6365 VPWR.n1150 VPWR.t3969 4.36035
R6366 VPWR.n1149 VPWR.t5292 4.36035
R6367 VPWR.n1149 VPWR.t6138 4.36035
R6368 VPWR.n1148 VPWR.t3798 4.36035
R6369 VPWR.n1145 VPWR.t1400 4.36035
R6370 VPWR.n1143 VPWR.t2753 4.36035
R6371 VPWR.n1132 VPWR.t2498 4.36035
R6372 VPWR.n1132 VPWR.t2843 4.36035
R6373 VPWR.n1123 VPWR.t1223 4.36035
R6374 VPWR.n1121 VPWR.t5025 4.36035
R6375 VPWR.n1119 VPWR.t5801 4.36035
R6376 VPWR.n1117 VPWR.t3388 4.36035
R6377 VPWR.n1115 VPWR.t2177 4.36035
R6378 VPWR.n1113 VPWR.t2534 4.36035
R6379 VPWR.n1111 VPWR.t2108 4.36035
R6380 VPWR.n1110 VPWR.t554 4.36035
R6381 VPWR.n679 VPWR.t3591 4.36035
R6382 VPWR.n678 VPWR.t5366 4.36035
R6383 VPWR.n675 VPWR.t1454 4.36035
R6384 VPWR.n674 VPWR.t5192 4.36035
R6385 VPWR.n658 VPWR.t718 4.36035
R6386 VPWR.n656 VPWR.t704 4.36035
R6387 VPWR.n654 VPWR.t2948 4.36035
R6388 VPWR.n652 VPWR.t4955 4.36035
R6389 VPWR.n650 VPWR.t4985 4.36035
R6390 VPWR.n647 VPWR.t4889 4.36035
R6391 VPWR.n641 VPWR.t1554 4.36035
R6392 VPWR.n639 VPWR.t571 4.36035
R6393 VPWR.n637 VPWR.t1160 4.36035
R6394 VPWR.n172 VPWR.t4098 4.36035
R6395 VPWR.n3111 VPWR.t2679 4.36035
R6396 VPWR.n3113 VPWR.t3272 4.36035
R6397 VPWR.n3116 VPWR.t449 4.36035
R6398 VPWR.n3118 VPWR.t5300 4.36035
R6399 VPWR.n3120 VPWR.t3645 4.36035
R6400 VPWR.n3122 VPWR.t5637 4.36035
R6401 VPWR.n3124 VPWR.t4486 4.36035
R6402 VPWR.n3126 VPWR.t331 4.36035
R6403 VPWR.n3128 VPWR.t5781 4.36035
R6404 VPWR.n3130 VPWR.t5332 4.36035
R6405 VPWR.n3143 VPWR.t2532 4.36035
R6406 VPWR.n3141 VPWR.t1756 4.36035
R6407 VPWR.n3139 VPWR.t722 4.36035
R6408 VPWR.n3137 VPWR.t710 4.36035
R6409 VPWR.n3135 VPWR.t1506 4.36035
R6410 VPWR.n3133 VPWR.t1828 4.36035
R6411 VPWR.n171 VPWR.t4944 4.36035
R6412 VPWR.n3156 VPWR.t2098 4.36035
R6413 VPWR.n3154 VPWR.t5834 4.36035
R6414 VPWR.n3152 VPWR.t4591 4.36035
R6415 VPWR.n3152 VPWR.t2492 4.36035
R6416 VPWR.n3151 VPWR.t2965 4.36035
R6417 VPWR.n3151 VPWR.t1902 4.36035
R6418 VPWR.n3150 VPWR.t2836 4.36035
R6419 VPWR.n3150 VPWR.t416 4.36035
R6420 VPWR.n3149 VPWR.t1644 4.36035
R6421 VPWR.n3149 VPWR.t4631 4.36035
R6422 VPWR.n3148 VPWR.t2422 4.36035
R6423 VPWR.n3148 VPWR.t732 4.36035
R6424 VPWR.n3147 VPWR.t5220 4.36035
R6425 VPWR.n3147 VPWR.t1736 4.36035
R6426 VPWR.n3146 VPWR.t3813 4.36035
R6427 VPWR.n3146 VPWR.t3804 4.36035
R6428 VPWR.n3145 VPWR.t5984 4.36035
R6429 VPWR.n3145 VPWR.t1973 4.36035
R6430 VPWR.n3155 VPWR.t5265 4.36035
R6431 VPWR.n3157 VPWR.t1606 4.36035
R6432 VPWR.n3132 VPWR.t3922 4.36035
R6433 VPWR.n3134 VPWR.t702 4.36035
R6434 VPWR.n3136 VPWR.t1961 4.36035
R6435 VPWR.n3138 VPWR.t1396 4.36035
R6436 VPWR.n3140 VPWR.t5415 4.36035
R6437 VPWR.n3142 VPWR.t3997 4.36035
R6438 VPWR.n3131 VPWR.t5100 4.36035
R6439 VPWR.n3129 VPWR.t4059 4.36035
R6440 VPWR.n3127 VPWR.t3500 4.36035
R6441 VPWR.n3125 VPWR.t2386 4.36035
R6442 VPWR.n3123 VPWR.t1852 4.36035
R6443 VPWR.n3121 VPWR.t4392 4.36035
R6444 VPWR.n3119 VPWR.t6350 4.36035
R6445 VPWR.n3117 VPWR.t6242 4.36035
R6446 VPWR.n3115 VPWR.t5575 4.36035
R6447 VPWR.n3112 VPWR.t5381 4.36035
R6448 VPWR.n3110 VPWR.t1386 4.36035
R6449 VPWR.n636 VPWR.t824 4.36035
R6450 VPWR.n638 VPWR.t6269 4.36035
R6451 VPWR.n640 VPWR.t1713 4.36035
R6452 VPWR.n643 VPWR.t5758 4.36035
R6453 VPWR.n645 VPWR.t4528 4.36035
R6454 VPWR.n646 VPWR.t4442 4.36035
R6455 VPWR.n649 VPWR.t4341 4.36035
R6456 VPWR.n651 VPWR.t4936 4.36035
R6457 VPWR.n653 VPWR.t994 4.36035
R6458 VPWR.n655 VPWR.t5862 4.36035
R6459 VPWR.n657 VPWR.t2480 4.36035
R6460 VPWR.n659 VPWR.t1951 4.36035
R6461 VPWR.n660 VPWR.t583 4.36035
R6462 VPWR.n662 VPWR.t4668 4.36035
R6463 VPWR.n664 VPWR.t3092 4.36035
R6464 VPWR.n676 VPWR.t1664 4.36035
R6465 VPWR.n1838 VPWR.t1 4.36035
R6466 VPWR.n1116 VPWR.t515 4.36035
R6467 VPWR.n1118 VPWR.t876 4.36035
R6468 VPWR.n1120 VPWR.t3676 4.36035
R6469 VPWR.n1133 VPWR.t5111 4.36035
R6470 VPWR.n1140 VPWR.t765 4.36035
R6471 VPWR.n1142 VPWR.t5152 4.36035
R6472 VPWR.n1144 VPWR.t3042 4.36035
R6473 VPWR.n1147 VPWR.t2779 4.36035
R6474 VPWR.n1155 VPWR.t3496 4.36035
R6475 VPWR.n1935 VPWR.t3851 4.36035
R6476 VPWR.n1933 VPWR.t1261 4.36035
R6477 VPWR.n1931 VPWR.t1675 4.36035
R6478 VPWR.n1929 VPWR.t632 4.36035
R6479 VPWR.n1927 VPWR.t2090 4.36035
R6480 VPWR.n2003 VPWR.t6078 4.36035
R6481 VPWR.n2001 VPWR.t5325 4.36035
R6482 VPWR.n2001 VPWR.t3057 4.36035
R6483 VPWR.n2000 VPWR.t2248 4.36035
R6484 VPWR.n2000 VPWR.t6161 4.36035
R6485 VPWR.n1999 VPWR.t1722 4.36035
R6486 VPWR.n1999 VPWR.t3051 4.36035
R6487 VPWR.n1998 VPWR.t5106 4.36035
R6488 VPWR.n1998 VPWR.t59 4.36035
R6489 VPWR.n1997 VPWR.t1990 4.36035
R6490 VPWR.n1997 VPWR.t4299 4.36035
R6491 VPWR.n1996 VPWR.t4067 4.36035
R6492 VPWR.n1996 VPWR.t4863 4.36035
R6493 VPWR.n1995 VPWR.t3860 4.36035
R6494 VPWR.n1995 VPWR.t5448 4.36035
R6495 VPWR.n1994 VPWR.t6452 4.36035
R6496 VPWR.n1994 VPWR.t4622 4.36035
R6497 VPWR.n1978 VPWR.t2767 4.36035
R6498 VPWR.n1976 VPWR.t1628 4.36035
R6499 VPWR.n1973 VPWR.t5845 4.36035
R6500 VPWR.n1971 VPWR.t4927 4.36035
R6501 VPWR.n1971 VPWR.t6074 4.36035
R6502 VPWR.n1957 VPWR.t2071 4.36035
R6503 VPWR.n1955 VPWR.t2852 4.36035
R6504 VPWR.n1951 VPWR.t4428 4.36035
R6505 VPWR.n2839 VPWR.t5559 4.36035
R6506 VPWR.n2841 VPWR.t4740 4.36035
R6507 VPWR.n2859 VPWR.t4790 4.36035
R6508 VPWR.n2859 VPWR.t2516 4.36035
R6509 VPWR.n2889 VPWR.t4046 4.36035
R6510 VPWR.n2888 VPWR.t5778 4.36035
R6511 VPWR.n2888 VPWR.t2942 4.36035
R6512 VPWR.n2887 VPWR.t2792 4.36035
R6513 VPWR.n2887 VPWR.t3733 4.36035
R6514 VPWR.n2886 VPWR.t7088 4.36035
R6515 VPWR.n2886 VPWR.t4713 4.36035
R6516 VPWR.n2885 VPWR.t1254 4.36035
R6517 VPWR.n2885 VPWR.t5579 4.36035
R6518 VPWR.n2884 VPWR.t4444 4.36035
R6519 VPWR.n2884 VPWR.t5354 4.36035
R6520 VPWR.n2883 VPWR.t5871 4.36035
R6521 VPWR.n2883 VPWR.t3512 4.36035
R6522 VPWR.n2882 VPWR.t2964 4.36035
R6523 VPWR.n2882 VPWR.t5744 4.36035
R6524 VPWR.n2881 VPWR.t1471 4.36035
R6525 VPWR.n2881 VPWR.t1082 4.36035
R6526 VPWR.n2890 VPWR.t563 4.36035
R6527 VPWR.n2893 VPWR.t4303 4.36035
R6528 VPWR.n2895 VPWR.t5277 4.36035
R6529 VPWR.n2896 VPWR.t686 4.36035
R6530 VPWR.n2898 VPWR.t2343 4.36035
R6531 VPWR.n2846 VPWR.t1311 4.36035
R6532 VPWR.n2845 VPWR.t978 4.36035
R6533 VPWR.n2844 VPWR.t5184 4.36035
R6534 VPWR.n2842 VPWR.t4957 4.36035
R6535 VPWR.n2840 VPWR.t2854 4.36035
R6536 VPWR.n2838 VPWR.t6454 4.36035
R6537 VPWR.n2836 VPWR.t364 4.36035
R6538 VPWR.n2833 VPWR.t3543 4.36035
R6539 VPWR.n1940 VPWR.t787 4.36035
R6540 VPWR.n1941 VPWR.t2994 4.36035
R6541 VPWR.n1943 VPWR.t4265 4.36035
R6542 VPWR.n1945 VPWR.t5512 4.36035
R6543 VPWR.n1947 VPWR.t2635 4.36035
R6544 VPWR.n1948 VPWR.t1281 4.36035
R6545 VPWR.n1950 VPWR.t1793 4.36035
R6546 VPWR.n1952 VPWR.t3625 4.36035
R6547 VPWR.n1954 VPWR.t2020 4.36035
R6548 VPWR.n1956 VPWR.t4646 4.36035
R6549 VPWR.n1958 VPWR.t5421 4.36035
R6550 VPWR.n1968 VPWR.t6328 4.36035
R6551 VPWR.n1970 VPWR.t5324 4.36035
R6552 VPWR.n1975 VPWR.t1193 4.36035
R6553 VPWR.n1993 VPWR.t5966 4.36035
R6554 VPWR.n1926 VPWR.t4065 4.36035
R6555 VPWR.n1928 VPWR.t1986 4.36035
R6556 VPWR.n1930 VPWR.t2536 4.36035
R6557 VPWR.n1932 VPWR.t1718 4.36035
R6558 VPWR.n1934 VPWR.t1673 4.36035
R6559 VPWR.n350 VPWR.t4196 4.36035
R6560 VPWR.n352 VPWR.t2143 4.36035
R6561 VPWR.n354 VPWR.t605 4.36035
R6562 VPWR.n356 VPWR.t1172 4.36035
R6563 VPWR.n358 VPWR.t1774 4.36035
R6564 VPWR.n2103 VPWR.t3516 4.36035
R6565 VPWR.n2105 VPWR.t5679 4.36035
R6566 VPWR.n2107 VPWR.t5769 4.36035
R6567 VPWR.n2110 VPWR.t4311 4.36035
R6568 VPWR.n2112 VPWR.t2518 4.36035
R6569 VPWR.n2114 VPWR.t2320 4.36035
R6570 VPWR.n2116 VPWR.t5700 4.36035
R6571 VPWR.n2118 VPWR.t6001 4.36035
R6572 VPWR.n2120 VPWR.t2010 4.36035
R6573 VPWR.n2122 VPWR.t4540 4.36035
R6574 VPWR.n2124 VPWR.t2219 4.36035
R6575 VPWR.n2127 VPWR.t591 4.36035
R6576 VPWR.n2127 VPWR.t3609 4.36035
R6577 VPWR.n2128 VPWR.t4770 4.36035
R6578 VPWR.n2128 VPWR.t3788 4.36035
R6579 VPWR.n2129 VPWR.t4308 4.36035
R6580 VPWR.n2129 VPWR.t5045 4.36035
R6581 VPWR.n2130 VPWR.t1782 4.36035
R6582 VPWR.n2130 VPWR.t5241 4.36035
R6583 VPWR.n2131 VPWR.t6039 4.36035
R6584 VPWR.n2135 VPWR.t4019 4.36035
R6585 VPWR.n2137 VPWR.t2145 4.36035
R6586 VPWR.n2139 VPWR.t497 4.36035
R6587 VPWR.n2142 VPWR.t5979 4.36035
R6588 VPWR.n2144 VPWR.t3226 4.36035
R6589 VPWR.n2146 VPWR.t4919 4.36035
R6590 VPWR.n2148 VPWR.t459 4.36035
R6591 VPWR.n2150 VPWR.t5771 4.36035
R6592 VPWR.n2152 VPWR.t4163 4.36035
R6593 VPWR.n2154 VPWR.t1845 4.36035
R6594 VPWR.n2156 VPWR.t3929 4.36035
R6595 VPWR.n2166 VPWR.t495 4.36035
R6596 VPWR.n2164 VPWR.t3608 4.36035
R6597 VPWR.n2162 VPWR.t5710 4.36035
R6598 VPWR.n2160 VPWR.t4239 4.36035
R6599 VPWR.n2158 VPWR.t3187 4.36035
R6600 VPWR.n2183 VPWR.t4546 4.36035
R6601 VPWR.n2181 VPWR.t5725 4.36035
R6602 VPWR.n2179 VPWR.t6160 4.36035
R6603 VPWR.n2177 VPWR.t3618 4.36035
R6604 VPWR.n2175 VPWR.t1225 4.36035
R6605 VPWR.n2175 VPWR.t4716 4.36035
R6606 VPWR.n2174 VPWR.t3567 4.36035
R6607 VPWR.n2174 VPWR.t4033 4.36035
R6608 VPWR.n2173 VPWR.t2713 4.36035
R6609 VPWR.n2173 VPWR.t1045 4.36035
R6610 VPWR.n2172 VPWR.t976 4.36035
R6611 VPWR.n2172 VPWR.t5341 4.36035
R6612 VPWR.n2171 VPWR.t349 4.36035
R6613 VPWR.n2171 VPWR.t1837 4.36035
R6614 VPWR.n2170 VPWR.t394 4.36035
R6615 VPWR.n2170 VPWR.t2461 4.36035
R6616 VPWR.n2169 VPWR.t3205 4.36035
R6617 VPWR.n2169 VPWR.t3227 4.36035
R6618 VPWR.n2168 VPWR.t5135 4.36035
R6619 VPWR.n2168 VPWR.t3038 4.36035
R6620 VPWR.n2178 VPWR.t4396 4.36035
R6621 VPWR.n2180 VPWR.t1475 4.36035
R6622 VPWR.n2182 VPWR.t682 4.36035
R6623 VPWR.n348 VPWR.t4354 4.36035
R6624 VPWR.n2159 VPWR.t3547 4.36035
R6625 VPWR.n2161 VPWR.t6283 4.36035
R6626 VPWR.n2163 VPWR.t2662 4.36035
R6627 VPWR.n2165 VPWR.t1550 4.36035
R6628 VPWR.n2157 VPWR.t428 4.36035
R6629 VPWR.n2155 VPWR.t3263 4.36035
R6630 VPWR.n2153 VPWR.t4032 4.36035
R6631 VPWR.n2151 VPWR.t3247 4.36035
R6632 VPWR.n2149 VPWR.t4362 4.36035
R6633 VPWR.n2147 VPWR.t1279 4.36035
R6634 VPWR.n2145 VPWR.t1450 4.36035
R6635 VPWR.n2143 VPWR.t2270 4.36035
R6636 VPWR.n2141 VPWR.t2715 4.36035
R6637 VPWR.n2138 VPWR.t3232 4.36035
R6638 VPWR.n2136 VPWR.t5822 4.36035
R6639 VPWR.n2133 VPWR.t1072 4.36035
R6640 VPWR.n2125 VPWR.t6180 4.36035
R6641 VPWR.n2123 VPWR.t4970 4.36035
R6642 VPWR.n2121 VPWR.t1134 4.36035
R6643 VPWR.n2119 VPWR.t757 4.36035
R6644 VPWR.n2117 VPWR.t6194 4.36035
R6645 VPWR.n2115 VPWR.t2430 4.36035
R6646 VPWR.n2113 VPWR.t4368 4.36035
R6647 VPWR.n2111 VPWR.t4848 4.36035
R6648 VPWR.n2109 VPWR.t724 4.36035
R6649 VPWR.n2106 VPWR.t3185 4.36035
R6650 VPWR.n2104 VPWR.t2757 4.36035
R6651 VPWR.n2102 VPWR.t4358 4.36035
R6652 VPWR.n357 VPWR.t1277 4.36035
R6653 VPWR.n355 VPWR.t1448 4.36035
R6654 VPWR.n353 VPWR.t4907 4.36035
R6655 VPWR.n351 VPWR.t1880 4.36035
R6656 VPWR.n349 VPWR.t5163 4.36035
R6657 VPWR.n287 VPWR.t1646 4.36035
R6658 VPWR.n289 VPWR.t1707 4.36035
R6659 VPWR.n291 VPWR.t1229 4.36035
R6660 VPWR.n293 VPWR.t5037 4.36035
R6661 VPWR.n295 VPWR.t4759 4.36035
R6662 VPWR.n298 VPWR.t2201 4.36035
R6663 VPWR.n300 VPWR.t4767 4.36035
R6664 VPWR.n302 VPWR.t3191 4.36035
R6665 VPWR.n305 VPWR.t4447 4.36035
R6666 VPWR.n307 VPWR.t3816 4.36035
R6667 VPWR.n309 VPWR.t2472 4.36035
R6668 VPWR.n311 VPWR.t2494 4.36035
R6669 VPWR.n313 VPWR.t5453 4.36035
R6670 VPWR.n315 VPWR.t3887 4.36035
R6671 VPWR.n317 VPWR.t4815 4.36035
R6672 VPWR.n319 VPWR.t4654 4.36035
R6673 VPWR.n330 VPWR.t1766 4.36035
R6674 VPWR.n328 VPWR.t4298 4.36035
R6675 VPWR.n326 VPWR.t4862 4.36035
R6676 VPWR.n324 VPWR.t4707 4.36035
R6677 VPWR.n322 VPWR.t2213 4.36035
R6678 VPWR.n285 VPWR.t745 4.36035
R6679 VPWR.n2273 VPWR.t6110 4.36035
R6680 VPWR.n2271 VPWR.t5061 4.36035
R6681 VPWR.n2269 VPWR.t3627 4.36035
R6682 VPWR.n2266 VPWR.t4513 4.36035
R6683 VPWR.n2264 VPWR.t3597 4.36035
R6684 VPWR.n2262 VPWR.t4590 4.36035
R6685 VPWR.n2260 VPWR.t4455 4.36035
R6686 VPWR.n2258 VPWR.t6209 4.36035
R6687 VPWR.n2256 VPWR.t3808 4.36035
R6688 VPWR.n2254 VPWR.t4025 4.36035
R6689 VPWR.n2252 VPWR.t1466 4.36035
R6690 VPWR.n2249 VPWR.t3818 4.36035
R6691 VPWR.n2247 VPWR.t489 4.36035
R6692 VPWR.n2245 VPWR.t2627 4.36035
R6693 VPWR.n2243 VPWR.t6192 4.36035
R6694 VPWR.n2241 VPWR.t4491 4.36035
R6695 VPWR.n347 VPWR.t4615 4.36035
R6696 VPWR.n345 VPWR.t4152 4.36035
R6697 VPWR.n343 VPWR.t1854 4.36035
R6698 VPWR.n341 VPWR.t1562 4.36035
R6699 VPWR.n339 VPWR.t1914 4.36035
R6700 VPWR.n339 VPWR.t581 4.36035
R6701 VPWR.n338 VPWR.t5451 4.36035
R6702 VPWR.n338 VPWR.t4101 4.36035
R6703 VPWR.n337 VPWR.t1392 4.36035
R6704 VPWR.n337 VPWR.t3109 4.36035
R6705 VPWR.n336 VPWR.t3079 4.36035
R6706 VPWR.n336 VPWR.t1336 4.36035
R6707 VPWR.n335 VPWR.t6326 4.36035
R6708 VPWR.n335 VPWR.t2528 4.36035
R6709 VPWR.n334 VPWR.t3386 4.36035
R6710 VPWR.n334 VPWR.t4575 4.36035
R6711 VPWR.n333 VPWR.t5742 4.36035
R6712 VPWR.n333 VPWR.t3981 4.36035
R6713 VPWR.n332 VPWR.t3903 4.36035
R6714 VPWR.n332 VPWR.t5647 4.36035
R6715 VPWR.n342 VPWR.t2842 4.36035
R6716 VPWR.n344 VPWR.t5273 4.36035
R6717 VPWR.n346 VPWR.t3169 4.36035
R6718 VPWR.n2240 VPWR.t6054 4.36035
R6719 VPWR.n2242 VPWR.t3354 4.36035
R6720 VPWR.n2244 VPWR.t4875 4.36035
R6721 VPWR.n2246 VPWR.t676 4.36035
R6722 VPWR.n2248 VPWR.t4915 4.36035
R6723 VPWR.n2251 VPWR.t4526 4.36035
R6724 VPWR.n2253 VPWR.t1655 4.36035
R6725 VPWR.n2255 VPWR.t3726 4.36035
R6726 VPWR.n2257 VPWR.t61 4.36035
R6727 VPWR.n2259 VPWR.t6219 4.36035
R6728 VPWR.n2261 VPWR.t4352 4.36035
R6729 VPWR.n2263 VPWR.t5631 4.36035
R6730 VPWR.n2265 VPWR.t6089 4.36035
R6731 VPWR.n2267 VPWR.t4009 4.36035
R6732 VPWR.n2270 VPWR.t3545 4.36035
R6733 VPWR.n2272 VPWR.t3214 4.36035
R6734 VPWR.n2274 VPWR.t3589 4.36035
R6735 VPWR.n321 VPWR.t1422 4.36035
R6736 VPWR.n323 VPWR.t2057 4.36035
R6737 VPWR.n325 VPWR.t5482 4.36035
R6738 VPWR.n327 VPWR.t6151 4.36035
R6739 VPWR.n329 VPWR.t5173 4.36035
R6740 VPWR.n320 VPWR.t5542 4.36035
R6741 VPWR.n318 VPWR.t4254 4.36035
R6742 VPWR.n316 VPWR.t945 4.36035
R6743 VPWR.n314 VPWR.t4941 4.36035
R6744 VPWR.n312 VPWR.t3365 4.36035
R6745 VPWR.n310 VPWR.t3775 4.36035
R6746 VPWR.n308 VPWR.t783 4.36035
R6747 VPWR.n306 VPWR.t3854 4.36035
R6748 VPWR.n304 VPWR.t3094 4.36035
R6749 VPWR.n301 VPWR.t5852 4.36035
R6750 VPWR.n299 VPWR.t1090 4.36035
R6751 VPWR.n297 VPWR.t2889 4.36035
R6752 VPWR.n294 VPWR.t5841 4.36035
R6753 VPWR.n292 VPWR.t1008 4.36035
R6754 VPWR.n290 VPWR.t2133 4.36035
R6755 VPWR.n288 VPWR.t4190 4.36035
R6756 VPWR.n286 VPWR.t3318 4.36035
R6757 VPWR.n2385 VPWR.t6202 4.36035
R6758 VPWR.n2388 VPWR.t1402 4.36035
R6759 VPWR.n2388 VPWR.t3234 4.36035
R6760 VPWR.n2387 VPWR.t5677 4.36035
R6761 VPWR.n2387 VPWR.t5035 4.36035
R6762 VPWR.n2386 VPWR.t2732 4.36035
R6763 VPWR.n2386 VPWR.t4827 4.36035
R6764 VPWR.n2384 VPWR.t1616 4.36035
R6765 VPWR.n2384 VPWR.t4371 4.36035
R6766 VPWR.n2392 VPWR.t6441 4.36035
R6767 VPWR.n2392 VPWR.t5820 4.36035
R6768 VPWR.n2391 VPWR.t7114 4.36035
R6769 VPWR.n2391 VPWR.t3455 4.36035
R6770 VPWR.n2390 VPWR.t6238 4.36035
R6771 VPWR.n2390 VPWR.t3433 4.36035
R6772 VPWR.n2389 VPWR.t5837 4.36035
R6773 VPWR.n2389 VPWR.t2341 4.36035
R6774 VPWR.n2396 VPWR.t3524 4.36035
R6775 VPWR.n2399 VPWR.t4445 4.36035
R6776 VPWR.n2399 VPWR.t4214 4.36035
R6777 VPWR.n2398 VPWR.t3539 4.36035
R6778 VPWR.n2398 VPWR.t996 4.36035
R6779 VPWR.n2397 VPWR.t6020 4.36035
R6780 VPWR.n2397 VPWR.t5506 4.36035
R6781 VPWR.n2395 VPWR.t1209 4.36035
R6782 VPWR.n2395 VPWR.t6186 4.36035
R6783 VPWR.n2403 VPWR.t5182 4.36035
R6784 VPWR.n2403 VPWR.t3690 4.36035
R6785 VPWR.n2402 VPWR.t3513 4.36035
R6786 VPWR.n2402 VPWR.t3103 4.36035
R6787 VPWR.n2401 VPWR.t4757 4.36035
R6788 VPWR.n2401 VPWR.t2840 4.36035
R6789 VPWR.n2400 VPWR.t5307 4.36035
R6790 VPWR.n2400 VPWR.t6113 4.36035
R6791 VPWR.n2407 VPWR.t3643 4.36035
R6792 VPWR.n2410 VPWR.t3378 4.36035
R6793 VPWR.n2410 VPWR.t4741 4.36035
R6794 VPWR.n2409 VPWR.t6136 4.36035
R6795 VPWR.n2409 VPWR.t4055 4.36035
R6796 VPWR.n2408 VPWR.t3858 4.36035
R6797 VPWR.n2408 VPWR.t3437 4.36035
R6798 VPWR.n2406 VPWR.t2780 4.36035
R6799 VPWR.n2406 VPWR.t892 4.36035
R6800 VPWR.n2414 VPWR.t5993 4.36035
R6801 VPWR.n2414 VPWR.t998 4.36035
R6802 VPWR.n2413 VPWR.t678 4.36035
R6803 VPWR.n2413 VPWR.t3248 4.36035
R6804 VPWR.n2412 VPWR.t3117 4.36035
R6805 VPWR.n2412 VPWR.t6181 4.36035
R6806 VPWR.n2411 VPWR.t2496 4.36035
R6807 VPWR.n2411 VPWR.t2929 4.36035
R6808 VPWR.n282 VPWR.t3032 4.36035
R6809 VPWR.n280 VPWR.t6084 4.36035
R6810 VPWR.n278 VPWR.t1250 4.36035
R6811 VPWR.n276 VPWR.t473 4.36035
R6812 VPWR.n274 VPWR.t3452 4.36035
R6813 VPWR.n2313 VPWR.t3948 4.36035
R6814 VPWR.n2311 VPWR.t2061 4.36035
R6815 VPWR.n2309 VPWR.t2450 4.36035
R6816 VPWR.n2306 VPWR.t4857 4.36035
R6817 VPWR.n2304 VPWR.t493 4.36035
R6818 VPWR.n2302 VPWR.t3856 4.36035
R6819 VPWR.n2300 VPWR.t1195 4.36035
R6820 VPWR.n2298 VPWR.t1926 4.36035
R6821 VPWR.n2296 VPWR.t2193 4.36035
R6822 VPWR.n2294 VPWR.t4544 4.36035
R6823 VPWR.n2292 VPWR.t6056 4.36035
R6824 VPWR.n2289 VPWR.t1418 4.36035
R6825 VPWR.n2287 VPWR.t3177 4.36035
R6826 VPWR.n2285 VPWR.t3467 4.36035
R6827 VPWR.n2283 VPWR.t4807 4.36035
R6828 VPWR.n2281 VPWR.t5360 4.36035
R6829 VPWR.n2279 VPWR.t4595 4.36035
R6830 VPWR.n2187 VPWR.t3036 4.36035
R6831 VPWR.n2189 VPWR.t6086 4.36035
R6832 VPWR.n2191 VPWR.t1248 4.36035
R6833 VPWR.n2194 VPWR.t5995 4.36035
R6834 VPWR.n2196 VPWR.t3195 4.36035
R6835 VPWR.n2198 VPWR.t4921 4.36035
R6836 VPWR.n2200 VPWR.t680 4.36035
R6837 VPWR.n2202 VPWR.t2452 4.36035
R6838 VPWR.n2204 VPWR.t5944 4.36035
R6839 VPWR.n2206 VPWR.t534 4.36035
R6840 VPWR.n2208 VPWR.t3713 4.36035
R6841 VPWR.n2218 VPWR.t2474 4.36035
R6842 VPWR.n2216 VPWR.t2300 4.36035
R6843 VPWR.n2214 VPWR.t5606 4.36035
R6844 VPWR.n2212 VPWR.t1184 4.36035
R6845 VPWR.n2210 VPWR.t3444 4.36035
R6846 VPWR.n2235 VPWR.t4505 4.36035
R6847 VPWR.n2233 VPWR.t1287 4.36035
R6848 VPWR.n2231 VPWR.t1410 4.36035
R6849 VPWR.n2229 VPWR.t548 4.36035
R6850 VPWR.n2227 VPWR.t6127 4.36035
R6851 VPWR.n2227 VPWR.t4726 4.36035
R6852 VPWR.n2226 VPWR.t4170 4.36035
R6853 VPWR.n2226 VPWR.t5195 4.36035
R6854 VPWR.n2225 VPWR.t4878 4.36035
R6855 VPWR.n2225 VPWR.t1053 4.36035
R6856 VPWR.n2224 VPWR.t3382 4.36035
R6857 VPWR.n2224 VPWR.t4051 4.36035
R6858 VPWR.n2223 VPWR.t4129 4.36035
R6859 VPWR.n2223 VPWR.t1420 4.36035
R6860 VPWR.n2222 VPWR.t6450 4.36035
R6861 VPWR.n2222 VPWR.t2465 4.36035
R6862 VPWR.n2221 VPWR.t1227 4.36035
R6863 VPWR.n2221 VPWR.t3196 4.36035
R6864 VPWR.n2220 VPWR.t347 4.36035
R6865 VPWR.n2220 VPWR.t3363 4.36035
R6866 VPWR.n2230 VPWR.t6445 4.36035
R6867 VPWR.n2232 VPWR.t6308 4.36035
R6868 VPWR.n2234 VPWR.t73 4.36035
R6869 VPWR.n2186 VPWR.t1681 4.36035
R6870 VPWR.n2211 VPWR.t3674 4.36035
R6871 VPWR.n2213 VPWR.t5510 4.36035
R6872 VPWR.n2215 VPWR.t5450 4.36035
R6873 VPWR.n2217 VPWR.t3783 4.36035
R6874 VPWR.n2209 VPWR.t5556 4.36035
R6875 VPWR.n2207 VPWR.t3538 4.36035
R6876 VPWR.n2205 VPWR.t2018 4.36035
R6877 VPWR.n2203 VPWR.t4644 4.36035
R6878 VPWR.n2201 VPWR.t808 4.36035
R6879 VPWR.n2199 VPWR.t1275 4.36035
R6880 VPWR.n2197 VPWR.t1679 4.36035
R6881 VPWR.n2195 VPWR.t1760 4.36035
R6882 VPWR.n2193 VPWR.t5767 4.36035
R6883 VPWR.n2190 VPWR.t2096 4.36035
R6884 VPWR.n2188 VPWR.t2426 4.36035
R6885 VPWR.n284 VPWR.t2250 4.36035
R6886 VPWR.n2280 VPWR.t4637 4.36035
R6887 VPWR.n2282 VPWR.t4459 4.36035
R6888 VPWR.n2284 VPWR.t3334 4.36035
R6889 VPWR.n2286 VPWR.t7124 4.36035
R6890 VPWR.n2288 VPWR.t2798 4.36035
R6891 VPWR.n2291 VPWR.t5108 4.36035
R6892 VPWR.n2293 VPWR.t2408 4.36035
R6893 VPWR.n2295 VPWR.t2230 4.36035
R6894 VPWR.n2297 VPWR.t5956 4.36035
R6895 VPWR.n2299 VPWR.t4930 4.36035
R6896 VPWR.n2301 VPWR.t392 4.36035
R6897 VPWR.n2303 VPWR.t7086 4.36035
R6898 VPWR.n2305 VPWR.t7141 4.36035
R6899 VPWR.n2307 VPWR.t499 4.36035
R6900 VPWR.n2310 VPWR.t3050 4.36035
R6901 VPWR.n2312 VPWR.t4641 4.36035
R6902 VPWR.n2314 VPWR.t830 4.36035
R6903 VPWR.n275 VPWR.t3380 4.36035
R6904 VPWR.n277 VPWR.t5669 4.36035
R6905 VPWR.n279 VPWR.t2924 4.36035
R6906 VPWR.n281 VPWR.t1671 4.36035
R6907 VPWR.n283 VPWR.t3551 4.36035
R6908 VPWR.n2322 VPWR.t4304 4.36035
R6909 VPWR.n2322 VPWR.t4011 4.36035
R6910 VPWR.n2321 VPWR.t5098 4.36035
R6911 VPWR.n2321 VPWR.t1580 4.36035
R6912 VPWR.n2320 VPWR.t579 4.36035
R6913 VPWR.n2320 VPWR.t1896 4.36035
R6914 VPWR.n2317 VPWR.t884 4.36035
R6915 VPWR.n2317 VPWR.t5987 4.36035
R6916 VPWR.n2381 VPWR.t5181 4.36035
R6917 VPWR.n2381 VPWR.t990 4.36035
R6918 VPWR.n2380 VPWR.t4266 4.36035
R6919 VPWR.n2380 VPWR.t1343 4.36035
R6920 VPWR.n2379 VPWR.t4754 4.36035
R6921 VPWR.n2379 VPWR.t3968 4.36035
R6922 VPWR.n2378 VPWR.t5078 4.36035
R6923 VPWR.n2378 VPWR.t5646 4.36035
R6924 VPWR.n2376 VPWR.t692 4.36035
R6925 VPWR.n2375 VPWR.t2856 4.36035
R6926 VPWR.n2374 VPWR.t4407 4.36035
R6927 VPWR.n2373 VPWR.t1578 4.36035
R6928 VPWR.n2372 VPWR.t3794 4.36035
R6929 VPWR.n2371 VPWR.t5083 4.36035
R6930 VPWR.n2370 VPWR.t5581 4.36035
R6931 VPWR.n2369 VPWR.t5812 4.36035
R6932 VPWR.n2367 VPWR.t4377 4.36035
R6933 VPWR.n2366 VPWR.t552 4.36035
R6934 VPWR.n2365 VPWR.t1349 4.36035
R6935 VPWR.n2364 VPWR.t2088 4.36035
R6936 VPWR.n2363 VPWR.t4860 4.36035
R6937 VPWR.n2361 VPWR.t1546 4.36035
R6938 VPWR.n2360 VPWR.t447 4.36035
R6939 VPWR.n2359 VPWR.t3522 4.36035
R6940 VPWR.n2357 VPWR.t1094 4.36035
R6941 VPWR.n2356 VPWR.t4078 4.36035
R6942 VPWR.n2355 VPWR.t4976 4.36035
R6943 VPWR.n2354 VPWR.t5375 4.36035
R6944 VPWR.n2353 VPWR.t5787 4.36035
R6945 VPWR.n2352 VPWR.t6122 4.36035
R6946 VPWR.n2351 VPWR.t1498 4.36035
R6947 VPWR.n2350 VPWR.t3939 4.36035
R6948 VPWR.n2348 VPWR.t1939 4.36035
R6949 VPWR.n2347 VPWR.t5066 4.36035
R6950 VPWR.n2346 VPWR.t5649 4.36035
R6951 VPWR.n2345 VPWR.t1803 4.36035
R6952 VPWR.n2344 VPWR.t3294 4.36035
R6953 VPWR.n2342 VPWR.t6237 4.36035
R6954 VPWR.n2341 VPWR.t6273 4.36035
R6955 VPWR.n2340 VPWR.t4364 4.36035
R6956 VPWR.n2338 VPWR.t5715 4.36035
R6957 VPWR.n2337 VPWR.t2460 4.36035
R6958 VPWR.n2336 VPWR.t5839 4.36035
R6959 VPWR.n2335 VPWR.t5280 4.36035
R6960 VPWR.n2334 VPWR.t2693 4.36035
R6961 VPWR.n2333 VPWR.t6051 4.36035
R6962 VPWR.n2332 VPWR.t5286 4.36035
R6963 VPWR.n2331 VPWR.t1830 4.36035
R6964 VPWR.n2015 VPWR.t4934 4.36035
R6965 VPWR.n2013 VPWR.t2777 4.36035
R6966 VPWR.n2011 VPWR.t2075 4.36035
R6967 VPWR.n2009 VPWR.t5027 4.36035
R6968 VPWR.n2007 VPWR.t661 4.36035
R6969 VPWR.n2052 VPWR.t3392 4.36035
R6970 VPWR.n2049 VPWR.t4122 4.36035
R6971 VPWR.n2047 VPWR.t1856 4.36035
R6972 VPWR.n2045 VPWR.t1889 4.36035
R6973 VPWR.n2043 VPWR.t556 4.36035
R6974 VPWR.n2041 VPWR.t714 4.36035
R6975 VPWR.n2039 VPWR.t5756 4.36035
R6976 VPWR.n2037 VPWR.t5938 4.36035
R6977 VPWR.n2035 VPWR.t984 4.36035
R6978 VPWR.n2032 VPWR.t370 4.36035
R6979 VPWR.n2018 VPWR.t3770 4.36035
R6980 VPWR.n2016 VPWR.t4057 4.36035
R6981 VPWR.n2711 VPWR.t6312 4.36035
R6982 VPWR.n2713 VPWR.t3390 4.36035
R6983 VPWR.n2715 VPWR.t3796 4.36035
R6984 VPWR.n2717 VPWR.t2141 4.36035
R6985 VPWR.n2727 VPWR.t5312 4.36035
R6986 VPWR.n2745 VPWR.t2719 4.36035
R6987 VPWR.n2743 VPWR.t2173 4.36035
R6988 VPWR.n2741 VPWR.t565 4.36035
R6989 VPWR.n2739 VPWR.t741 4.36035
R6990 VPWR.n2737 VPWR.t6106 4.36035
R6991 VPWR.n2735 VPWR.t6018 4.36035
R6992 VPWR.n2733 VPWR.t1502 4.36035
R6993 VPWR.n2731 VPWR.t6325 4.36035
R6994 VPWR.n2827 VPWR.t4337 4.36035
R6995 VPWR.n2824 VPWR.t5960 4.36035
R6996 VPWR.n2822 VPWR.t5334 4.36035
R6997 VPWR.n2820 VPWR.t771 4.36035
R6998 VPWR.n2818 VPWR.t5538 4.36035
R6999 VPWR.n2816 VPWR.t3063 4.36035
R7000 VPWR.n2814 VPWR.t2833 4.36035
R7001 VPWR.n2812 VPWR.t6104 4.36035
R7002 VPWR.n2810 VPWR.t5428 4.36035
R7003 VPWR.n2807 VPWR.t1180 4.36035
R7004 VPWR.n2807 VPWR.t577 4.36035
R7005 VPWR.n2806 VPWR.t1979 4.36035
R7006 VPWR.n2806 VPWR.t5347 4.36035
R7007 VPWR.n2805 VPWR.t6348 4.36035
R7008 VPWR.n2805 VPWR.t3977 4.36035
R7009 VPWR.n2804 VPWR.t4476 4.36035
R7010 VPWR.n2804 VPWR.t327 4.36035
R7011 VPWR.n2784 VPWR.t4268 4.36035
R7012 VPWR.n2778 VPWR.t1556 4.36035
R7013 VPWR.n2776 VPWR.t573 4.36035
R7014 VPWR.n2774 VPWR.t2442 4.36035
R7015 VPWR.n2772 VPWR.t593 4.36035
R7016 VPWR.n2770 VPWR.t2147 4.36035
R7017 VPWR.n2768 VPWR.t1483 4.36035
R7018 VPWR.n2766 VPWR.t4572 4.36035
R7019 VPWR.n2764 VPWR.t5302 4.36035
R7020 VPWR.n2760 VPWR.t3394 4.36035
R7021 VPWR.n2758 VPWR.t652 4.36035
R7022 VPWR.n2758 VPWR.t5638 4.36035
R7023 VPWR.n2757 VPWR.t418 4.36035
R7024 VPWR.n2757 VPWR.t3668 4.36035
R7025 VPWR.n2756 VPWR.t3697 4.36035
R7026 VPWR.n2756 VPWR.t5038 4.36035
R7027 VPWR.n2755 VPWR.t4854 4.36035
R7028 VPWR.n2755 VPWR.t4765 4.36035
R7029 VPWR.n2754 VPWR.t4164 4.36035
R7030 VPWR.n2754 VPWR.t2906 4.36035
R7031 VPWR.n2753 VPWR.t1935 4.36035
R7032 VPWR.n2753 VPWR.t3994 4.36035
R7033 VPWR.n2752 VPWR.t767 4.36035
R7034 VPWR.n2752 VPWR.t2041 4.36035
R7035 VPWR.n2751 VPWR.t931 4.36035
R7036 VPWR.n2751 VPWR.t2305 4.36035
R7037 VPWR.n2761 VPWR.t3800 4.36035
R7038 VPWR.n2765 VPWR.t4120 4.36035
R7039 VPWR.n2767 VPWR.t816 4.36035
R7040 VPWR.n2769 VPWR.t2106 4.36035
R7041 VPWR.n2771 VPWR.t3715 4.36035
R7042 VPWR.n2773 VPWR.t2191 4.36035
R7043 VPWR.n2775 VPWR.t5760 4.36035
R7044 VPWR.n2777 VPWR.t4275 4.36035
R7045 VPWR.n2780 VPWR.t872 4.36035
R7046 VPWR.n2781 VPWR.t7116 4.36035
R7047 VPWR.n2783 VPWR.t5958 4.36035
R7048 VPWR.n2785 VPWR.t986 4.36035
R7049 VPWR.n2787 VPWR.t1504 4.36035
R7050 VPWR.n2790 VPWR.t2065 4.36035
R7051 VPWR.n2791 VPWR.t5748 4.36035
R7052 VPWR.n2792 VPWR.t3822 4.36035
R7053 VPWR.n2794 VPWR.t1564 4.36035
R7054 VPWR.n2798 VPWR.t1351 4.36035
R7055 VPWR.n2800 VPWR.t3012 4.36035
R7056 VPWR.n2802 VPWR.t2256 4.36035
R7057 VPWR.n2803 VPWR.t4577 4.36035
R7058 VPWR.n2809 VPWR.t2313 4.36035
R7059 VPWR.n2811 VPWR.t603 4.36035
R7060 VPWR.n2813 VPWR.t4519 4.36035
R7061 VPWR.n2815 VPWR.t7070 4.36035
R7062 VPWR.n2817 VPWR.t1642 4.36035
R7063 VPWR.n2819 VPWR.t1123 4.36035
R7064 VPWR.n2821 VPWR.t3954 4.36035
R7065 VPWR.n2823 VPWR.t3761 4.36035
R7066 VPWR.n2825 VPWR.t1060 4.36035
R7067 VPWR.n192 VPWR.t4574 4.36035
R7068 VPWR.n2732 VPWR.t5504 4.36035
R7069 VPWR.n2734 VPWR.t1885 4.36035
R7070 VPWR.n2736 VPWR.t2701 4.36035
R7071 VPWR.n2738 VPWR.t5904 4.36035
R7072 VPWR.n2740 VPWR.t3419 4.36035
R7073 VPWR.n2742 VPWR.t4664 4.36035
R7074 VPWR.n2744 VPWR.t7084 4.36035
R7075 VPWR.n2730 VPWR.t7132 4.36035
R7076 VPWR.n2728 VPWR.t5247 4.36035
R7077 VPWR.n2714 VPWR.t3763 4.36035
R7078 VPWR.n194 VPWR.t4769 4.36035
R7079 VPWR.n2017 VPWR.t7068 4.36035
R7080 VPWR.n2031 VPWR.t5294 4.36035
R7081 VPWR.n2034 VPWR.t5368 4.36035
R7082 VPWR.n2036 VPWR.t4846 4.36035
R7083 VPWR.n2038 VPWR.t313 4.36035
R7084 VPWR.n2040 VPWR.t870 4.36035
R7085 VPWR.n2042 VPWR.t2383 4.36035
R7086 VPWR.n2044 VPWR.t2157 4.36035
R7087 VPWR.n2046 VPWR.t2412 4.36035
R7088 VPWR.n2048 VPWR.t1345 4.36035
R7089 VPWR.n2050 VPWR.t1041 4.36035
R7090 VPWR.n2006 VPWR.t4017 4.36035
R7091 VPWR.n2008 VPWR.t3250 4.36035
R7092 VPWR.n2010 VPWR.t1816 4.36035
R7093 VPWR.n2012 VPWR.t6436 4.36035
R7094 VPWR.n2014 VPWR.t6457 4.36035
R7095 VPWR.n2064 VPWR.t5206 4.36035
R7096 VPWR.n2062 VPWR.t5900 4.36035
R7097 VPWR.n2060 VPWR.t619 4.36035
R7098 VPWR.n2058 VPWR.t3088 4.36035
R7099 VPWR.n2056 VPWR.t6231 4.36035
R7100 VPWR.n2097 VPWR.t410 4.36035
R7101 VPWR.n2095 VPWR.t1614 4.36035
R7102 VPWR.n2093 VPWR.t4626 4.36035
R7103 VPWR.n2091 VPWR.t1872 4.36035
R7104 VPWR.n2091 VPWR.t4378 4.36035
R7105 VPWR.n2090 VPWR.t5275 4.36035
R7106 VPWR.n2090 VPWR.t5878 4.36035
R7107 VPWR.n2089 VPWR.t1612 4.36035
R7108 VPWR.n2089 VPWR.t5259 4.36035
R7109 VPWR.n2088 VPWR.t4405 4.36035
R7110 VPWR.n2088 VPWR.t2677 4.36035
R7111 VPWR.n2087 VPWR.t5684 4.36035
R7112 VPWR.n2087 VPWR.t810 4.36035
R7113 VPWR.n2086 VPWR.t941 4.36035
R7114 VPWR.n2086 VPWR.t3814 4.36035
R7115 VPWR.n2083 VPWR.t2710 4.36035
R7116 VPWR.n2081 VPWR.t5850 4.36035
R7117 VPWR.n2691 VPWR.t5407 4.36035
R7118 VPWR.n2689 VPWR.t2763 4.36035
R7119 VPWR.n2687 VPWR.t4705 4.36035
R7120 VPWR.n2684 VPWR.t388 4.36035
R7121 VPWR.n2684 VPWR.t4736 4.36035
R7122 VPWR.n2683 VPWR.t4839 4.36035
R7123 VPWR.n2680 VPWR.t5892 4.36035
R7124 VPWR.n2678 VPWR.t1481 4.36035
R7125 VPWR.n2676 VPWR.t5729 4.36035
R7126 VPWR.n2674 VPWR.t812 4.36035
R7127 VPWR.n2672 VPWR.t4917 4.36035
R7128 VPWR.n2670 VPWR.t5150 4.36035
R7129 VPWR.n2667 VPWR.t3415 4.36035
R7130 VPWR.n2665 VPWR.t2996 4.36035
R7131 VPWR.n2663 VPWR.t3080 4.36035
R7132 VPWR.n2663 VPWR.t1807 4.36035
R7133 VPWR.n2662 VPWR.t4853 4.36035
R7134 VPWR.n2662 VPWR.t5554 4.36035
R7135 VPWR.n2661 VPWR.t4731 4.36035
R7136 VPWR.n2661 VPWR.t1632 4.36035
R7137 VPWR.n2660 VPWR.t2421 4.36035
R7138 VPWR.n2660 VPWR.t1510 4.36035
R7139 VPWR.n2659 VPWR.t5543 4.36035
R7140 VPWR.n2659 VPWR.t1560 4.36035
R7141 VPWR.n2658 VPWR.t4306 4.36035
R7142 VPWR.n2658 VPWR.t4942 4.36035
R7143 VPWR.n2657 VPWR.t67 4.36035
R7144 VPWR.n2657 VPWR.t4139 4.36035
R7145 VPWR.n2654 VPWR.t3657 4.36035
R7146 VPWR.n2652 VPWR.t4002 4.36035
R7147 VPWR.n2652 VPWR.t1148 4.36035
R7148 VPWR.n2651 VPWR.t5310 4.36035
R7149 VPWR.n2651 VPWR.t3641 4.36035
R7150 VPWR.n2650 VPWR.t1895 4.36035
R7151 VPWR.n2650 VPWR.t6135 4.36035
R7152 VPWR.n2649 VPWR.t3704 4.36035
R7153 VPWR.n2649 VPWR.t4356 4.36035
R7154 VPWR.n2648 VPWR.t700 4.36035
R7155 VPWR.n2648 VPWR.t2722 4.36035
R7156 VPWR.n2647 VPWR.t451 4.36035
R7157 VPWR.n2647 VPWR.t2220 4.36035
R7158 VPWR.n2646 VPWR.t5064 4.36035
R7159 VPWR.n2646 VPWR.t5031 4.36035
R7160 VPWR.n254 VPWR.t3648 4.36035
R7161 VPWR.n254 VPWR.t424 4.36035
R7162 VPWR.n253 VPWR.t2926 4.36035
R7163 VPWR.n250 VPWR.t4319 4.36035
R7164 VPWR.n248 VPWR.t2434 4.36035
R7165 VPWR.n246 VPWR.t3719 4.36035
R7166 VPWR.n244 VPWR.t2053 4.36035
R7167 VPWR.n242 VPWR.t2712 4.36035
R7168 VPWR.n240 VPWR.t2374 4.36035
R7169 VPWR.n238 VPWR.t2633 4.36035
R7170 VPWR.n235 VPWR.t3768 4.36035
R7171 VPWR.n232 VPWR.t1650 4.36035
R7172 VPWR.n230 VPWR.t3885 4.36035
R7173 VPWR.n228 VPWR.t5773 4.36035
R7174 VPWR.n226 VPWR.t1566 4.36035
R7175 VPWR.n224 VPWR.t5069 4.36035
R7176 VPWR.n222 VPWR.t5377 4.36035
R7177 VPWR.n220 VPWR.t1967 4.36035
R7178 VPWR.n217 VPWR.t5964 4.36035
R7179 VPWR.n215 VPWR.t3602 4.36035
R7180 VPWR.n215 VPWR.t2012 4.36035
R7181 VPWR.n214 VPWR.t3427 4.36035
R7182 VPWR.n214 VPWR.t1347 4.36035
R7183 VPWR.n213 VPWR.t1969 4.36035
R7184 VPWR.n213 VPWR.t3197 4.36035
R7185 VPWR.n212 VPWR.t3952 4.36035
R7186 VPWR.n212 VPWR.t4257 4.36035
R7187 VPWR.n211 VPWR.t1975 4.36035
R7188 VPWR.n211 VPWR.t2981 4.36035
R7189 VPWR.n210 VPWR.t7142 4.36035
R7190 VPWR.n210 VPWR.t1496 4.36035
R7191 VPWR.n209 VPWR.t1570 4.36035
R7192 VPWR.n209 VPWR.t4271 4.36035
R7193 VPWR.n208 VPWR.t2131 4.36035
R7194 VPWR.n208 VPWR.t1544 4.36035
R7195 VPWR.n218 VPWR.t5105 4.36035
R7196 VPWR.n221 VPWR.t3706 4.36035
R7197 VPWR.n223 VPWR.t1534 4.36035
R7198 VPWR.n225 VPWR.t2847 4.36035
R7199 VPWR.n227 VPWR.t4925 4.36035
R7200 VPWR.n229 VPWR.t4394 4.36035
R7201 VPWR.n231 VPWR.t611 4.36035
R7202 VPWR.n233 VPWR.t3653 4.36035
R7203 VPWR.n237 VPWR.t5167 4.36035
R7204 VPWR.n239 VPWR.t5383 4.36035
R7205 VPWR.n241 VPWR.t1305 4.36035
R7206 VPWR.n243 VPWR.t828 4.36035
R7207 VPWR.n245 VPWR.t2845 4.36035
R7208 VPWR.n247 VPWR.t5042 4.36035
R7209 VPWR.n249 VPWR.t1416 4.36035
R7210 VPWR.n251 VPWR.t2645 4.36035
R7211 VPWR.n2656 VPWR.t521 4.36035
R7212 VPWR.n2666 VPWR.t2476 4.36035
R7213 VPWR.n2668 VPWR.t386 4.36035
R7214 VPWR.n2671 VPWR.t3027 4.36035
R7215 VPWR.n2673 VPWR.t4635 4.36035
R7216 VPWR.n2675 VPWR.t4457 4.36035
R7217 VPWR.n2677 VPWR.t3332 4.36035
R7218 VPWR.n2679 VPWR.t7122 4.36035
R7219 VPWR.n2681 VPWR.t5230 4.36035
R7220 VPWR.n2686 VPWR.t1452 4.36035
R7221 VPWR.n2688 VPWR.t992 4.36035
R7222 VPWR.n2690 VPWR.t5224 4.36035
R7223 VPWR.n2692 VPWR.t2264 4.36035
R7224 VPWR.n2694 VPWR.t6156 4.36035
R7225 VPWR.n2696 VPWR.t5484 4.36035
R7226 VPWR.n2698 VPWR.t4666 4.36035
R7227 VPWR.n2082 VPWR.t2811 4.36035
R7228 VPWR.n2085 VPWR.t5655 4.36035
R7229 VPWR.n2094 VPWR.t5942 4.36035
R7230 VPWR.n2096 VPWR.t5689 4.36035
R7231 VPWR.n2055 VPWR.t739 4.36035
R7232 VPWR.n2057 VPWR.t5940 4.36035
R7233 VPWR.n2059 VPWR.t3145 4.36035
R7234 VPWR.n2061 VPWR.t1000 4.36035
R7235 VPWR.n2063 VPWR.t4070 4.36035
R7236 VPWR.n459 VPWR.t5445 4.36035
R7237 VPWR.n490 VPWR.t5327 4.36035
R7238 VPWR.n500 VPWR.t5088 4.36035
R7239 VPWR.n3033 VPWR.t3781 4.36035
R7240 VPWR.n3035 VPWR.t4895 4.36035
R7241 VPWR.n3037 VPWR.t2080 4.36035
R7242 VPWR.n3039 VPWR.t2909 4.36035
R7243 VPWR.n3041 VPWR.t1179 4.36035
R7244 VPWR.n3054 VPWR.t4648 4.36035
R7245 VPWR.n3052 VPWR.t5562 4.36035
R7246 VPWR.n3050 VPWR.t2939 4.36035
R7247 VPWR.n3048 VPWR.t3615 4.36035
R7248 VPWR.n3046 VPWR.t4711 4.36035
R7249 VPWR.n3044 VPWR.t3459 4.36035
R7250 VPWR.n173 VPWR.t5645 4.36035
R7251 VPWR.n3104 VPWR.t5954 4.36035
R7252 VPWR.n3102 VPWR.t2026 4.36035
R7253 VPWR.n3099 VPWR.t4826 4.36035
R7254 VPWR.n3097 VPWR.t5336 4.36035
R7255 VPWR.n3095 VPWR.t3510 4.36035
R7256 VPWR.n3093 VPWR.t2444 4.36035
R7257 VPWR.n3091 VPWR.t2724 4.36035
R7258 VPWR.n3089 VPWR.t1648 4.36035
R7259 VPWR.n3087 VPWR.t2820 4.36035
R7260 VPWR.n3085 VPWR.t5436 4.36035
R7261 VPWR.n3082 VPWR.t1716 4.36035
R7262 VPWR.n3080 VPWR.t5946 4.36035
R7263 VPWR.n3078 VPWR.t4200 4.36035
R7264 VPWR.n3076 VPWR.t4901 4.36035
R7265 VPWR.n3074 VPWR.t2014 4.36035
R7266 VPWR.n3072 VPWR.t5751 4.36035
R7267 VPWR.n3070 VPWR.t4633 4.36035
R7268 VPWR.n3067 VPWR.t599 4.36035
R7269 VPWR.n3065 VPWR.t2376 4.36035
R7270 VPWR.n3063 VPWR.t382 4.36035
R7271 VPWR.n3063 VPWR.t3562 4.36035
R7272 VPWR.n3062 VPWR.t6100 4.36035
R7273 VPWR.n3062 VPWR.t1697 4.36035
R7274 VPWR.n3061 VPWR.t3030 4.36035
R7275 VPWR.n3061 VPWR.t2490 4.36035
R7276 VPWR.n3060 VPWR.t894 4.36035
R7277 VPWR.n3060 VPWR.t4749 4.36035
R7278 VPWR.n3059 VPWR.t2983 4.36035
R7279 VPWR.n3059 VPWR.t3359 4.36035
R7280 VPWR.n3058 VPWR.t5547 4.36035
R7281 VPWR.n3058 VPWR.t6137 4.36035
R7282 VPWR.n3057 VPWR.t339 4.36035
R7283 VPWR.n3057 VPWR.t2468 4.36035
R7284 VPWR.n3056 VPWR.t1658 4.36035
R7285 VPWR.n3056 VPWR.t2384 4.36035
R7286 VPWR.n3066 VPWR.t3964 4.36035
R7287 VPWR.n3068 VPWR.t4597 4.36035
R7288 VPWR.n3071 VPWR.t1004 4.36035
R7289 VPWR.n3073 VPWR.t5732 4.36035
R7290 VPWR.n3075 VPWR.t3918 4.36035
R7291 VPWR.n3077 VPWR.t2550 4.36035
R7292 VPWR.n3079 VPWR.t3557 4.36035
R7293 VPWR.n3081 VPWR.t2675 4.36035
R7294 VPWR.n3084 VPWR.t3211 4.36035
R7295 VPWR.n3086 VPWR.t1799 4.36035
R7296 VPWR.n3088 VPWR.t4728 4.36035
R7297 VPWR.n3090 VPWR.t4180 4.36035
R7298 VPWR.n3092 VPWR.t4425 4.36035
R7299 VPWR.n3094 VPWR.t2252 4.36035
R7300 VPWR.n3096 VPWR.t4333 4.36035
R7301 VPWR.n3098 VPWR.t1891 4.36035
R7302 VPWR.n3100 VPWR.t2222 4.36035
R7303 VPWR.n3103 VPWR.t3123 4.36035
R7304 VPWR.n3105 VPWR.t4951 4.36035
R7305 VPWR.n3043 VPWR.t3044 4.36035
R7306 VPWR.n3045 VPWR.t2215 4.36035
R7307 VPWR.n3047 VPWR.t6188 4.36035
R7308 VPWR.n3049 VPWR.t4035 4.36035
R7309 VPWR.n3051 VPWR.t1371 4.36035
R7310 VPWR.n3053 VPWR.t2877 4.36035
R7311 VPWR.n3042 VPWR.t2137 4.36035
R7312 VPWR.n3040 VPWR.t3847 4.36035
R7313 VPWR.n3038 VPWR.t1002 4.36035
R7314 VPWR.n3036 VPWR.t4074 4.36035
R7315 VPWR.n3034 VPWR.t6302 4.36035
R7316 VPWR.n3032 VPWR.t3728 4.36035
R7317 VPWR.n3030 VPWR.t5764 4.36035
R7318 VPWR.n3028 VPWR.t5222 4.36035
R7319 VPWR.n3027 VPWR.t4542 4.36035
R7320 VPWR.n3024 VPWR.t4718 4.36035
R7321 VPWR.n553 VPWR.t2197 4.36035
R7322 VPWR.n555 VPWR.t5619 4.36035
R7323 VPWR.n556 VPWR.t5797 4.36035
R7324 VPWR.n569 VPWR.t4850 4.36035
R7325 VPWR.n570 VPWR.t4270 4.36035
R7326 VPWR.n1851 VPWR.t3055 4.36035
R7327 VPWR.n1862 VPWR.t1748 4.36035
R7328 VPWR.n1864 VPWR.t1850 4.36035
R7329 VPWR.n1866 VPWR.t1945 4.36035
R7330 VPWR.n1867 VPWR.t5165 4.36035
R7331 VPWR.n1869 VPWR.t6249 4.36035
R7332 VPWR.n497 VPWR.t4096 4.36035
R7333 VPWR.n460 VPWR.t5403 4.36035
R7334 VPWR.n361 VPWR.t1182 4.36035
R7335 VPWR.n367 VPWR.t3802 4.36035
R7336 VPWR.n365 VPWR.t4809 4.36035
R7337 VPWR.n363 VPWR.t4579 4.36035
R7338 VPWR.n1911 VPWR.t2322 4.36035
R7339 VPWR.n1905 VPWR.t5316 4.36035
R7340 VPWR.n1903 VPWR.t3621 4.36035
R7341 VPWR.n1901 VPWR.t5349 4.36035
R7342 VPWR.n1886 VPWR.t1965 4.36035
R7343 VPWR.n455 VPWR.t2512 4.36035
R7344 VPWR.n441 VPWR.t5583 4.36035
R7345 VPWR.n439 VPWR.t3777 4.36035
R7346 VPWR.n437 VPWR.t3404 4.36035
R7347 VPWR.n436 VPWR.t2454 4.36035
R7348 VPWR.n425 VPWR.t2254 4.36035
R7349 VPWR.n422 VPWR.t4662 4.36035
R7350 VPWR.n2930 VPWR.t2818 4.36035
R7351 VPWR.n2930 VPWR.t1832 4.36035
R7352 VPWR.n2931 VPWR.t5328 4.36035
R7353 VPWR.n2931 VPWR.t487 4.36035
R7354 VPWR.n2932 VPWR.t6434 4.36035
R7355 VPWR.n2932 VPWR.t5877 4.36035
R7356 VPWR.n2937 VPWR.t3199 4.36035
R7357 VPWR.n2938 VPWR.t6169 4.36035
R7358 VPWR.n3012 VPWR.t4617 4.36035
R7359 VPWR.n3010 VPWR.t3010 4.36035
R7360 VPWR.n3008 VPWR.t2985 4.36035
R7361 VPWR.n3006 VPWR.t5682 4.36035
R7362 VPWR.n3004 VPWR.t2328 4.36035
R7363 VPWR.n3002 VPWR.t2296 4.36035
R7364 VPWR.n3000 VPWR.t4501 4.36035
R7365 VPWR.n2998 VPWR.t4887 4.36035
R7366 VPWR.n2996 VPWR.t567 4.36035
R7367 VPWR.n2995 VPWR.t6300 4.36035
R7368 VPWR.n2994 VPWR.t4517 4.36035
R7369 VPWR.n2993 VPWR.t3245 4.36035
R7370 VPWR.n2992 VPWR.t3686 4.36035
R7371 VPWR.n2991 VPWR.t6235 4.36035
R7372 VPWR.n2989 VPWR.t5948 4.36035
R7373 VPWR.n2988 VPWR.t3741 4.36035
R7374 VPWR.n2986 VPWR.t1500 4.36035
R7375 VPWR.n2985 VPWR.t3747 4.36035
R7376 VPWR.n2984 VPWR.t1893 4.36035
R7377 VPWR.n2983 VPWR.t3845 4.36035
R7378 VPWR.n2982 VPWR.t5373 4.36035
R7379 VPWR.n2981 VPWR.t6183 4.36035
R7380 VPWR.n2980 VPWR.t5055 4.36035
R7381 VPWR.n2979 VPWR.t1025 4.36035
R7382 VPWR.n2977 VPWR.t4587 4.36035
R7383 VPWR.n2976 VPWR.t1809 4.36035
R7384 VPWR.n2975 VPWR.t2884 4.36035
R7385 VPWR.n2974 VPWR.t1074 4.36035
R7386 VPWR.n2973 VPWR.t1818 4.36035
R7387 VPWR.n2972 VPWR.t2470 4.36035
R7388 VPWR.n2970 VPWR.t1006 4.36035
R7389 VPWR.n2969 VPWR.t865 4.36035
R7390 VPWR.n2967 VPWR.t3528 4.36035
R7391 VPWR.n2966 VPWR.t3688 4.36035
R7392 VPWR.n2965 VPWR.t2130 4.36035
R7393 VPWR.n2964 VPWR.t4339 4.36035
R7394 VPWR.n2963 VPWR.t2309 4.36035
R7395 VPWR.n2962 VPWR.t4277 4.36035
R7396 VPWR.n2961 VPWR.t1088 4.36035
R7397 VPWR.n2960 VPWR.t3927 4.36035
R7398 VPWR.n3001 VPWR.t2345 4.36035
R7399 VPWR.n3003 VPWR.t4023 4.36035
R7400 VPWR.n3005 VPWR.t85 4.36035
R7401 VPWR.n3007 VPWR.t6359 4.36035
R7402 VPWR.n3009 VPWR.t2721 4.36035
R7403 VPWR.n3011 VPWR.t3865 4.36035
R7404 VPWR.n3014 VPWR.t6134 4.36035
R7405 VPWR.n3016 VPWR.t1977 4.36035
R7406 VPWR.n3019 VPWR.t83 4.36035
R7407 VPWR.n2936 VPWR.t886 4.36035
R7408 VPWR.n2933 VPWR.t6347 4.36035
R7409 VPWR.n438 VPWR.t3549 4.36035
R7410 VPWR.n440 VPWR.t2815 4.36035
R7411 VPWR.n442 VPWR.t5236 4.36035
R7412 VPWR.n1902 VPWR.t7076 4.36035
R7413 VPWR.n1904 VPWR.t1720 4.36035
R7414 VPWR.n1906 VPWR.t5667 4.36035
R7415 VPWR.n1908 VPWR.t4891 4.36035
R7416 VPWR.n1910 VPWR.t1064 4.36035
R7417 VPWR.n1912 VPWR.t1576 4.36035
R7418 VPWR.n1914 VPWR.t471 4.36035
R7419 VPWR.n1916 VPWR.t2875 4.36035
R7420 VPWR.n1919 VPWR.t3447 4.36035
R7421 VPWR.n1921 VPWR.t7126 4.36035
R7422 VPWR.n360 VPWR.t1058 4.36035
R7423 VPWR.n364 VPWR.t5008 4.36035
R7424 VPWR.n366 VPWR.t1373 4.36035
R7425 VPWR.n368 VPWR.t4824 4.36035
R7426 VPWR.n362 VPWR.t4404 4.36035
R7427 VPWR.n268 VPWR.t1433 4.36035
R7428 VPWR.n268 VPWR.t4230 4.36035
R7429 VPWR.n269 VPWR.t6360 4.36035
R7430 VPWR.n269 VPWR.t1176 4.36035
R7431 VPWR.n270 VPWR.t690 4.36035
R7432 VPWR.n270 VPWR.t5882 4.36035
R7433 VPWR.n271 VPWR.t3013 4.36035
R7434 VPWR.n271 VPWR.t2510 4.36035
R7435 VPWR.n272 VPWR.t5245 4.36035
R7436 VPWR.n272 VPWR.t5983 4.36035
R7437 VPWR.n2458 VPWR.t863 4.36035
R7438 VPWR.n2458 VPWR.t4191 4.36035
R7439 VPWR.n2459 VPWR.t3895 4.36035
R7440 VPWR.n2462 VPWR.t307 4.36035
R7441 VPWR.n2464 VPWR.t6148 4.36035
R7442 VPWR.n3702 VPWR.t5288 4.36035
R7443 VPWR.n3704 VPWR.t4375 4.36035
R7444 VPWR.n3705 VPWR.t4294 4.36035
R7445 VPWR.n3705 VPWR.t4131 4.36035
R7446 VPWR.n3684 VPWR.t3111 4.36035
R7447 VPWR.n3684 VPWR.t5094 4.36035
R7448 VPWR.n3713 VPWR.t1244 4.36035
R7449 VPWR.n3713 VPWR.t3440 4.36035
R7450 VPWR.n3712 VPWR.t1297 4.36035
R7451 VPWR.n3712 VPWR.t4659 4.36035
R7452 VPWR.n3711 VPWR.t2904 4.36035
R7453 VPWR.n3711 VPWR.t1540 4.36035
R7454 VPWR.n3710 VPWR.t965 4.36035
R7455 VPWR.n3710 VPWR.t1656 4.36035
R7456 VPWR.n3709 VPWR.t530 4.36035
R7457 VPWR.n3709 VPWR.t3178 4.36035
R7458 VPWR.n3708 VPWR.t3077 4.36035
R7459 VPWR.n3708 VPWR.t4287 4.36035
R7460 VPWR.n3703 VPWR.t3343 4.36035
R7461 VPWR.n3701 VPWR.t5296 4.36035
R7462 VPWR.n3699 VPWR.t6112 4.36035
R7463 VPWR.n3698 VPWR.t5864 4.36035
R7464 VPWR.n3697 VPWR.t4733 4.36035
R7465 VPWR.n3696 VPWR.t2631 4.36035
R7466 VPWR.n3695 VPWR.t6185 4.36035
R7467 VPWR.n3694 VPWR.t5502 4.36035
R7468 VPWR.n3692 VPWR.t1092 4.36035
R7469 VPWR.n3691 VPWR.t4777 4.36035
R7470 VPWR.n3690 VPWR.t1435 4.36035
R7471 VPWR.n3689 VPWR.t857 4.36035
R7472 VPWR.n3688 VPWR.t2988 4.36035
R7473 VPWR.n3687 VPWR.t5379 4.36035
R7474 VPWR.n60 VPWR.t1822 4.36035
R7475 VPWR.n3757 VPWR.t955 4.36035
R7476 VPWR.n3759 VPWR.t2424 4.36035
R7477 VPWR.n3760 VPWR.t917 4.36035
R7478 VPWR.n3761 VPWR.t6438 4.36035
R7479 VPWR.n3762 VPWR.t561 4.36035
R7480 VPWR.n3763 VPWR.t2977 4.36035
R7481 VPWR.n3764 VPWR.t7093 4.36035
R7482 VPWR.n3765 VPWR.t3135 4.36035
R7483 VPWR.n3766 VPWR.t5518 4.36035
R7484 VPWR.n3768 VPWR.t5651 4.36035
R7485 VPWR.n3769 VPWR.t75 4.36035
R7486 VPWR.n3770 VPWR.t1199 4.36035
R7487 VPWR.n3771 VPWR.t3779 4.36035
R7488 VPWR.n3772 VPWR.t5389 4.36035
R7489 VPWR.n3773 VPWR.t5267 4.36035
R7490 VPWR.n3774 VPWR.t3606 4.36035
R7491 VPWR.n38 VPWR.t6119 4.36035
R7492 VPWR.n55 VPWR.t3700 4.36035
R7493 VPWR.n54 VPWR.t2971 4.36035
R7494 VPWR.n53 VPWR.t7091 4.36035
R7495 VPWR.n52 VPWR.t3867 4.36035
R7496 VPWR.n51 VPWR.t4241 4.36035
R7497 VPWR.n50 VPWR.t3504 4.36035
R7498 VPWR.n49 VPWR.t785 4.36035
R7499 VPWR.n48 VPWR.t3682 4.36035
R7500 VPWR.n46 VPWR.t3376 4.36035
R7501 VPWR.n45 VPWR.t3439 4.36035
R7502 VPWR.n44 VPWR.t2568 4.36035
R7503 VPWR.n43 VPWR.t5735 4.36035
R7504 VPWR.n42 VPWR.t3759 4.36035
R7505 VPWR.n41 VPWR.t2689 4.36035
R7506 VPWR.n40 VPWR.t6223 4.36035
R7507 VPWR.n7 VPWR.t4947 4.36035
R7508 VPWR.n3819 VPWR.t2155 4.36035
R7509 VPWR.n3820 VPWR.t5793 4.36035
R7510 VPWR.n3821 VPWR.t4345 4.36035
R7511 VPWR.n3822 VPWR.t597 4.36035
R7512 VPWR.n3823 VPWR.t3276 4.36035
R7513 VPWR.n3824 VPWR.t2266 4.36035
R7514 VPWR.n3825 VPWR.t3328 4.36035
R7515 VPWR.n3826 VPWR.t2334 4.36035
R7516 VPWR.n3828 VPWR.t4536 4.36035
R7517 VPWR.n3829 VPWR.t3487 4.36035
R7518 VPWR.n3830 VPWR.t380 4.36035
R7519 VPWR.n3831 VPWR.t2006 4.36035
R7520 VPWR.n3832 VPWR.t749 4.36035
R7521 VPWR.n3833 VPWR.t3812 4.36035
R7522 VPWR.n3834 VPWR.t2817 4.36035
R7523 VPWR.n3835 VPWR.t4811 4.36035
R7524 VPWR.n2624 VPWR.t6449 4.36035
R7525 VPWR.n2625 VPWR.t2102 4.36035
R7526 VPWR.n2626 VPWR.t726 4.36035
R7527 VPWR.n2627 VPWR.t4897 4.36035
R7528 VPWR.n2628 VPWR.t4029 4.36035
R7529 VPWR.n2629 VPWR.t832 4.36035
R7530 VPWR.n2630 VPWR.t2804 4.36035
R7531 VPWR.n2631 VPWR.t2084 4.36035
R7532 VPWR.n2633 VPWR.t1776 4.36035
R7533 VPWR.n2634 VPWR.t1138 4.36035
R7534 VPWR.n2635 VPWR.t3555 4.36035
R7535 VPWR.n2636 VPWR.t2809 4.36035
R7536 VPWR.n2637 VPWR.t6353 4.36035
R7537 VPWR.n2638 VPWR.t3161 4.36035
R7538 VPWR.n2639 VPWR.t861 4.36035
R7539 VPWR.n2640 VPWR.t319 4.36035
R7540 VPWR.n256 VPWR.t4789 4.36035
R7541 VPWR.n2612 VPWR.t5578 4.36035
R7542 VPWR.n2613 VPWR.t826 4.36035
R7543 VPWR.n2614 VPWR.t3133 4.36035
R7544 VPWR.n2615 VPWR.t501 4.36035
R7545 VPWR.n2616 VPWR.t1016 4.36035
R7546 VPWR.n2617 VPWR.t1117 4.36035
R7547 VPWR.n2618 VPWR.t640 4.36035
R7548 VPWR.n2611 VPWR.t5130 4.36035
R7549 VPWR.n2610 VPWR.t5854 4.36035
R7550 VPWR.n2609 VPWR.t5691 4.36035
R7551 VPWR.n2608 VPWR.t3320 4.36035
R7552 VPWR.n2607 VPWR.t4289 4.36035
R7553 VPWR.n2606 VPWR.t1572 4.36035
R7554 VPWR.n2605 VPWR.t1963 4.36035
R7555 VPWR.n2604 VPWR.t6014 4.36035
R7556 VPWR.n258 VPWR.t6323 4.36035
R7557 VPWR.n2483 VPWR.t2749 4.36035
R7558 VPWR.n2484 VPWR.t2935 4.36035
R7559 VPWR.n2485 VPWR.t1039 4.36035
R7560 VPWR.n2486 VPWR.t2697 4.36035
R7561 VPWR.n2487 VPWR.t5894 4.36035
R7562 VPWR.n2488 VPWR.t3739 4.36035
R7563 VPWR.n2489 VPWR.t4658 4.36035
R7564 VPWR.n2491 VPWR.t5171 4.36035
R7565 VPWR.n2492 VPWR.t453 4.36035
R7566 VPWR.n2493 VPWR.t5199 4.36035
R7567 VPWR.n2494 VPWR.t2928 4.36035
R7568 VPWR.n2495 VPWR.t4453 4.36035
R7569 VPWR.n2496 VPWR.t1240 4.36035
R7570 VPWR.n2497 VPWR.t1309 4.36035
R7571 VPWR.n2498 VPWR.t4373 4.36035
R7572 VPWR.n265 VPWR.t868 4.36035
R7573 VPWR.n2472 VPWR.t626 4.36035
R7574 VPWR.n2473 VPWR.t1440 4.36035
R7575 VPWR.n2474 VPWR.t5860 4.36035
R7576 VPWR.n2475 VPWR.t4624 4.36035
R7577 VPWR.n2476 VPWR.t7120 4.36035
R7578 VPWR.n2477 VPWR.t4953 4.36035
R7579 VPWR.n2478 VPWR.t988 4.36035
R7580 VPWR.n2471 VPWR.t3384 4.36035
R7581 VPWR.n2470 VPWR.t65 4.36035
R7582 VPWR.n2469 VPWR.t2668 4.36035
R7583 VPWR.n2468 VPWR.t4198 4.36035
R7584 VPWR.n2467 VPWR.t2975 4.36035
R7585 VPWR.n2465 VPWR.t846 4.36035
R7586 VPWR.n2463 VPWR.t5033 4.36035
R7587 VPWR.n2461 VPWR.t773 4.36035
R7588 VPWR.n2425 VPWR.t2199 4.36035
R7589 VPWR.n2423 VPWR.t1754 4.36035
R7590 VPWR.n2421 VPWR.t834 4.36035
R7591 VPWR.n2419 VPWR.t378 4.36035
R7592 VPWR.n2417 VPWR.t5968 4.36035
R7593 VPWR.n2452 VPWR.t840 4.36035
R7594 VPWR.n2450 VPWR.t6120 4.36035
R7595 VPWR.n2450 VPWR.t5362 4.36035
R7596 VPWR.n2449 VPWR.t4102 4.36035
R7597 VPWR.n2449 VPWR.t1098 4.36035
R7598 VPWR.n2448 VPWR.t1341 4.36035
R7599 VPWR.n2448 VPWR.t1010 4.36035
R7600 VPWR.n2447 VPWR.t4945 4.36035
R7601 VPWR.n2447 VPWR.t1283 4.36035
R7602 VPWR.n2444 VPWR.t855 4.36035
R7603 VPWR.n2442 VPWR.t769 4.36035
R7604 VPWR.n2440 VPWR.t3655 4.36035
R7605 VPWR.n2438 VPWR.t4784 4.36035
R7606 VPWR.n2436 VPWR.t6012 4.36035
R7607 VPWR.n2436 VPWR.t2100 4.36035
R7608 VPWR.n2435 VPWR.t2566 4.36035
R7609 VPWR.n2435 VPWR.t1772 4.36035
R7610 VPWR.n2434 VPWR.t5081 4.36035
R7611 VPWR.n2434 VPWR.t822 4.36035
R7612 VPWR.n2433 VPWR.t2552 4.36035
R7613 VPWR.n2433 VPWR.t4475 4.36035
R7614 VPWR.n2432 VPWR.t4487 4.36035
R7615 VPWR.n2432 VPWR.t1066 4.36035
R7616 VPWR.n2431 VPWR.t5500 4.36035
R7617 VPWR.n2431 VPWR.t763 4.36035
R7618 VPWR.n2430 VPWR.t5200 4.36035
R7619 VPWR.n2430 VPWR.t457 4.36035
R7620 VPWR.n263 VPWR.t1236 4.36035
R7621 VPWR.n263 VPWR.t915 4.36035
R7622 VPWR.n2504 VPWR.t4619 4.36035
R7623 VPWR.n2507 VPWR.t4440 4.36035
R7624 VPWR.n2509 VPWR.t3905 4.36035
R7625 VPWR.n2511 VPWR.t4949 4.36035
R7626 VPWR.n2513 VPWR.t532 4.36035
R7627 VPWR.n2516 VPWR.t2686 4.36035
R7628 VPWR.n2516 VPWR.t2887 4.36035
R7629 VPWR.n2517 VPWR.t2937 4.36035
R7630 VPWR.n2517 VPWR.t5474 4.36035
R7631 VPWR.n2518 VPWR.t2946 4.36035
R7632 VPWR.n2518 VPWR.t3613 4.36035
R7633 VPWR.n2519 VPWR.t1780 4.36035
R7634 VPWR.n2532 VPWR.t2055 4.36035
R7635 VPWR.n2530 VPWR.t6251 4.36035
R7636 VPWR.n2528 VPWR.t3165 4.36035
R7637 VPWR.n2526 VPWR.t4913 4.36035
R7638 VPWR.n2524 VPWR.t3877 4.36035
R7639 VPWR.n2522 VPWR.t4021 4.36035
R7640 VPWR.n2520 VPWR.t4639 4.36035
R7641 VPWR.n2598 VPWR.t1724 4.36035
R7642 VPWR.n2596 VPWR.t4746 4.36035
R7643 VPWR.n2596 VPWR.t4147 4.36035
R7644 VPWR.n2595 VPWR.t2911 4.36035
R7645 VPWR.n2595 VPWR.t3494 4.36035
R7646 VPWR.n2594 VPWR.t3312 4.36035
R7647 VPWR.n2594 VPWR.t3086 4.36035
R7648 VPWR.n2593 VPWR.t2807 4.36035
R7649 VPWR.n2593 VPWR.t2195 4.36035
R7650 VPWR.n2592 VPWR.t5754 4.36035
R7651 VPWR.n2592 VPWR.t3128 4.36035
R7652 VPWR.n2589 VPWR.t3243 4.36035
R7653 VPWR.n2587 VPWR.t3593 4.36035
R7654 VPWR.n2585 VPWR.t2717 4.36035
R7655 VPWR.n2583 VPWR.t2236 4.36035
R7656 VPWR.n2583 VPWR.t5473 4.36035
R7657 VPWR.n2582 VPWR.t7072 4.36035
R7658 VPWR.n2582 VPWR.t5875 4.36035
R7659 VPWR.n2581 VPWR.t6356 4.36035
R7660 VPWR.n2581 VPWR.t4932 4.36035
R7661 VPWR.n2580 VPWR.t925 4.36035
R7662 VPWR.n2580 VPWR.t3408 4.36035
R7663 VPWR.n2579 VPWR.t5148 4.36035
R7664 VPWR.n2579 VPWR.t1252 4.36035
R7665 VPWR.n2578 VPWR.t4547 4.36035
R7666 VPWR.n2578 VPWR.t2410 4.36035
R7667 VPWR.n2577 VPWR.t5399 4.36035
R7668 VPWR.n2577 VPWR.t2073 4.36035
R7669 VPWR.n2576 VPWR.t5897 4.36035
R7670 VPWR.n2576 VPWR.t5309 4.36035
R7671 VPWR.n2574 VPWR.t1843 4.36035
R7672 VPWR.n2571 VPWR.t2268 4.36035
R7673 VPWR.n2569 VPWR.t1018 4.36035
R7674 VPWR.n2567 VPWR.t1992 4.36035
R7675 VPWR.n2565 VPWR.t1096 4.36035
R7676 VPWR.n2563 VPWR.t3025 4.36035
R7677 VPWR.n2560 VPWR.t4534 4.36035
R7678 VPWR.n2560 VPWR.t2104 4.36035
R7679 VPWR.n2559 VPWR.t628 4.36035
R7680 VPWR.n2559 VPWR.t5557 4.36035
R7681 VPWR.n2558 VPWR.t1984 4.36035
R7682 VPWR.n2555 VPWR.t636 4.36035
R7683 VPWR.n2553 VPWR.t396 4.36035
R7684 VPWR.n2551 VPWR.t4775 4.36035
R7685 VPWR.n2549 VPWR.t1558 4.36035
R7686 VPWR.n2547 VPWR.t1812 4.36035
R7687 VPWR.n2545 VPWR.t4751 4.36035
R7688 VPWR.n2543 VPWR.t5228 4.36035
R7689 VPWR.n0 VPWR.t759 4.36035
R7690 VPWR.n2 VPWR.t2315 4.36035
R7691 VPWR.n2 VPWR.t4295 4.36035
R7692 VPWR.n11 VPWR.t3426 4.36035
R7693 VPWR.n11 VPWR.t913 4.36035
R7694 VPWR.n12 VPWR.t1810 4.36035
R7695 VPWR.n12 VPWR.t674 4.36035
R7696 VPWR.n13 VPWR.t5683 4.36035
R7697 VPWR.n13 VPWR.t4301 4.36035
R7698 VPWR.n14 VPWR.t1714 4.36035
R7699 VPWR.n14 VPWR.t1703 4.36035
R7700 VPWR.n15 VPWR.t4855 4.36035
R7701 VPWR.n15 VPWR.t575 4.36035
R7702 VPWR.n18 VPWR.t1174 4.36035
R7703 VPWR.n20 VPWR.t2094 4.36035
R7704 VPWR.n29 VPWR.t1115 4.36035
R7705 VPWR.n29 VPWR.t3441 4.36035
R7706 VPWR.n28 VPWR.t1701 4.36035
R7707 VPWR.n28 VPWR.t3857 4.36035
R7708 VPWR.n27 VPWR.t1824 4.36035
R7709 VPWR.n27 VPWR.t3563 4.36035
R7710 VPWR.n26 VPWR.t2691 4.36035
R7711 VPWR.n26 VPWR.t3832 4.36035
R7712 VPWR.n25 VPWR.t4263 4.36035
R7713 VPWR.n25 VPWR.t4756 4.36035
R7714 VPWR.n24 VPWR.t5736 4.36035
R7715 VPWR.n24 VPWR.t3692 4.36035
R7716 VPWR.n23 VPWR.t3137 4.36035
R7717 VPWR.n23 VPWR.t4099 4.36035
R7718 VPWR.n22 VPWR.t5973 4.36035
R7719 VPWR.n22 VPWR.t6009 4.36035
R7720 VPWR.n21 VPWR.t1878 4.36035
R7721 VPWR.n3812 VPWR.t6091 4.36035
R7722 VPWR.n3810 VPWR.t5746 4.36035
R7723 VPWR.n3808 VPWR.t5472 4.36035
R7724 VPWR.n3806 VPWR.t6257 4.36035
R7725 VPWR.n3804 VPWR.t1303 4.36035
R7726 VPWR.n3802 VPWR.t1805 4.36035
R7727 VPWR.n3799 VPWR.t2973 4.36035
R7728 VPWR.n3799 VPWR.t4290 4.36035
R7729 VPWR.n3798 VPWR.t6023 4.36035
R7730 VPWR.n3795 VPWR.t3959 4.36035
R7731 VPWR.n3793 VPWR.t5458 4.36035
R7732 VPWR.n3791 VPWR.t1870 4.36035
R7733 VPWR.n3789 VPWR.t5103 4.36035
R7734 VPWR.n3787 VPWR.t4216 4.36035
R7735 VPWR.n3785 VPWR.t6267 4.36035
R7736 VPWR.n3783 VPWR.t467 4.36035
R7737 VPWR.n3781 VPWR.t519 4.36035
R7738 VPWR.n3779 VPWR.t4928 4.36035
R7739 VPWR.n3779 VPWR.t2043 4.36035
R7740 VPWR.n36 VPWR.t4613 4.36035
R7741 VPWR.n36 VPWR.t5982 4.36035
R7742 VPWR.n65 VPWR.t5664 4.36035
R7743 VPWR.n65 VPWR.t1191 4.36035
R7744 VPWR.n66 VPWR.t7079 4.36035
R7745 VPWR.n66 VPWR.t1187 4.36035
R7746 VPWR.n67 VPWR.t2978 4.36035
R7747 VPWR.n67 VPWR.t2625 4.36035
R7748 VPWR.n68 VPWR.t953 4.36035
R7749 VPWR.n68 VPWR.t5576 4.36035
R7750 VPWR.n69 VPWR.t3619 4.36035
R7751 VPWR.n69 VPWR.t1146 4.36035
R7752 VPWR.n72 VPWR.t1100 4.36035
R7753 VPWR.n74 VPWR.t4939 4.36035
R7754 VPWR.n74 VPWR.t1630 4.36035
R7755 VPWR.n75 VPWR.t3842 4.36035
R7756 VPWR.n75 VPWR.t2607 4.36035
R7757 VPWR.n76 VPWR.t1485 4.36035
R7758 VPWR.n76 VPWR.t1980 4.36035
R7759 VPWR.n77 VPWR.t4582 4.36035
R7760 VPWR.n77 VPWR.t1285 4.36035
R7761 VPWR.n78 VPWR.t2989 4.36035
R7762 VPWR.n78 VPWR.t390 4.36035
R7763 VPWR.n79 VPWR.t5687 4.36035
R7764 VPWR.n79 VPWR.t513 4.36035
R7765 VPWR.n80 VPWR.t2882 4.36035
R7766 VPWR.n80 VPWR.t1552 4.36035
R7767 VPWR.n81 VPWR.t6226 4.36035
R7768 VPWR.n81 VPWR.t550 4.36035
R7769 VPWR.n82 VPWR.t4745 4.36035
R7770 VPWR.n62 VPWR.t5226 4.36035
R7771 VPWR.n3751 VPWR.t1542 4.36035
R7772 VPWR.n3749 VPWR.t4292 4.36035
R7773 VPWR.n3747 VPWR.t3518 4.36035
R7774 VPWR.n3745 VPWR.t4923 4.36035
R7775 VPWR.n3743 VPWR.t4350 4.36035
R7776 VPWR.n3741 VPWR.t1820 4.36035
R7777 VPWR.n3738 VPWR.t663 4.36035
R7778 VPWR.n3735 VPWR.t4503 4.36035
R7779 VPWR.n3733 VPWR.t814 4.36035
R7780 VPWR.n3731 VPWR.t432 4.36035
R7781 VPWR.n3729 VPWR.t4402 4.36035
R7782 VPWR.n3727 VPWR.t2790 4.36035
R7783 VPWR.n3725 VPWR.t3695 4.36035
R7784 VPWR.n3723 VPWR.t5080 4.36035
R7785 VPWR.n3721 VPWR.t6011 4.36035
R7786 VPWR.n3719 VPWR.t4250 4.36035
R7787 VPWR.n3719 VPWR.t5802 4.36035
R7788 VPWR.n3718 VPWR.t1374 4.36035
R7789 VPWR.n3718 VPWR.t650 4.36035
R7790 VPWR.n94 VPWR.t2280 4.36035
R7791 VPWR.n94 VPWR.t4885 4.36035
R7792 VPWR.n93 VPWR.t77 4.36035
R7793 VPWR.n93 VPWR.t3707 4.36035
R7794 VPWR.n92 VPWR.t637 4.36035
R7795 VPWR.n92 VPWR.t357 4.36035
R7796 VPWR.n91 VPWR.t4730 4.36035
R7797 VPWR.n91 VPWR.t1301 4.36035
R7798 VPWR.n90 VPWR.t1470 4.36035
R7799 VPWR.n90 VPWR.t1365 4.36035
R7800 VPWR.n89 VPWR.t1508 4.36035
R7801 VPWR.n89 VPWR.t3126 4.36035
R7802 VPWR.n3722 VPWR.t2311 4.36035
R7803 VPWR.n3724 VPWR.t2372 4.36035
R7804 VPWR.n3726 VPWR.t2211 4.36035
R7805 VPWR.n3728 VPWR.t6197 4.36035
R7806 VPWR.n3730 VPWR.t345 4.36035
R7807 VPWR.n3732 VPWR.t3526 4.36035
R7808 VPWR.n3734 VPWR.t5843 4.36035
R7809 VPWR.n3736 VPWR.t6206 4.36035
R7810 VPWR.n3740 VPWR.t5536 4.36035
R7811 VPWR.n3742 VPWR.t2683 4.36035
R7812 VPWR.n3744 VPWR.t455 4.36035
R7813 VPWR.n3746 VPWR.t4735 4.36035
R7814 VPWR.n3748 VPWR.t4779 4.36035
R7815 VPWR.n3750 VPWR.t4141 4.36035
R7816 VPWR.n3752 VPWR.t6124 4.36035
R7817 VPWR.n83 VPWR.t4556 4.36035
R7818 VPWR.n70 VPWR.t5727 4.36035
R7819 VPWR.n3782 VPWR.t5364 4.36035
R7820 VPWR.n3784 VPWR.t1043 4.36035
R7821 VPWR.n3786 VPWR.t6225 4.36035
R7822 VPWR.n3788 VPWR.t5478 4.36035
R7823 VPWR.n3790 VPWR.t5686 4.36035
R7824 VPWR.n3792 VPWR.t3553 4.36035
R7825 VPWR.n3794 VPWR.t368 4.36035
R7826 VPWR.n3796 VPWR.t957 4.36035
R7827 VPWR.n3801 VPWR.t6295 4.36035
R7828 VPWR.n3803 VPWR.t1662 4.36035
R7829 VPWR.n3805 VPWR.t5697 4.36035
R7830 VPWR.n3807 VPWR.t4027 4.36035
R7831 VPWR.n3809 VPWR.t7139 4.36035
R7832 VPWR.n3811 VPWR.t6432 4.36035
R7833 VPWR.n3813 VPWR.t2038 4.36035
R7834 VPWR.n19 VPWR.t3259 4.36035
R7835 VPWR.n16 VPWR.t3937 4.36035
R7836 VPWR.n2542 VPWR.t6080 4.36035
R7837 VPWR.n2544 VPWR.t4782 4.36035
R7838 VPWR.n2546 VPWR.t617 4.36035
R7839 VPWR.n2548 VPWR.t5234 4.36035
R7840 VPWR.n2550 VPWR.t853 4.36035
R7841 VPWR.n2552 VPWR.t5441 4.36035
R7842 VPWR.n2554 VPWR.t4813 4.36035
R7843 VPWR.n2556 VPWR.t3330 4.36035
R7844 VPWR.n2562 VPWR.t4899 4.36035
R7845 VPWR.n2564 VPWR.t3520 4.36035
R7846 VPWR.n2566 VPWR.t1634 4.36035
R7847 VPWR.n2568 VPWR.t420 4.36035
R7848 VPWR.n2570 VPWR.t4738 4.36035
R7849 VPWR.n2572 VPWR.t2243 4.36035
R7850 VPWR.n2586 VPWR.t2069 4.36035
R7851 VPWR.n2588 VPWR.t4753 4.36035
R7852 VPWR.n2591 VPWR.t630 4.36035
R7853 VPWR.n260 VPWR.t4416 4.36035
R7854 VPWR.n2521 VPWR.t5867 4.36035
R7855 VPWR.n2523 VPWR.t3875 4.36035
R7856 VPWR.n2525 VPWR.t2613 4.36035
R7857 VPWR.n2527 VPWR.t6093 4.36035
R7858 VPWR.n2529 VPWR.t5830 4.36035
R7859 VPWR.n2531 VPWR.t4763 4.36035
R7860 VPWR.n2533 VPWR.t6204 4.36035
R7861 VPWR.n2514 VPWR.t2139 4.36035
R7862 VPWR.n2512 VPWR.t4104 4.36035
R7863 VPWR.n2510 VPWR.t4166 4.36035
R7864 VPWR.n2508 VPWR.t5330 4.36035
R7865 VPWR.n2506 VPWR.t1376 4.36035
R7866 VPWR.n2439 VPWR.t3084 4.36035
R7867 VPWR.n2441 VPWR.t2063 4.36035
R7868 VPWR.n2443 VPWR.t4176 4.36035
R7869 VPWR.n2446 VPWR.t4772 4.36035
R7870 VPWR.n2453 VPWR.t5762 4.36035
R7871 VPWR.n2418 VPWR.t4553 4.36035
R7872 VPWR.n2420 VPWR.t712 4.36035
R7873 VPWR.n2422 VPWR.t2813 4.36035
R7874 VPWR.n2424 VPWR.t2116 4.36035
R7875 VPWR.n2426 VPWR.t4489 4.36035
R7876 VPWR.n3700 VPWR.n3685 4.35925
R7877 VPWR.n2466 VPWR.n266 4.35925
R7878 VPWR.t1210 VPWR.n3450 4.35924
R7879 VPWR.t5523 VPWR.n3465 4.35924
R7880 VPWR.t2387 VPWR.n3480 4.35924
R7881 VPWR.t2111 VPWR.n3495 4.35924
R7882 VPWR.t2671 VPWR.n3510 4.35924
R7883 VPWR.t2787 VPWR.n3525 4.35924
R7884 VPWR.t2329 VPWR.n3540 4.35924
R7885 VPWR.t4972 VPWR.n3555 4.35924
R7886 VPWR.t1733 VPWR.n3570 4.35924
R7887 VPWR.t2742 VPWR.n3585 4.35924
R7888 VPWR.t7101 VPWR.n3600 4.35924
R7889 VPWR.t2785 VPWR.n3615 4.35924
R7890 VPWR.t3924 VPWR.n3630 4.35924
R7891 VPWR.t80 VPWR.n3645 4.35924
R7892 VPWR.t3722 VPWR.n3660 4.35924
R7893 VPWR.t4346 VPWR.n3675 4.35924
R7894 VPWR.n1341 VPWR.n1276 4.35924
R7895 VPWR.n1211 VPWR.n1172 4.35924
R7896 VPWR VPWR.n1087 4.35924
R7897 VPWR VPWR.t4045 4.35924
R7898 VPWR.n2108 VPWR.t5768 4.35924
R7899 VPWR.n303 VPWR.t3190 4.35924
R7900 VPWR.t6201 VPWR 4.35924
R7901 VPWR.t3523 VPWR 4.35924
R7902 VPWR.t3642 VPWR 4.35924
R7903 VPWR.n2308 VPWR.t2449 4.35924
R7904 VPWR.n2051 VPWR.t3391 4.35924
R7905 VPWR.n2092 VPWR.n2065 4.35924
R7906 VPWR.n475 VPWR.n458 4.35924
R7907 VPWR VPWR.n371 4.35924
R7908 VPWR.n2460 VPWR.n267 4.35924
R7909 VPWR.n2451 VPWR.n2427 4.35924
R7910 VPWR.n3385 VPWR.n101 4.35923
R7911 VPWR.n3414 VPWR.n98 4.35923
R7912 VPWR VPWR.n954 4.35923
R7913 VPWR.n1009 VPWR.n935 4.35923
R7914 VPWR.n1359 VPWR.n1035 4.35923
R7915 VPWR.n1460 VPWR.n1389 4.35923
R7916 VPWR.n1429 VPWR.n1400 4.35923
R7917 VPWR.n3354 VPWR.n3353 4.35923
R7918 VPWR.n865 VPWR.n853 4.35923
R7919 VPWR.n895 VPWR.n833 4.35923
R7920 VPWR.n1325 VPWR.t4523 4.35923
R7921 VPWR.n1295 VPWR.t4468 4.35923
R7922 VPWR.n1655 VPWR.n822 4.35923
R7923 VPWR.n3301 VPWR.n3262 4.35923
R7924 VPWR.n1240 VPWR.t3906 4.35923
R7925 VPWR.n1686 VPWR.n735 4.35923
R7926 VPWR.n3255 VPWR.n3254 4.35923
R7927 VPWR.n3175 VPWR.t3202 4.35923
R7928 VPWR.n3205 VPWR.n143 4.35923
R7929 VPWR.n1799 VPWR.n1783 4.35923
R7930 VPWR.n1191 VPWR.n1175 4.35923
R7931 VPWR.n1728 VPWR.n724 4.35923
R7932 VPWR.n1778 VPWR.n1777 4.35923
R7933 VPWR.n648 VPWR.t4340 4.35923
R7934 VPWR.t5099 VPWR.n3144 4.35923
R7935 VPWR.n681 VPWR.n628 4.35923
R7936 VPWR.n1829 VPWR.n612 4.35923
R7937 VPWR.n1107 VPWR.n1093 4.35923
R7938 VPWR.n1141 VPWR.n1088 4.35923
R7939 VPWR.n1992 VPWR.n1936 4.35923
R7940 VPWR.n1953 VPWR.t2019 4.35923
R7941 VPWR.n2861 VPWR.n2860 4.35923
R7942 VPWR.n2903 VPWR.n2874 4.35923
R7943 VPWR.n2126 VPWR.t6179 4.35923
R7944 VPWR.t427 VPWR.n2167 4.35923
R7945 VPWR.t5541 VPWR.n331 4.35923
R7946 VPWR.n2250 VPWR.t4525 4.35923
R7947 VPWR.n2290 VPWR.t5107 4.35923
R7948 VPWR.t5555 VPWR.n2219 4.35923
R7949 VPWR.n2368 VPWR.n2327 4.35923
R7950 VPWR.n2358 VPWR.n2328 4.35923
R7951 VPWR.n2349 VPWR.n2329 4.35923
R7952 VPWR.n2339 VPWR.n2330 4.35923
R7953 VPWR.n2324 VPWR.n2323 4.35923
R7954 VPWR.n2779 VPWR.t871 4.35923
R7955 VPWR.n2033 VPWR.t5367 4.35923
R7956 VPWR.t7131 VPWR.n2746 4.35923
R7957 VPWR.n2808 VPWR.t2312 4.35923
R7958 VPWR.n2084 VPWR.n2066 4.35923
R7959 VPWR.n2685 VPWR.n199 4.35923
R7960 VPWR.n2655 VPWR.n202 4.35923
R7961 VPWR.n236 VPWR.n205 4.35923
R7962 VPWR.t2136 VPWR.n3055 4.35923
R7963 VPWR.n3083 VPWR.t3210 4.35923
R7964 VPWR.n558 VPWR.n541 4.35923
R7965 VPWR.n1861 VPWR.t1747 4.35923
R7966 VPWR.n588 VPWR.n525 4.35923
R7967 VPWR.n511 VPWR.n510 4.35923
R7968 VPWR.n2997 VPWR.n2956 4.35923
R7969 VPWR.n2987 VPWR.n2957 4.35923
R7970 VPWR.n2978 VPWR.n2958 4.35923
R7971 VPWR.n2968 VPWR.n2959 4.35923
R7972 VPWR.n3013 VPWR.t6133 4.35923
R7973 VPWR.n2929 VPWR.n180 4.35923
R7974 VPWR.n2951 VPWR.n2950 4.35923
R7975 VPWR.n405 VPWR.n395 4.35923
R7976 VPWR.n429 VPWR.n378 4.35923
R7977 VPWR.n416 VPWR.n385 4.35923
R7978 VPWR.n370 VPWR.n369 4.35923
R7979 VPWR.n1913 VPWR.t470 4.35923
R7980 VPWR.n1895 VPWR.n372 4.35923
R7981 VPWR.n445 VPWR.n374 4.35923
R7982 VPWR.n2445 VPWR.n2428 4.35923
R7983 VPWR.n2515 VPWR.n261 4.35923
R7984 VPWR.n2590 VPWR.n2537 4.35923
R7985 VPWR.n2561 VPWR.n2540 4.35923
R7986 VPWR.n17 VPWR.n10 4.35923
R7987 VPWR.n3800 VPWR.n33 4.35923
R7988 VPWR.n71 VPWR.n64 4.35923
R7989 VPWR.n3739 VPWR.n86 4.35923
R7990 VPWR.n2377 VPWR.n2326 4.35916
R7991 VPWR.n2999 VPWR.n2955 4.35916
R7992 VPWR.n1509 VPWR.n1508 4.35914
R7993 VPWR.n1507 VPWR.n1506 4.35914
R7994 VPWR.n1489 VPWR.n1022 4.35914
R7995 VPWR.n1482 VPWR.n1026 4.35914
R7996 VPWR.n1474 VPWR.n1029 4.35914
R7997 VPWR.n1069 VPWR.n1064 4.35914
R7998 VPWR.n1077 VPWR.n1059 4.35914
R7999 VPWR.n1545 VPWR.n1542 4.35914
R8000 VPWR.n1553 VPWR.n1535 4.35914
R8001 VPWR.n1562 VPWR.n1534 4.35914
R8002 VPWR.n1571 VPWR.n1570 4.35914
R8003 VPWR.n1573 VPWR.n1572 4.35914
R8004 VPWR.n1582 VPWR.n1526 4.35914
R8005 VPWR.n1591 VPWR.n1525 4.35914
R8006 VPWR.n1599 VPWR.n1524 4.35914
R8007 VPWR.n1523 VPWR.n1018 4.35914
R8008 VPWR.n1522 VPWR.n1521 4.35914
R8009 VPWR.n1621 VPWR.n923 4.35914
R8010 VPWR.n1637 VPWR.n912 4.35914
R8011 VPWR.n1608 VPWR.n929 4.35914
R8012 VPWR.n1005 VPWR.n938 4.35914
R8013 VPWR.n994 VPWR.n947 4.35914
R8014 VPWR.n966 VPWR.n965 4.35914
R8015 VPWR.n981 VPWR.n955 4.35914
R8016 VPWR.n3435 VPWR.n3434 4.35914
R8017 VPWR.n3416 VPWR.n97 4.35914
R8018 VPWR.n3397 VPWR.n99 4.35914
R8019 VPWR.n3387 VPWR.n100 4.35914
R8020 VPWR.n1424 VPWR.n1406 4.35914
R8021 VPWR.n1451 VPWR.n1392 4.35914
R8022 VPWR.n1468 VPWR.n1386 4.35914
R8023 VPWR.n1385 VPWR.n1384 4.35914
R8024 VPWR.n1350 VPWR.n1038 4.35914
R8025 VPWR.n1668 VPWR.n819 4.35914
R8026 VPWR.n1309 VPWR.n1278 4.35914
R8027 VPWR.n878 VPWR.n846 4.35914
R8028 VPWR.n3324 VPWR.n115 4.35914
R8029 VPWR.n3369 VPWR.n3355 4.35914
R8030 VPWR.n3312 VPWR.n3256 4.35914
R8031 VPWR.n3228 VPWR.n128 4.35914
R8032 VPWR.n3286 VPWR.n3269 4.35914
R8033 VPWR.n783 VPWR.n756 4.35914
R8034 VPWR.n815 VPWR.n743 4.35914
R8035 VPWR.n1703 VPWR.n729 4.35914
R8036 VPWR.n1260 VPWR.n1229 4.35914
R8037 VPWR.n1744 VPWR.n714 4.35914
R8038 VPWR.n1715 VPWR.n725 4.35914
R8039 VPWR.n1811 VPWR.n1779 4.35914
R8040 VPWR.n3218 VPWR.n136 4.35914
R8041 VPWR.n3191 VPWR.n151 4.35914
R8042 VPWR.n165 VPWR.t2793 4.35914
R8043 VPWR.n1122 VPWR.t1222 4.35914
R8044 VPWR.n694 VPWR.n624 4.35914
R8045 VPWR.n1841 VPWR.n604 4.35914
R8046 VPWR.n665 VPWR.n632 4.35914
R8047 VPWR.n3153 VPWR.t5833 4.35914
R8048 VPWR.n3114 VPWR.t3271 4.35914
R8049 VPWR.n2916 VPWR.n2866 4.35914
R8050 VPWR.n2832 VPWR.n187 4.35914
R8051 VPWR.n1972 VPWR.n1937 4.35914
R8052 VPWR.n2002 VPWR.t6077 4.35914
R8053 VPWR.n2176 VPWR.t3617 4.35914
R8054 VPWR.n2140 VPWR.t496 4.35914
R8055 VPWR.n340 VPWR.t1561 4.35914
R8056 VPWR.n2268 VPWR.t3626 4.35914
R8057 VPWR.n2228 VPWR.t547 4.35914
R8058 VPWR.n2192 VPWR.t1247 4.35914
R8059 VPWR.n2319 VPWR.n2318 4.35914
R8060 VPWR.n2826 VPWR.t4336 4.35914
R8061 VPWR.n2712 VPWR.n193 4.35914
R8062 VPWR.n2759 VPWR.t3393 4.35914
R8063 VPWR.n216 VPWR.n207 4.35914
R8064 VPWR.n234 VPWR.n206 4.35914
R8065 VPWR.n252 VPWR.n204 4.35914
R8066 VPWR.n2653 VPWR.n203 4.35914
R8067 VPWR.n2664 VPWR.n201 4.35914
R8068 VPWR.n2682 VPWR.n200 4.35914
R8069 VPWR.n2700 VPWR.n198 4.35914
R8070 VPWR.n2080 VPWR.t5849 4.35914
R8071 VPWR.n1877 VPWR.n512 4.35914
R8072 VPWR.n598 VPWR.n523 4.35914
R8073 VPWR.n3026 VPWR.n176 4.35914
R8074 VPWR.n573 VPWR.n535 4.35914
R8075 VPWR.n3064 VPWR.t2375 4.35914
R8076 VPWR.n3101 VPWR.t2025 4.35914
R8077 VPWR.n454 VPWR.n373 4.35914
R8078 VPWR.n421 VPWR.n381 4.35914
R8079 VPWR.n2925 VPWR.n181 4.35914
R8080 VPWR.n3018 VPWR.n2953 4.35914
R8081 VPWR.n3693 VPWR.n3686 4.35914
R8082 VPWR.n3758 VPWR.n59 4.35914
R8083 VPWR.n3767 VPWR.n58 4.35914
R8084 VPWR.n57 VPWR.n56 4.35914
R8085 VPWR.n47 VPWR.n39 4.35914
R8086 VPWR.n3818 VPWR.n6 4.35914
R8087 VPWR.n3827 VPWR.n5 4.35914
R8088 VPWR.n2622 VPWR.n4 4.35914
R8089 VPWR.n2632 VPWR.n2623 4.35914
R8090 VPWR.n2641 VPWR.n2621 4.35914
R8091 VPWR.n2620 VPWR.n2619 4.35914
R8092 VPWR.n2603 VPWR.n257 4.35914
R8093 VPWR.n2490 VPWR.n2482 4.35914
R8094 VPWR.n2499 VPWR.n2481 4.35914
R8095 VPWR.n2480 VPWR.n2479 4.35914
R8096 VPWR.n3707 VPWR.n3706 4.35914
R8097 VPWR.n3720 VPWR.n88 4.35914
R8098 VPWR.n3737 VPWR.n87 4.35914
R8099 VPWR.n85 VPWR.n84 4.35914
R8100 VPWR.n73 VPWR.n63 4.35914
R8101 VPWR.n3780 VPWR.n35 4.35914
R8102 VPWR.n3797 VPWR.n34 4.35914
R8103 VPWR.n32 VPWR.n9 4.35914
R8104 VPWR.n31 VPWR.n30 4.35914
R8105 VPWR.n3840 VPWR.n1 4.35914
R8106 VPWR.n2557 VPWR.n2541 4.35914
R8107 VPWR.n2573 VPWR.n2539 4.35914
R8108 VPWR.n2584 VPWR.n2538 4.35914
R8109 VPWR.n2597 VPWR.n2536 4.35914
R8110 VPWR.n2535 VPWR.n2534 4.35914
R8111 VPWR.n2505 VPWR.n262 4.35914
R8112 VPWR.n2437 VPWR.n2429 4.35914
R8113 VPWR VPWR.n920 4.35913
R8114 VPWR VPWR.t3170 4.35913
R8115 VPWR VPWR.n2325 4.35913
R8116 VPWR.n1431 VPWR.t2681 4.35083
R8117 VPWR.n1327 VPWR.t5059 4.35083
R8118 VPWR.n863 VPWR.t6775 4.35083
R8119 VPWR.n1235 VPWR.t1170 4.35083
R8120 VPWR.n3201 VPWR.t6679 4.35083
R8121 VPWR.n1808 VPWR.t5600 4.35083
R8122 VPWR.n592 VPWR.t202 4.35083
R8123 VPWR.n1574 VPWR.t6673 4.34469
R8124 VPWR.n1594 VPWR.t5832 4.34469
R8125 VPWR.n1598 VPWR.t109 4.34469
R8126 VPWR.n1518 VPWR.t3560 4.34469
R8127 VPWR.n1519 VPWR.t5928 4.34469
R8128 VPWR.n1520 VPWR.t5932 4.34469
R8129 VPWR.n1486 VPWR.t2771 4.34469
R8130 VPWR.n1475 VPWR.t6765 4.34469
R8131 VPWR.n1462 VPWR.t5816 4.34469
R8132 VPWR.n1445 VPWR.t6761 4.34469
R8133 VPWR.n1612 VPWR.t107 4.34469
R8134 VPWR.n1012 VPWR.t44 4.34469
R8135 VPWR.n3380 VPWR.t2587 4.34469
R8136 VPWR.n983 VPWR.t1259 4.34469
R8137 VPWR.n989 VPWR.t4882 4.34469
R8138 VPWR.n991 VPWR.t1162 4.34469
R8139 VPWR.n1443 VPWR.t2769 4.34469
R8140 VPWR.n1446 VPWR.t3490 4.34469
R8141 VPWR.n1294 VPWR.t3678 4.34469
R8142 VPWR.n1288 VPWR.t3680 4.34469
R8143 VPWR.n1286 VPWR.t2773 4.34469
R8144 VPWR.n1665 VPWR.t909 4.34469
R8145 VPWR.n1661 VPWR.t644 4.34469
R8146 VPWR.n1660 VPWR.t2448 4.34469
R8147 VPWR.n1649 VPWR.t6809 4.34469
R8148 VPWR.n3334 VPWR.t1255 4.34469
R8149 VPWR.n859 VPWR.t980 4.34469
R8150 VPWR.n880 VPWR.t111 4.34469
R8151 VPWR.n1659 VPWR.t646 4.34469
R8152 VPWR.n1705 VPWR.t5739 4.34469
R8153 VPWR.n1681 VPWR.t5847 4.34469
R8154 VPWR.n808 VPWR.t117 4.34469
R8155 VPWR.n771 VPWR.t209 4.34469
R8156 VPWR.n3237 VPWR.t113 4.34469
R8157 VPWR.n3252 VPWR.t982 4.34469
R8158 VPWR.n3304 VPWR.t3634 4.34469
R8159 VPWR.n3311 VPWR.t6992 4.34469
R8160 VPWR.n3315 VPWR.t2955 4.34469
R8161 VPWR.n770 VPWR.t6864 4.34469
R8162 VPWR.n1701 VPWR.t335 4.34469
R8163 VPWR.n1193 VPWR.t2596 4.34469
R8164 VPWR.n1189 VPWR.t2728 4.34469
R8165 VPWR.n1181 VPWR.t4720 4.34469
R8166 VPWR.n1756 VPWR.t126 4.34469
R8167 VPWR.n1810 VPWR.t6425 4.34469
R8168 VPWR.n1806 VPWR.t5881 4.34469
R8169 VPWR.n1801 VPWR.t2167 4.34469
R8170 VPWR.n3209 VPWR.t476 4.34469
R8171 VPWR.n1108 VPWR.t937 4.34469
R8172 VPWR.n689 VPWR.t1762 4.34469
R8173 VPWR.n686 VPWR.t1289 4.34469
R8174 VPWR.n667 VPWR.t6374 4.34469
R8175 VPWR.n673 VPWR.t5540 4.34469
R8176 VPWR.n677 VPWR.t6588 4.34469
R8177 VPWR.n687 VPWR.t6600 4.34469
R8178 VPWR.n691 VPWR.t2649 4.34469
R8179 VPWR.n2843 VPWR.t4467 4.34469
R8180 VPWR.n2914 VPWR.t5044 4.34469
R8181 VPWR.n2782 VPWR.t4551 4.34469
R8182 VPWR.n600 VPWR.t185 4.34469
R8183 VPWR.n571 VPWR.t6953 4.34469
R8184 VPWR.n554 VPWR.t4474 4.34469
R8185 VPWR.n547 VPWR.t2332 4.34469
R8186 VPWR.n597 VPWR.t133 4.34469
R8187 VPWR.n2941 VPWR.t2576 4.34469
R8188 VPWR.n2946 VPWR.t2703 4.34469
R8189 VPWR.n2949 VPWR.t5447 4.34469
R8190 VPWR.n2939 VPWR.t2707 4.34469
R8191 VPWR.n2928 VPWR.t5568 4.34469
R8192 VPWR.n1458 VPWR.t4603 4.32513
R8193 VPWR.n1454 VPWR.t4601 4.32513
R8194 VPWR.n1453 VPWR.t6279 4.32513
R8195 VPWR.n1457 VPWR.t6281 4.32513
R8196 VPWR.n1459 VPWR.t2656 4.32513
R8197 VPWR.n1463 VPWR.t2658 4.32513
R8198 VPWR.n1299 VPWR.t1427 4.32513
R8199 VPWR.n1299 VPWR.t5203 4.32513
R8200 VPWR.n1297 VPWR.t1425 4.32513
R8201 VPWR.n1297 VPWR.t5202 4.32513
R8202 VPWR.n1450 VPWR.t5040 4.32122
R8203 VPWR.n1563 VPWR.t4124 4.31388
R8204 VPWR.n1566 VPWR.t5873 4.31388
R8205 VPWR.n1569 VPWR.t5304 4.31388
R8206 VPWR.n1532 VPWR.t2591 4.31388
R8207 VPWR.n1583 VPWR.t2149 4.31388
R8208 VPWR.n1586 VPWR.t2307 4.31388
R8209 VPWR.n1592 VPWR.t2581 4.31388
R8210 VPWR.n1593 VPWR.t5387 4.31388
R8211 VPWR.n1601 VPWR.t7108 4.30388
R8212 VPWR.n3327 VPWR.t6403 4.30388
R8213 VPWR.n1317 VPWR.t4094 4.30388
R8214 VPWR.n3232 VPWR.t6528 4.30388
R8215 VPWR.n3251 VPWR.t4210 4.30388
R8216 VPWR.n3299 VPWR.t4522 4.30388
R8217 VPWR.n3243 VPWR.t6967 4.30388
R8218 VPWR.n3225 VPWR.t6770 4.30388
R8219 VPWR.n1807 VPWR.t974 4.30388
R8220 VPWR.n2910 VPWR.t6961 4.30388
R8221 VPWR.n2801 VPWR.t2765 4.30388
R8222 VPWR.n594 VPWR.t5004 4.30388
R8223 VPWR.n589 VPWR.t3274 4.30388
R8224 VPWR.n595 VPWR.t5161 4.30388
R8225 VPWR.n404 VPWR.t3402 4.30388
R8226 VPWR.n1054 VPWR.t1738 4.30165
R8227 VPWR.n1042 VPWR.t1525 4.30165
R8228 VPWR.n1046 VPWR.t5719 4.30165
R8229 VPWR.n1050 VPWR.t2570 4.30165
R8230 VPWR.n1357 VPWR.t4869 4.30165
R8231 VPWR.n1360 VPWR.t5936 4.30165
R8232 VPWR.n1364 VPWR.t2484 4.30165
R8233 VPWR.n1467 VPWR.t2153 4.30165
R8234 VPWR.n1355 VPWR.t3790 4.30165
R8235 VPWR.n1349 VPWR.t5661 4.30165
R8236 VPWR.n1051 VPWR.t1742 4.30165
R8237 VPWR.n1047 VPWR.t1213 4.30165
R8238 VPWR.n1041 VPWR.t1529 4.30165
R8239 VPWR.n1275 VPWR.t3278 4.30165
R8240 VPWR.n1271 VPWR.t2274 4.30165
R8241 VPWR.n1271 VPWR.t2913 4.30165
R8242 VPWR.n1268 VPWR.t3711 4.30165
R8243 VPWR.n1343 VPWR.t4382 4.30165
R8244 VPWR.n1337 VPWR.t4865 4.30165
R8245 VPWR.n1334 VPWR.t3096 4.30165
R8246 VPWR.n1308 VPWR.t1955 4.30165
R8247 VPWR.n1306 VPWR.t3508 4.30165
R8248 VPWR.n1305 VPWR.t3883 4.30165
R8249 VPWR.n1333 VPWR.t3151 4.30165
R8250 VPWR.n1340 VPWR.t921 4.30165
R8251 VPWR.n1269 VPWR.t5723 4.30165
R8252 VPWR.n1272 VPWR.t1941 4.30165
R8253 VPWR.n1224 VPWR.t2879 4.30165
R8254 VPWR.n1223 VPWR.t2184 4.30165
R8255 VPWR.n1219 VPWR.t2278 4.30165
R8256 VPWR.n1261 VPWR.t2486 4.30165
R8257 VPWR.n1255 VPWR.t3891 4.30165
R8258 VPWR.n1253 VPWR.t2224 4.30165
R8259 VPWR.n1698 VPWR.t2747 4.30165
R8260 VPWR.n1696 VPWR.t4834 4.30165
R8261 VPWR.n1704 VPWR.t4430 4.30165
R8262 VPWR.n1248 VPWR.t1070 4.30165
R8263 VPWR.n1252 VPWR.t6060 4.30165
R8264 VPWR.n1254 VPWR.t6062 4.30165
R8265 VPWR.n1221 VPWR.t1104 4.30165
R8266 VPWR.n1225 VPWR.t5627 4.30165
R8267 VPWR.n1226 VPWR.t5623 4.30165
R8268 VPWR.n1169 VPWR.t842 4.30165
R8269 VPWR.n1165 VPWR.t4478 4.30165
R8270 VPWR.n1164 VPWR.t4484 4.30165
R8271 VPWR.n1160 VPWR.t905 4.30165
R8272 VPWR.n1212 VPWR.t4281 4.30165
R8273 VPWR.n1205 VPWR.t5411 4.30165
R8274 VPWR.n1204 VPWR.t1273 4.30165
R8275 VPWR.n1714 VPWR.t4438 4.30165
R8276 VPWR.n1718 VPWR.t1051 4.30165
R8277 VPWR.n1719 VPWR.t1588 4.30165
R8278 VPWR.n1713 VPWR.t1317 4.30165
R8279 VPWR.n726 VPWR.t1319 4.30165
R8280 VPWR.n1180 VPWR.t3059 4.30165
R8281 VPWR.n1185 VPWR.t2126 4.30165
R8282 VPWR.n1186 VPWR.t4156 4.30165
R8283 VPWR.n1190 VPWR.t1687 4.30165
R8284 VPWR.n1194 VPWR.t6246 4.30165
R8285 VPWR.n1197 VPWR.t2395 4.30165
R8286 VPWR.n1200 VPWR.t2399 4.30165
R8287 VPWR.n1203 VPWR.t1868 4.30165
R8288 VPWR.n1210 VPWR.t3587 4.30165
R8289 VPWR.n1213 VPWR.t1078 4.30165
R8290 VPWR.n1161 VPWR.t6175 4.30165
R8291 VPWR.n1168 VPWR.t7106 4.30165
R8292 VPWR.n1085 VPWR.t2526 4.30165
R8293 VPWR.n1085 VPWR.t6176 4.30165
R8294 VPWR.n1084 VPWR.t3737 4.30165
R8295 VPWR.n1084 VPWR.t5906 4.30165
R8296 VPWR.n1156 VPWR.t4509 4.30165
R8297 VPWR.n1148 VPWR.t1860 4.30165
R8298 VPWR.n1137 VPWR.t1586 4.30165
R8299 VPWR.n1134 VPWR.t1683 4.30165
R8300 VPWR.n1129 VPWR.t542 4.30165
R8301 VPWR.n1127 VPWR.t5614 4.30165
R8302 VPWR.n1128 VPWR.t536 4.30165
R8303 VPWR.n1138 VPWR.t3975 4.30165
R8304 VPWR.n1082 VPWR.t5910 4.30165
R8305 VPWR.n1988 VPWR.t5886 4.30165
R8306 VPWR.n1984 VPWR.t3000 4.30165
R8307 VPWR.n1982 VPWR.t2370 4.30165
R8308 VPWR.n1967 VPWR.t3073 4.30165
R8309 VPWR.n1964 VPWR.t5693 4.30165
R8310 VPWR.n1963 VPWR.t4412 4.30165
R8311 VPWR.n1959 VPWR.t2120 4.30165
R8312 VPWR.n1962 VPWR.t5528 4.30165
R8313 VPWR.n1979 VPWR.t5890 4.30165
R8314 VPWR.n1983 VPWR.t6255 4.30165
R8315 VPWR.n1987 VPWR.t6132 4.30165
R8316 VPWR.n1989 VPWR.t1388 4.30165
R8317 VPWR.n2131 VPWR.t5602 4.30165
R8318 VPWR.n2028 VPWR.t3173 4.30165
R8319 VPWR.n2026 VPWR.t1406 4.30165
R8320 VPWR.n2022 VPWR.t4532 4.30165
R8321 VPWR.n2722 VPWR.t609 4.30165
R8322 VPWR.n2724 VPWR.t1119 4.30165
R8323 VPWR.n2727 VPWR.t5952 4.30165
R8324 VPWR.n2723 VPWR.t5992 4.30165
R8325 VPWR.n2719 VPWR.t1125 4.30165
R8326 VPWR.n2718 VPWR.t5322 4.30165
R8327 VPWR.n2021 VPWR.t1604 4.30165
R8328 VPWR.n2025 VPWR.t2203 4.30165
R8329 VPWR.n2027 VPWR.t2209 4.30165
R8330 VPWR.n2077 VPWR.t6005 4.30165
R8331 VPWR.n2075 VPWR.t1369 4.30165
R8332 VPWR.n2071 VPWR.t5134 4.30165
R8333 VPWR.n2705 VPWR.t3572 4.30165
R8334 VPWR.n2703 VPWR.t1514 4.30165
R8335 VPWR.n2699 VPWR.t1518 4.30165
R8336 VPWR.n2695 VPWR.t2917 4.30165
R8337 VPWR.n2704 VPWR.t2364 4.30165
R8338 VPWR.n2067 VPWR.t4063 4.30165
R8339 VPWR.n2068 VPWR.t4650 4.30165
R8340 VPWR.n2072 VPWR.t967 4.30165
R8341 VPWR.n2078 VPWR.t5128 4.30165
R8342 VPWR.n463 VPWR.t2827 4.30165
R8343 VPWR.n464 VPWR.t2829 4.30165
R8344 VPWR.n468 VPWR.t1640 4.30165
R8345 VPWR.n474 VPWR.t3115 4.30165
R8346 VPWR.n478 VPWR.t4145 4.30165
R8347 VPWR.n482 VPWR.t6163 4.30165
R8348 VPWR.n486 VPWR.t507 4.30165
R8349 VPWR.n495 VPWR.t1732 4.30165
R8350 VPWR.n506 VPWR.t4722 4.30165
R8351 VPWR.n505 VPWR.t5340 4.30165
R8352 VPWR.n500 VPWR.t3337 4.30165
R8353 VPWR.n457 VPWR.t5608 4.30165
R8354 VPWR.n1879 VPWR.t1709 4.30165
R8355 VPWR.n1879 VPWR.t2605 4.30165
R8356 VPWR.n1878 VPWR.t2601 4.30165
R8357 VPWR.n1872 VPWR.t5177 4.30165
R8358 VPWR.n1873 VPWR.t3423 4.30165
R8359 VPWR.n503 VPWR.t3989 4.30165
R8360 VPWR.n504 VPWR.t734 4.30165
R8361 VPWR.n496 VPWR.t1728 4.30165
R8362 VPWR.n492 VPWR.t2870 4.30165
R8363 VPWR.n489 VPWR.t4499 4.30165
R8364 VPWR.n487 VPWR.t5188 4.30165
R8365 VPWR.n483 VPWR.t509 4.30165
R8366 VPWR.n479 VPWR.t4607 4.30165
R8367 VPWR.n473 VPWR.t751 4.30165
R8368 VPWR.n469 VPWR.t1492 4.30165
R8369 VPWR.n462 VPWR.t6316 4.30165
R8370 VPWR.n1923 VPWR.t3463 4.30165
R8371 VPWR.n1920 VPWR.t309 4.30165
R8372 VPWR.n1917 VPWR.t3121 4.30165
R8373 VPWR.n1909 VPWR.t1768 4.30165
R8374 VPWR.n1897 VPWR.t3153 4.30165
R8375 VPWR.n1891 VPWR.t5826 4.30165
R8376 VPWR.n1890 VPWR.t2503 4.30165
R8377 VPWR.n451 VPWR.t2862 4.30165
R8378 VPWR.n450 VPWR.t2860 4.30165
R8379 VPWR.n444 VPWR.t3069 4.30165
R8380 VPWR.n444 VPWR.t3421 4.30165
R8381 VPWR.n448 VPWR.t5493 4.30165
R8382 VPWR.n449 VPWR.t5113 4.30165
R8383 VPWR.n1888 VPWR.t1489 4.30165
R8384 VPWR.n1889 VPWR.t4841 4.30165
R8385 VPWR.n1896 VPWR.t5785 4.30165
R8386 VPWR.n1898 VPWR.t5073 4.30165
R8387 VPWR.n1432 VPWR.t2440 4.29774
R8388 VPWR.n1419 VPWR.t836 4.29774
R8389 VPWR.n1007 VPWR.t7137 4.29774
R8390 VPWR.n993 VPWR.t4400 4.29774
R8391 VPWR.n1004 VPWR.t3218 4.29774
R8392 VPWR.n1015 VPWR.t3534 4.29774
R8393 VPWR.n1618 VPWR.t2049 4.29774
R8394 VPWR.n1422 VPWR.t4451 4.29774
R8395 VPWR.n1647 VPWR.t6304 4.29774
R8396 VPWR.n3332 VPWR.t613 4.29774
R8397 VPWR.n898 VPWR.t5806 4.29774
R8398 VPWR.n796 VPWR.t3374 4.29774
R8399 VPWR.n782 VPWR.t820 4.29774
R8400 VPWR.n3314 VPWR.t949 4.29774
R8401 VPWR.n3303 VPWR.t4007 4.29774
R8402 VPWR.n793 VPWR.t4108 4.29774
R8403 VPWR.n1680 VPWR.t2260 4.29774
R8404 VPWR.n134 VPWR.t3869 4.29774
R8405 VPWR.n3203 VPWR.t4204 4.29774
R8406 VPWR.n3192 VPWR.t5856 4.29774
R8407 VPWR.n3213 VPWR.t2784 4.29774
R8408 VPWR.n1798 VPWR.t2022 4.29774
R8409 VPWR.n672 VPWR.t5673 4.29774
R8410 VPWR.n1105 VPWR.t1295 4.29774
R8411 VPWR.n2835 VPWR.t2895 4.29774
R8412 VPWR.n2919 VPWR.t585 4.29774
R8413 VPWR.n2902 VPWR.t5704 4.29774
R8414 VPWR.n2908 VPWR.t6265 4.29774
R8415 VPWR.n2857 VPWR.t4172 4.29774
R8416 VPWR.n2788 VPWR.t5249 4.29774
R8417 VPWR.n1863 VPWR.t3252 4.29774
R8418 VPWR.n548 VPWR.t6036 4.29774
R8419 VPWR.n415 VPWR.t1908 4.29774
R8420 VPWR.n2948 VPWR.t1752 4.29774
R8421 VPWR.n414 VPWR.t1922 4.29774
R8422 VPWR.n426 VPWR.t4564 4.29774
R8423 VPWR.n1075 VPWR.t6142 4.28209
R8424 VPWR.n1052 VPWR.t1110 4.28209
R8425 VPWR.n1619 VPWR.t4965 4.28209
R8426 VPWR.n975 VPWR.t5019 4.28209
R8427 VPWR.n1630 VPWR.t4182 4.28209
R8428 VPWR.n3347 VPWR.t6047 4.28209
R8429 VPWR.n3292 VPWR.t404 4.28209
R8430 VPWR.n1478 VPWR.t4670 4.27035
R8431 VPWR.n1629 VPWR.t6691 4.27035
R8432 VPWR.n814 VPWR.t3004 4.27035
R8433 VPWR.n1729 VPWR.t6547 4.27035
R8434 VPWR.n1771 VPWR.t292 4.27035
R8435 VPWR.n695 VPWR.t6918 4.27035
R8436 VPWR.n1027 VPWR.t4672 3.91054
R8437 VPWR.n1061 VPWR.t6146 3.91054
R8438 VPWR.n1037 VPWR.t1106 3.91054
R8439 VPWR.n921 VPWR.t4961 3.91054
R8440 VPWR.n914 VPWR.t4186 3.91054
R8441 VPWR.n745 VPWR.t3006 3.91054
R8442 VPWR.n911 VPWR.t6705 3.7566
R8443 VPWR.n2644 VPWR.n2643 3.5285
R8444 VPWR.n3837 VPWR.n3 3.5285
R8445 VPWR.t5752 VPWR.t6410 3.52369
R8446 VPWR.t6099 VPWR.t6065 3.47272
R8447 VPWR.t6866 VPWR 3.47272
R8448 VPWR VPWR.t668 3.47272
R8449 VPWR.t6908 VPWR 3.47272
R8450 VPWR VPWR.t6729 3.47272
R8451 VPWR.t4690 VPWR.t6006 3.47272
R8452 VPWR VPWR.t5117 3.47272
R8453 VPWR VPWR.t6527 3.47272
R8454 VPWR VPWR.t6966 3.47272
R8455 VPWR VPWR.t6510 3.47272
R8456 VPWR VPWR.t2595 3.47272
R8457 VPWR.t5012 VPWR 3.47272
R8458 VPWR.t3348 VPWR 3.47272
R8459 VPWR VPWR.t3401 3.47272
R8460 VPWR.n1370 VPWR.t6794 3.40237
R8461 VPWR.n1370 VPWR.t7095 3.40237
R8462 VPWR.n761 VPWR.t6526 3.40237
R8463 VPWR.n761 VPWR.t3478 3.40237
R8464 VPWR.n124 VPWR.t4559 3.40237
R8465 VPWR.n124 VPWR.t6969 3.40237
R8466 VPWR.n2867 VPWR.t6827 3.40237
R8467 VPWR.n2867 VPWR.t3396 3.40237
R8468 VPWR.n2870 VPWR.t6956 3.40237
R8469 VPWR.n2870 VPWR.t6427 3.40237
R8470 VPWR.n542 VPWR.t3347 3.40237
R8471 VPWR.n542 VPWR.t6610 3.40237
R8472 VPWR.n1383 VPWR.n1367 3.28037
R8473 VPWR.n1382 VPWR.n1368 3.28037
R8474 VPWR.n968 VPWR.n961 3.28037
R8475 VPWR.n1754 VPWR.n706 3.28037
R8476 VPWR.n596 VPWR.n524 3.28037
R8477 VPWR.n829 VPWR.t3141 3.15624
R8478 VPWR.n713 VPWR.t274 3.07367
R8479 VPWR.n711 VPWR.t264 3.07367
R8480 VPWR.n709 VPWR.t256 3.07367
R8481 VPWR.n708 VPWR.t6843 3.07367
R8482 VPWR.n710 VPWR.t6839 3.07367
R8483 VPWR.n712 VPWR.t6837 3.07367
R8484 VPWR.n610 VPWR.t272 3.07367
R8485 VPWR.n609 VPWR.t248 3.07367
R8486 VPWR.n608 VPWR.t246 3.07367
R8487 VPWR.n1393 VPWR.t7063 3.03383
R8488 VPWR.n1393 VPWR.t6217 3.03383
R8489 VPWR.n625 VPWR.t3916 3.03383
R8490 VPWR.n625 VPWR.t2379 3.03383
R8491 VPWR.n539 VPWR.t6378 3.03383
R8492 VPWR.n539 VPWR.t961 3.03383
R8493 VPWR.n382 VPWR.t4801 3.03383
R8494 VPWR.n382 VPWR.t5154 3.03383
R8495 VPWR.n3331 VPWR.n111 2.96671
R8496 VPWR.n1678 VPWR.n738 2.96671
R8497 VPWR.n1104 VPWR.n1095 2.96671
R8498 VPWR.n644 VPWR.n635 2.96671
R8499 VPWR.n1381 VPWR.n1369 2.95895
R8500 VPWR.n816 VPWR.n740 2.95895
R8501 VPWR.n1742 VPWR.n716 2.95895
R8502 VPWR.n1837 VPWR.n607 2.95895
R8503 VPWR.n1102 VPWR.n1096 2.95895
R8504 VPWR.n1378 VPWR.n1371 2.95583
R8505 VPWR.n131 VPWR.n130 2.95583
R8506 VPWR.n3239 VPWR.n126 2.95583
R8507 VPWR.n2913 VPWR.n2868 2.95583
R8508 VPWR.n2912 VPWR.n2869 2.95583
R8509 VPWR.n550 VPWR.n543 2.95583
R8510 VPWR.n986 VPWR.n950 2.85289
R8511 VPWR.n1702 VPWR.n730 2.85289
R8512 VPWR.n1700 VPWR.n731 2.85289
R8513 VPWR.n1195 VPWR.n1174 2.85289
R8514 VPWR.n1187 VPWR.n1176 2.85289
R8515 VPWR.n1800 VPWR.n1781 2.85289
R8516 VPWR.n671 VPWR.n629 2.85289
R8517 VPWR.n549 VPWR.n544 2.85289
R8518 VPWR.n561 VPWR.n540 2.85289
R8519 VPWR.n2942 VPWR.n179 2.85289
R8520 VPWR.n396 VPWR.t2952 2.82433
R8521 VPWR.n746 VPWR.t6983 2.82302
R8522 VPWR.n971 VPWR.n959 2.79028
R8523 VPWR.n969 VPWR.n960 2.79028
R8524 VPWR.n3342 VPWR.n3340 2.79028
R8525 VPWR.n107 VPWR.n106 2.79028
R8526 VPWR.n3287 VPWR.n3266 2.79028
R8527 VPWR.n3285 VPWR.n3270 2.79028
R8528 VPWR.n1023 VPWR.t2114 2.73703
R8529 VPWR.n918 VPWR.t3230 2.73703
R8530 VPWR.n1603 VPWR.n1019 2.72094
R8531 VPWR.n1514 VPWR.n1020 2.72094
R8532 VPWR.n1615 VPWR.n925 2.72094
R8533 VPWR.n1016 VPWR.n930 2.72094
R8534 VPWR.n3377 VPWR.n103 2.72094
R8535 VPWR.n1626 VPWR.n919 2.72094
R8536 VPWR.n897 VPWR.n831 2.72094
R8537 VPWR.n872 VPWR.n849 2.72094
R8538 VPWR.n1677 VPWR.n739 2.72094
R8539 VPWR.n427 VPWR.n380 2.72094
R8540 VPWR.n418 VPWR.n383 2.72094
R8541 VPWR.n730 VPWR.t4836 2.63984
R8542 VPWR.n731 VPWR.t1592 2.63984
R8543 VPWR.n1174 VPWR.t5409 2.63984
R8544 VPWR.n1176 VPWR.t1584 2.63984
R8545 VPWR.n943 VPWR.t6773 2.61116
R8546 VPWR.n748 VPWR.t188 2.61116
R8547 VPWR.n851 VPWR.t7003 2.55888
R8548 VPWR.n1765 VPWR.t5591 2.55888
R8549 VPWR.n529 VPWR.t4993 2.55888
R8550 VPWR.n959 VPWR.t5017 2.51646
R8551 VPWR.n3340 VPWR.t6045 2.51646
R8552 VPWR.n3266 VPWR.t400 2.51646
R8553 VPWR.n959 VPWR.t1949 2.37087
R8554 VPWR.n3340 VPWR.t3672 2.37087
R8555 VPWR.n3266 VPWR.t1338 2.37087
R8556 VPWR.n851 VPWR.t5145 2.3374
R8557 VPWR.n1765 VPWR.t36 2.3374
R8558 VPWR.n529 VPWR.t3021 2.3374
R8559 VPWR.t4978 VPWR.t6909 2.31531
R8560 VPWR.n1399 VPWR.t5050 2.2755
R8561 VPWR.n1409 VPWR.t2162 2.2755
R8562 VPWR.n937 VPWR.t2284 2.2755
R8563 VPWR.n948 VPWR.t5219 2.2755
R8564 VPWR.n940 VPWR.t5052 2.2755
R8565 VPWR.n931 VPWR.t3530 2.2755
R8566 VPWR.n924 VPWR.t672 2.2755
R8567 VPWR.n1408 VPWR.t5480 2.2755
R8568 VPWR.n824 VPWR.t1652 2.2755
R8569 VPWR.n110 VPWR.t2520 2.2755
R8570 VPWR.n832 VPWR.t1012 2.2755
R8571 VPWR.n751 VPWR.t2960 2.2755
R8572 VPWR.n757 VPWR.t5463 2.2755
R8573 VPWR.n123 VPWR.t3659 2.2755
R8574 VPWR.n3259 VPWR.t5836 2.2755
R8575 VPWR.n752 VPWR.t4106 2.2755
R8576 VPWR.n737 VPWR.t2258 2.2755
R8577 VPWR.n135 VPWR.t5915 2.2755
R8578 VPWR.n145 VPWR.t463 2.2755
R8579 VPWR.n152 VPWR.t4072 2.2755
R8580 VPWR.n139 VPWR.t3163 2.2755
R8581 VPWR.n1784 VPWR.t1669 2.2755
R8582 VPWR.n630 VPWR.t688 2.2755
R8583 VPWR.n1094 VPWR.t2286 2.2755
R8584 VPWR.n186 VPWR.t5426 2.2755
R8585 VPWR.n2851 VPWR.t333 2.2755
R8586 VPWR.n2875 VPWR.t1332 2.2755
R8587 VPWR.n2871 VPWR.t1797 2.2755
R8588 VPWR.n2848 VPWR.t3207 2.2755
R8589 VPWR.n2750 VPWR.t1456 2.2755
R8590 VPWR.n515 VPWR.t878 2.2755
R8591 VPWR.n545 VPWR.t2241 2.2755
R8592 VPWR.n386 VPWR.t3082 2.2755
R8593 VPWR.n2943 VPWR.t4048 2.2755
R8594 VPWR.n387 VPWR.t2463 2.2755
R8595 VPWR.n379 VPWR.t2738 2.2755
R8596 VPWR.n1394 VPWR.t5585 2.25159
R8597 VPWR.n623 VPWR.t5629 2.25159
R8598 VPWR.n538 VPWR.t5824 2.25159
R8599 VPWR.n384 VPWR.t7100 2.25159
R8600 VPWR.n1027 VPWR.t11 2.22001
R8601 VPWR.n1061 VPWR.t7051 2.22001
R8602 VPWR.n1037 VPWR.t6344 2.22001
R8603 VPWR.n1411 VPWR.t6699 2.22001
R8604 VPWR.n1411 VPWR.t6701 2.22001
R8605 VPWR.n921 VPWR.t6520 2.22001
R8606 VPWR.n914 VPWR.t1691 2.22001
R8607 VPWR.n745 VPWR.t6743 2.22001
R8608 VPWR.n713 VPWR.t260 2.22001
R8609 VPWR.n711 VPWR.t262 2.22001
R8610 VPWR.n709 VPWR.t250 2.22001
R8611 VPWR.n708 VPWR.t6845 2.22001
R8612 VPWR.n710 VPWR.t6835 2.22001
R8613 VPWR.n712 VPWR.t6833 2.22001
R8614 VPWR.n610 VPWR.t268 2.22001
R8615 VPWR.n609 VPWR.t254 2.22001
R8616 VPWR.n608 VPWR.t252 2.22001
R8617 VPWR.n835 VPWR.t2349 2.15435
R8618 VPWR.n837 VPWR.t6532 2.15435
R8619 VPWR.n837 VPWR.t6539 2.15435
R8620 VPWR.n838 VPWR.t2362 2.15435
R8621 VPWR.n839 VPWR.t6534 2.15435
R8622 VPWR.n839 VPWR.t3475 2.15435
R8623 VPWR.n841 VPWR.t6965 2.15435
R8624 VPWR.n841 VPWR.t6974 2.15435
R8625 VPWR.n842 VPWR.t3485 2.15435
R8626 VPWR.n842 VPWR.t3480 2.15435
R8627 VPWR.n843 VPWR.t6978 2.15435
R8628 VPWR.n843 VPWR.t6976 2.15435
R8629 VPWR.n856 VPWR.t6409 2.15435
R8630 VPWR.n857 VPWR.t6847 2.15435
R8631 VPWR.n857 VPWR.t6853 2.15435
R8632 VPWR.n118 VPWR.t6413 2.15435
R8633 VPWR.n117 VPWR.t6849 2.15435
R8634 VPWR.n117 VPWR.t4086 2.15435
R8635 VPWR.n116 VPWR.t2561 2.15435
R8636 VPWR.n116 VPWR.t2558 2.15435
R8637 VPWR.n113 VPWR.t4088 2.15435
R8638 VPWR.n113 VPWR.t4083 2.15435
R8639 VPWR.n112 VPWR.t2563 2.15435
R8640 VPWR.n112 VPWR.t2556 2.15435
R8641 VPWR.n1780 VPWR.t6289 2.15435
R8642 VPWR.n1780 VPWR.t2165 2.15435
R8643 VPWR.n627 VPWR.t6605 2.15435
R8644 VPWR.n627 VPWR.t6594 2.15435
R8645 VPWR.n518 VPWR.t4793 2.15435
R8646 VPWR.n518 VPWR.t5006 2.15435
R8647 VPWR.n519 VPWR.t4325 2.15435
R8648 VPWR.n519 VPWR.t3300 2.15435
R8649 VPWR.n521 VPWR.t3296 2.15435
R8650 VPWR.n521 VPWR.t4327 2.15435
R8651 VPWR.n522 VPWR.t5000 2.15435
R8652 VPWR.n522 VPWR.t4805 2.15435
R8653 VPWR.n537 VPWR.t5121 2.15435
R8654 VPWR.n537 VPWR.t6891 2.15435
R8655 VPWR.n1396 VPWR.t6751 2.10455
R8656 VPWR.n1396 VPWR.t6948 2.10455
R8657 VPWR.n1401 VPWR.t6759 2.10455
R8658 VPWR.n1401 VPWR.t7061 2.10455
R8659 VPWR.n942 VPWR.t6368 2.10455
R8660 VPWR.n942 VPWR.t6483 2.10455
R8661 VPWR.n951 VPWR.t159 2.10455
R8662 VPWR.n951 VPWR.t6481 2.10455
R8663 VPWR.n102 VPWR.t139 2.10455
R8664 VPWR.n102 VPWR.t6491 2.10455
R8665 VPWR.n944 VPWR.t6868 2.10455
R8666 VPWR.n944 VPWR.t6479 2.10455
R8667 VPWR.n936 VPWR.t97 2.10455
R8668 VPWR.n936 VPWR.t6487 2.10455
R8669 VPWR.n927 VPWR.t7057 2.10455
R8670 VPWR.n927 VPWR.t6469 2.10455
R8671 VPWR.n1412 VPWR.t7042 2.10455
R8672 VPWR.n1412 VPWR.t6493 2.10455
R8673 VPWR.n828 VPWR.t7097 2.10455
R8674 VPWR.n828 VPWR.t6499 2.10455
R8675 VPWR.n3356 VPWR.t6906 2.10455
R8676 VPWR.n3356 VPWR.t6495 2.10455
R8677 VPWR.n3338 VPWR.t103 2.10455
R8678 VPWR.n3338 VPWR.t6477 2.10455
R8679 VPWR.n836 VPWR.t6614 2.10455
R8680 VPWR.n836 VPWR.t6648 2.10455
R8681 VPWR.n754 VPWR.t144 2.10455
R8682 VPWR.n754 VPWR.t6654 2.10455
R8683 VPWR.n759 VPWR.t223 2.10455
R8684 VPWR.n759 VPWR.t6652 2.10455
R8685 VPWR.n3258 VPWR.t6339 2.10455
R8686 VPWR.n3258 VPWR.t6485 2.10455
R8687 VPWR.n3272 VPWR.t6384 2.10455
R8688 VPWR.n3272 VPWR.t6467 2.10455
R8689 VPWR.n3264 VPWR.t7007 2.10455
R8690 VPWR.n3264 VPWR.t6473 2.10455
R8691 VPWR.n747 VPWR.t6767 2.10455
R8692 VPWR.n747 VPWR.t176 2.10455
R8693 VPWR.n734 VPWR.t6755 2.10455
R8694 VPWR.n734 VPWR.t6370 2.10455
R8695 VPWR.n138 VPWR.t38 2.10455
R8696 VPWR.n138 VPWR.t6489 2.10455
R8697 VPWR.n148 VPWR.t6740 2.10455
R8698 VPWR.n148 VPWR.t6475 2.10455
R8699 VPWR.n154 VPWR.t7028 2.10455
R8700 VPWR.n154 VPWR.t6465 2.10455
R8701 VPWR.n144 VPWR.t6389 2.10455
R8702 VPWR.n144 VPWR.t6471 2.10455
R8703 VPWR.n1786 VPWR.t6397 2.10455
R8704 VPWR.n1786 VPWR.t6664 2.10455
R8705 VPWR.n633 VPWR.t155 2.10455
R8706 VPWR.n633 VPWR.t6660 2.10455
R8707 VPWR.n1089 VPWR.t6747 2.10455
R8708 VPWR.n1089 VPWR.t26 2.10455
R8709 VPWR.n1939 VPWR.t6757 2.10455
R8710 VPWR.n1939 VPWR.t128 2.10455
R8711 VPWR.n2847 VPWR.t6650 2.10455
R8712 VPWR.n2847 VPWR.t6461 2.10455
R8713 VPWR.n2878 VPWR.t92 2.10455
R8714 VPWR.n2878 VPWR.t6646 2.10455
R8715 VPWR.n2876 VPWR.t6944 2.10455
R8716 VPWR.n2876 VPWR.t6656 2.10455
R8717 VPWR.n185 VPWR.t7045 2.10455
R8718 VPWR.n185 VPWR.t6662 2.10455
R8719 VPWR.n2747 VPWR.t6644 2.10455
R8720 VPWR.n2747 VPWR.t164 2.10455
R8721 VPWR.n513 VPWR.t6745 2.10455
R8722 VPWR.n513 VPWR.t6597 2.10455
R8723 VPWR.n174 VPWR.t99 2.10455
R8724 VPWR.n174 VPWR.t6666 2.10455
R8725 VPWR.n390 VPWR.t200 2.10455
R8726 VPWR.n390 VPWR.t6668 2.10455
R8727 VPWR.n2954 VPWR.t51 2.10455
R8728 VPWR.n2954 VPWR.t6658 2.10455
R8729 VPWR.n391 VPWR.t7033 2.10455
R8730 VPWR.n391 VPWR.t6642 2.10455
R8731 VPWR.n375 VPWR.t6763 2.10455
R8732 VPWR.n375 VPWR.t6416 2.10455
R8733 VPWR.n605 VPWR.t3304 2.08822
R8734 VPWR.n701 VPWR.t2458 2.07457
R8735 VPWR.n606 VPWR.t6712 2.07457
R8736 VPWR.n1019 VPWR.t1205 2.06607
R8737 VPWR.n1019 VPWR.t1203 2.06607
R8738 VPWR.n1020 VPWR.t3665 2.06607
R8739 VPWR.n1020 VPWR.t3663 2.06607
R8740 VPWR.n1028 VPWR.t4674 2.06607
R8741 VPWR.n1060 VPWR.t6140 2.06607
R8742 VPWR.n1039 VPWR.t1112 2.06607
R8743 VPWR.n922 VPWR.t4959 2.06607
R8744 VPWR.n925 VPWR.t6334 2.06607
R8745 VPWR.n925 VPWR.t6336 2.06607
R8746 VPWR.n930 VPWR.t150 2.06607
R8747 VPWR.n930 VPWR.t152 2.06607
R8748 VPWR.n919 VPWR.t5922 2.06607
R8749 VPWR.n919 VPWR.t5920 2.06607
R8750 VPWR.n916 VPWR.t4188 2.06607
R8751 VPWR.n830 VPWR.t3143 2.06607
R8752 VPWR.n849 VPWR.t2034 2.06607
R8753 VPWR.n849 VPWR.t2032 2.06607
R8754 VPWR.n744 VPWR.t3002 2.06607
R8755 VPWR.n723 VPWR.t6555 2.06607
R8756 VPWR.n722 VPWR.t6573 2.06607
R8757 VPWR.n721 VPWR.t6565 2.06607
R8758 VPWR.n720 VPWR.t6561 2.06607
R8759 VPWR.n719 VPWR.t6559 2.06607
R8760 VPWR.n718 VPWR.t6551 2.06607
R8761 VPWR.n717 VPWR.t6549 2.06607
R8762 VPWR.n1764 VPWR.t290 2.06607
R8763 VPWR.n1762 VPWR.t236 2.06607
R8764 VPWR.n1761 VPWR.t278 2.06607
R8765 VPWR.n702 VPWR.t280 2.06607
R8766 VPWR.n703 VPWR.t282 2.06607
R8767 VPWR.n704 VPWR.t284 2.06607
R8768 VPWR.n705 VPWR.t238 2.06607
R8769 VPWR.n622 VPWR.t6926 2.06607
R8770 VPWR.n620 VPWR.t6922 2.06607
R8771 VPWR.n619 VPWR.t6934 2.06607
R8772 VPWR.n617 VPWR.t6936 2.06607
R8773 VPWR.n616 VPWR.t6914 2.06607
R8774 VPWR.n615 VPWR.t6916 2.06607
R8775 VPWR.n613 VPWR.t6928 2.06607
R8776 VPWR.n943 VPWR.t888 2.03739
R8777 VPWR.n748 VPWR.t1620 2.03739
R8778 VPWR.n960 VPWR.t1947 1.92643
R8779 VPWR.n106 VPWR.t3670 1.92643
R8780 VPWR.n3270 VPWR.t1340 1.92643
R8781 VPWR.n958 VPWR.t414 1.84822
R8782 VPWR.n958 VPWR.t5671 1.84822
R8783 VPWR.n1372 VPWR.t315 1.84822
R8784 VPWR.n1372 VPWR.t3755 1.84822
R8785 VPWR.n847 VPWR.t794 1.84822
R8786 VPWR.n847 VPWR.t798 1.84822
R8787 VPWR.n848 VPWR.t7001 1.84822
R8788 VPWR.n848 VPWR.t6997 1.84822
R8789 VPWR.n850 VPWR.t796 1.84822
R8790 VPWR.n850 VPWR.t800 1.84822
R8791 VPWR.n821 VPWR.t7036 1.84822
R8792 VPWR.n821 VPWR.t4223 1.84822
R8793 VPWR.n820 VPWR.t4221 1.84822
R8794 VPWR.n820 VPWR.t6502 1.84822
R8795 VPWR.n129 VPWR.t6541 1.84822
R8796 VPWR.n129 VPWR.t2358 1.84822
R8797 VPWR.n127 VPWR.t2351 1.84822
R8798 VPWR.n127 VPWR.t6530 1.84822
R8799 VPWR.n125 VPWR.t7110 1.84822
R8800 VPWR.n125 VPWR.t6971 1.84822
R8801 VPWR.n3245 VPWR.t4212 1.84822
R8802 VPWR.n3245 VPWR.t174 1.84822
R8803 VPWR.n3244 VPWR.t168 1.84822
R8804 VPWR.n3244 VPWR.t4208 1.84822
R8805 VPWR.n1766 VPWR.t2546 1.84822
R8806 VPWR.n1766 VPWR.t2538 1.84822
R8807 VPWR.n698 VPWR.t5595 1.84822
R8808 VPWR.n698 VPWR.t5597 1.84822
R8809 VPWR.n700 VPWR.t2544 1.84822
R8810 VPWR.n700 VPWR.t2540 1.84822
R8811 VPWR.n1097 VPWR.t6807 1.84822
R8812 VPWR.n1097 VPWR.t1267 1.84822
R8813 VPWR.n626 VPWR.t4820 1.84822
R8814 VPWR.n626 VPWR.t4232 1.84822
R8815 VPWR.n531 VPWR.t232 1.84822
R8816 VPWR.n531 VPWR.t230 1.84822
R8817 VPWR.n532 VPWR.t4989 1.84822
R8818 VPWR.n532 VPWR.t4991 1.84822
R8819 VPWR.n533 VPWR.t234 1.84822
R8820 VPWR.n533 VPWR.t228 1.84822
R8821 VPWR.n536 VPWR.t6824 1.84822
R8822 VPWR.n536 VPWR.t6893 1.84822
R8823 VPWR.n520 VPWR.t4321 1.84822
R8824 VPWR.n520 VPWR.t3298 1.84822
R8825 VPWR.n397 VPWR.t6708 1.84822
R8826 VPWR.n397 VPWR.t6805 1.84822
R8827 VPWR.n2501 VPWR.n264 1.7645
R8828 VPWR.n2601 VPWR.n259 1.7645
R8829 VPWR.n1063 VPWR.t5653 1.75837
R8830 VPWR.n1062 VPWR.t2530 1.75837
R8831 VPWR.n956 VPWR.t1361 1.75837
R8832 VPWR.n1023 VPWR.t89 1.73383
R8833 VPWR.n918 VPWR.t5930 1.73383
R8834 VPWR.n103 VPWR.t4390 1.72898
R8835 VPWR.n831 VPWR.t4050 1.72898
R8836 VPWR.n739 VPWR.t2478 1.72898
R8837 VPWR.n380 VPWR.t469 1.72898
R8838 VPWR.n383 VPWR.t3611 1.72898
R8839 VPWR.n605 VPWR.t3306 1.7198
R8840 VPWR.n746 VPWR.t775 1.68569
R8841 VPWR.n396 VPWR.t4700 1.68569
R8842 VPWR.n911 VPWR.t6695 1.67844
R8843 VPWR.n852 VPWR.t5143 1.6626
R8844 VPWR.n852 VPWR.t5139 1.6626
R8845 VPWR.n1763 VPWR.t32 1.6626
R8846 VPWR.n1763 VPWR.t34 1.6626
R8847 VPWR.n527 VPWR.t3017 1.6626
R8848 VPWR.n527 VPWR.t3023 1.6626
R8849 VPWR.n1021 VPWR.t6228 1.66185
R8850 VPWR.n1034 VPWR.t3410 1.66185
R8851 VPWR.n840 VPWR.t2086 1.66185
R8852 VPWR.n147 VPWR.t5708 1.66185
R8853 VPWR.n2872 VPWR.t2036 1.65985
R8854 VPWR.n602 VPWR.t6803 1.61112
R8855 VPWR.n602 VPWR.t6796 1.61112
R8856 VPWR.n526 VPWR.t6798 1.61112
R8857 VPWR.n526 VPWR.t6811 1.61112
R8858 VPWR.n950 VPWR.t5063 1.5575
R8859 VPWR.n1781 VPWR.t2067 1.5575
R8860 VPWR.n629 VPWR.t3224 1.5575
R8861 VPWR.n544 VPWR.t3935 1.5575
R8862 VPWR.n540 VPWR.t5147 1.5575
R8863 VPWR.n179 VPWR.t2002 1.5575
R8864 VPWR.n715 VPWR.t6571 1.52029
R8865 VPWR.n707 VPWR.t240 1.52029
R8866 VPWR.n611 VPWR.t6930 1.52029
R8867 VPWR.n855 VPWR.t3578 1.51717
R8868 VPWR.n855 VPWR.t3583 1.51717
R8869 VPWR.n854 VPWR.t3580 1.51717
R8870 VPWR.n854 VPWR.t3576 1.51717
R8871 VPWR.n1387 VPWR.t5269 1.49844
R8872 VPWR.n1387 VPWR.t5810 1.49844
R8873 VPWR.n1395 VPWR.t1035 1.49844
R8874 VPWR.n1395 VPWR.t2609 1.49844
R8875 VPWR.n1036 VPWR.t4871 1.49844
R8876 VPWR.n1036 VPWR.t6880 1.49844
R8877 VPWR.n1277 VPWR.t1215 1.49844
R8878 VPWR.n1277 VPWR.t6872 1.49844
R8879 VPWR.n823 VPWR.t3730 1.49844
R8880 VPWR.n823 VPWR.t212 1.49844
R8881 VPWR.n701 VPWR.t2456 1.49844
R8882 VPWR.n606 VPWR.t6714 1.49844
R8883 VPWR.n1028 VPWR.t4676 1.4923
R8884 VPWR.n1060 VPWR.t6144 1.4923
R8885 VPWR.n1039 VPWR.t1108 1.4923
R8886 VPWR.n1390 VPWR.t4599 1.4923
R8887 VPWR.n1390 VPWR.t4605 1.4923
R8888 VPWR.n913 VPWR.t6697 1.4923
R8889 VPWR.n913 VPWR.t6689 1.4923
R8890 VPWR.n915 VPWR.t6683 1.4923
R8891 VPWR.n915 VPWR.t6687 1.4923
R8892 VPWR.n917 VPWR.t6693 1.4923
R8893 VPWR.n917 VPWR.t6685 1.4923
R8894 VPWR.n922 VPWR.t4963 1.4923
R8895 VPWR.n957 VPWR.t5015 1.4923
R8896 VPWR.n957 VPWR.t5023 1.4923
R8897 VPWR.n916 VPWR.t4184 1.4923
R8898 VPWR.n1391 VPWR.t6277 1.4923
R8899 VPWR.n1391 VPWR.t6275 1.4923
R8900 VPWR.n1388 VPWR.t2653 1.4923
R8901 VPWR.n1388 VPWR.t2660 1.4923
R8902 VPWR.n1280 VPWR.t1431 1.4923
R8903 VPWR.n1280 VPWR.t1429 1.4923
R8904 VPWR.n1279 VPWR.t5201 1.4923
R8905 VPWR.n1279 VPWR.t5204 1.4923
R8906 VPWR.n829 VPWR.t3599 1.4923
R8907 VPWR.n830 VPWR.t3139 1.4923
R8908 VPWR.n3339 VPWR.t6041 1.4923
R8909 VPWR.n3339 VPWR.t6049 1.4923
R8910 VPWR.n730 VPWR.t5741 1.4923
R8911 VPWR.n732 VPWR.t3881 1.4923
R8912 VPWR.n732 VPWR.t7024 1.4923
R8913 VPWR.n744 VPWR.t3008 1.4923
R8914 VPWR.n3265 VPWR.t402 1.4923
R8915 VPWR.n3265 VPWR.t406 1.4923
R8916 VPWR.n733 VPWR.t4436 1.4923
R8917 VPWR.n733 VPWR.t7009 1.4923
R8918 VPWR.n731 VPWR.t337 1.4923
R8919 VPWR.n1173 VPWR.t7026 1.4923
R8920 VPWR.n1173 VPWR.t1862 1.4923
R8921 VPWR.n1174 VPWR.t2594 1.4923
R8922 VPWR.n1176 VPWR.t2730 1.4923
R8923 VPWR.n1177 VPWR.t4160 1.4923
R8924 VPWR.n1177 VPWR.t7019 1.4923
R8925 VPWR.n723 VPWR.t6553 1.4923
R8926 VPWR.n722 VPWR.t6569 1.4923
R8927 VPWR.n721 VPWR.t6567 1.4923
R8928 VPWR.n720 VPWR.t6563 1.4923
R8929 VPWR.n719 VPWR.t6557 1.4923
R8930 VPWR.n718 VPWR.t6545 1.4923
R8931 VPWR.n717 VPWR.t6543 1.4923
R8932 VPWR.n1764 VPWR.t294 1.4923
R8933 VPWR.n1762 VPWR.t242 1.4923
R8934 VPWR.n1761 VPWR.t276 1.4923
R8935 VPWR.n702 VPWR.t286 1.4923
R8936 VPWR.n703 VPWR.t288 1.4923
R8937 VPWR.n704 VPWR.t296 1.4923
R8938 VPWR.n705 VPWR.t298 1.4923
R8939 VPWR.n622 VPWR.t6920 1.4923
R8940 VPWR.n620 VPWR.t6938 1.4923
R8941 VPWR.n619 VPWR.t6940 1.4923
R8942 VPWR.n617 VPWR.t6910 1.4923
R8943 VPWR.n616 VPWR.t6912 1.4923
R8944 VPWR.n615 VPWR.t6924 1.4923
R8945 VPWR.n613 VPWR.t6932 1.4923
R8946 VPWR.n1371 VPWR.t5 1.44083
R8947 VPWR.n111 VPWR.t2228 1.44083
R8948 VPWR.n738 VPWR.t4126 1.44083
R8949 VPWR.n130 VPWR.t3183 1.44083
R8950 VPWR.n126 VPWR.t1084 1.44083
R8951 VPWR.n1095 VPWR.t5394 1.44083
R8952 VPWR.n635 VPWR.t3849 1.44083
R8953 VPWR.n2868 VPWR.t6030 1.44083
R8954 VPWR.n2869 VPWR.t899 1.44083
R8955 VPWR.n543 VPWR.t2393 1.44083
R8956 VPWR.n1369 VPWR.t971 1.43493
R8957 VPWR.n740 VPWR.t1022 1.43493
R8958 VPWR.n716 VPWR.t1795 1.43493
R8959 VPWR.n607 VPWR.t850 1.43493
R8960 VPWR.n1096 VPWR.t441 1.43493
R8961 VPWR.n1367 VPWR.t6082 1.2628
R8962 VPWR.n1368 VPWR.t5123 1.2628
R8963 VPWR.n961 VPWR.t6066 1.2628
R8964 VPWR.n706 VPWR.t2806 1.2628
R8965 VPWR.n524 VPWR.t1168 1.2628
R8966 VPWR VPWR.t6577 1.15791
R8967 VPWR.t6990 VPWR.t4201 1.15791
R8968 VPWR.n964 VPWR.n963 1.07151
R8969 VPWR.n953 VPWR.n952 1.07151
R8970 VPWR.n1403 VPWR.n1402 1.07151
R8971 VPWR.n827 VPWR.n826 1.07151
R8972 VPWR.n3261 VPWR.n3260 1.07151
R8973 VPWR.n150 VPWR.n149 1.07151
R8974 VPWR.n946 VPWR.n945 0.993319
R8975 VPWR.n934 VPWR.n933 0.993319
R8976 VPWR.n1405 VPWR.n1404 0.993319
R8977 VPWR.n845 VPWR.n844 0.993319
R8978 VPWR.n3268 VPWR.n3267 0.993319
R8979 VPWR.n742 VPWR.n741 0.993319
R8980 VPWR.n1840 VPWR.n1839 0.77675
R8981 VPWR.n1058 VPWR.n1057 0.7625
R8982 VPWR.n1068 VPWR.n1067 0.7625
R8983 VPWR.n1485 VPWR.n1484 0.7625
R8984 VPWR.n1472 VPWR.n1032 0.75725
R8985 VPWR.n1067 VPWR.n1032 0.668
R8986 VPWR.n1514 VPWR.n1513 0.665
R8987 VPWR.n1603 VPWR.n1602 0.665
R8988 VPWR.n2855 VPWR.n2854 0.6455
R8989 VPWR.n2853 VPWR.n2852 0.6455
R8990 VPWR.n393 VPWR.n392 0.639539
R8991 VPWR.n1515 VPWR 0.635
R8992 VPWR.n1604 VPWR 0.635
R8993 VPWR.n429 VPWR 0.5885
R8994 VPWR.n412 VPWR.n411 0.5735
R8995 VPWR.n1511 VPWR.n1510 0.5405
R8996 VPWR.n2906 VPWR.n2905 0.5405
R8997 VPWR.n3357 VPWR.t3448 0.539645
R8998 VPWR.n155 VPWR.t2956 0.539645
R8999 VPWR.n1091 VPWR.t6069 0.536735
R9000 VPWR VPWR.n1070 0.5015
R9001 VPWR.n410 VPWR.n409 0.4895
R9002 VPWR VPWR.n3201 0.48725
R9003 VPWR.n1002 VPWR.n1001 0.4745
R9004 VPWR.n795 VPWR.n794 0.4625
R9005 VPWR.n1484 VPWR 0.46025
R9006 VPWR.n1616 VPWR.n1615 0.4535
R9007 VPWR VPWR.n864 0.4535
R9008 VPWR VPWR.n998 0.44675
R9009 VPWR.n896 VPWR 0.44225
R9010 VPWR.n3215 VPWR.n3214 0.4415
R9011 VPWR.n1346 VPWR.n1345 0.4415
R9012 VPWR.n1345 VPWR.n1265 0.4415
R9013 VPWR.n1265 VPWR.n1216 0.4415
R9014 VPWR.n1216 VPWR.n1158 0.4415
R9015 VPWR.n1158 VPWR.n359 0.4415
R9016 VPWR.n1925 VPWR.n359 0.4415
R9017 VPWR.n2005 VPWR.n1925 0.4415
R9018 VPWR.n2054 VPWR.n2005 0.4415
R9019 VPWR.n2099 VPWR.n2054 0.4415
R9020 VPWR.n2100 VPWR.n2099 0.4415
R9021 VPWR.n2100 VPWR.n273 0.4415
R9022 VPWR.n2316 VPWR.n273 0.4415
R9023 VPWR.n2383 VPWR.n2316 0.4415
R9024 VPWR.n2394 VPWR.n2383 0.4415
R9025 VPWR.n2405 VPWR.n2394 0.4415
R9026 VPWR.n2416 VPWR.n2405 0.4415
R9027 VPWR.n2456 VPWR.n2416 0.4415
R9028 VPWR.n2456 VPWR.n2455 0.4415
R9029 VPWR.n1471 VPWR.n727 0.4415
R9030 VPWR.n1708 VPWR.n727 0.4415
R9031 VPWR.n1709 VPWR.n1708 0.4415
R9032 VPWR.n1709 VPWR.n456 0.4415
R9033 VPWR.n1882 VPWR.n456 0.4415
R9034 VPWR.n1883 VPWR.n1882 0.4415
R9035 VPWR.n1883 VPWR.n195 0.4415
R9036 VPWR.n2709 VPWR.n195 0.4415
R9037 VPWR.n2709 VPWR.n2708 0.4415
R9038 VPWR.n2708 VPWR.n196 0.4415
R9039 VPWR.n2276 VPWR.n196 0.4415
R9040 VPWR.n2277 VPWR.n2276 0.4415
R9041 VPWR.n2277 VPWR.n264 0.4415
R9042 VPWR.n2502 VPWR.n2501 0.4415
R9043 VPWR.n1674 VPWR.n817 0.4415
R9044 VPWR.n1675 VPWR.n1674 0.4415
R9045 VPWR.n1675 VPWR.n601 0.4415
R9046 VPWR.n1845 VPWR.n601 0.4415
R9047 VPWR.n1846 VPWR.n1845 0.4415
R9048 VPWR.n1846 VPWR.n190 0.4415
R9049 VPWR.n2830 VPWR.n190 0.4415
R9050 VPWR.n2830 VPWR.n2829 0.4415
R9051 VPWR.n2829 VPWR.n191 0.4415
R9052 VPWR.n2185 VPWR.n191 0.4415
R9053 VPWR.n2238 VPWR.n2185 0.4415
R9054 VPWR.n2238 VPWR.n2237 0.4415
R9055 VPWR.n2237 VPWR.n259 0.4415
R9056 VPWR.n2601 VPWR.n2600 0.4415
R9057 VPWR.n1641 VPWR.n1640 0.4415
R9058 VPWR.n1641 VPWR.n697 0.4415
R9059 VPWR.n1816 VPWR.n697 0.4415
R9060 VPWR.n1817 VPWR.n1816 0.4415
R9061 VPWR.n1817 VPWR.n182 0.4415
R9062 VPWR.n2922 VPWR.n182 0.4415
R9063 VPWR.n2922 VPWR.n2921 0.4415
R9064 VPWR.n2921 VPWR.n183 0.4415
R9065 VPWR.n2644 VPWR.n183 0.4415
R9066 VPWR.n2643 VPWR.n255 0.4415
R9067 VPWR.n1606 VPWR.n132 0.4415
R9068 VPWR.n3223 VPWR.n132 0.4415
R9069 VPWR.n3223 VPWR.n3222 0.4415
R9070 VPWR.n3222 VPWR.n133 0.4415
R9071 VPWR.n3022 VPWR.n133 0.4415
R9072 VPWR.n3022 VPWR.n3021 0.4415
R9073 VPWR.n3021 VPWR.n178 0.4415
R9074 VPWR.n2762 VPWR.n178 0.4415
R9075 VPWR.n2762 VPWR.n3 0.4415
R9076 VPWR.n3838 VPWR.n3837 0.4415
R9077 VPWR.n3318 VPWR.n120 0.4415
R9078 VPWR.n3318 VPWR.n3317 0.4415
R9079 VPWR.n3317 VPWR.n121 0.4415
R9080 VPWR.n3108 VPWR.n121 0.4415
R9081 VPWR.n3108 VPWR.n3107 0.4415
R9082 VPWR.n3107 VPWR.n8 0.4415
R9083 VPWR.n3816 VPWR.n3815 0.4415
R9084 VPWR.n3374 VPWR.n3373 0.4415
R9085 VPWR.n3373 VPWR.n105 0.4415
R9086 VPWR.n3160 VPWR.n105 0.4415
R9087 VPWR.n3160 VPWR.n3159 0.4415
R9088 VPWR.n3159 VPWR.n170 0.4415
R9089 VPWR.n170 VPWR.n37 0.4415
R9090 VPWR.n3777 VPWR.n3776 0.4415
R9091 VPWR.n3458 VPWR.n3443 0.4415
R9092 VPWR.n3473 VPWR.n3458 0.4415
R9093 VPWR.n3488 VPWR.n3473 0.4415
R9094 VPWR.n3503 VPWR.n3488 0.4415
R9095 VPWR.n3518 VPWR.n3503 0.4415
R9096 VPWR.n3533 VPWR.n3518 0.4415
R9097 VPWR.n3548 VPWR.n3533 0.4415
R9098 VPWR.n3563 VPWR.n3548 0.4415
R9099 VPWR.n3578 VPWR.n3563 0.4415
R9100 VPWR.n3593 VPWR.n3578 0.4415
R9101 VPWR.n3608 VPWR.n3593 0.4415
R9102 VPWR.n3623 VPWR.n3608 0.4415
R9103 VPWR.n3638 VPWR.n3623 0.4415
R9104 VPWR.n3653 VPWR.n3638 0.4415
R9105 VPWR.n3668 VPWR.n3653 0.4415
R9106 VPWR.n3683 VPWR.n3668 0.4415
R9107 VPWR.n3715 VPWR.n3683 0.4415
R9108 VPWR.n3716 VPWR.n3715 0.4415
R9109 VPWR.n3755 VPWR.n3754 0.4415
R9110 VPWR VPWR.n898 0.4325
R9111 VPWR.n582 VPWR 0.422
R9112 VPWR VPWR.n3193 0.4175
R9113 VPWR VPWR.n866 0.3935
R9114 VPWR VPWR.n3207 0.3905
R9115 VPWR.n1057 VPWR 0.377
R9116 VPWR.n1614 VPWR.n1613 0.377
R9117 VPWR VPWR.n1447 0.3755
R9118 VPWR.n1011 VPWR 0.37325
R9119 VPWR.n3310 VPWR 0.37325
R9120 VPWR VPWR.n1444 0.37175
R9121 VPWR.n3451 VPWR 0.3665
R9122 VPWR.n3466 VPWR 0.3665
R9123 VPWR.n3481 VPWR 0.3665
R9124 VPWR.n3496 VPWR 0.3665
R9125 VPWR.n3511 VPWR 0.3665
R9126 VPWR.n3526 VPWR 0.3665
R9127 VPWR.n3541 VPWR 0.3665
R9128 VPWR.n3556 VPWR 0.3665
R9129 VPWR.n3571 VPWR 0.3665
R9130 VPWR.n3586 VPWR 0.3665
R9131 VPWR.n3601 VPWR 0.3665
R9132 VPWR.n3616 VPWR 0.3665
R9133 VPWR.n3631 VPWR 0.3665
R9134 VPWR.n3646 VPWR 0.3665
R9135 VPWR.n3661 VPWR 0.3665
R9136 VPWR.n3676 VPWR 0.3665
R9137 VPWR VPWR.n1541 0.3665
R9138 VPWR.n3436 VPWR 0.3665
R9139 VPWR.n3359 VPWR 0.3665
R9140 VPWR VPWR.n1234 0.3665
R9141 VPWR.n3274 VPWR 0.3665
R9142 VPWR.n157 VPWR 0.3665
R9143 VPWR.n3145 VPWR 0.3665
R9144 VPWR.n2881 VPWR 0.3665
R9145 VPWR.n2168 VPWR 0.3665
R9146 VPWR.n332 VPWR 0.3665
R9147 VPWR.n2389 VPWR 0.3665
R9148 VPWR.n2400 VPWR 0.3665
R9149 VPWR.n2411 VPWR 0.3665
R9150 VPWR.n2220 VPWR 0.3665
R9151 VPWR.n2331 VPWR 0.3665
R9152 VPWR.n2751 VPWR 0.3665
R9153 VPWR.n208 VPWR 0.3665
R9154 VPWR.n3056 VPWR 0.3665
R9155 VPWR.n2960 VPWR 0.3665
R9156 VPWR.n3708 VPWR 0.3665
R9157 VPWR.n89 VPWR 0.3665
R9158 VPWR VPWR.n1497 0.365
R9159 VPWR.n1516 VPWR 0.365
R9160 VPWR.n1546 VPWR 0.365
R9161 VPWR.n908 VPWR 0.365
R9162 VPWR VPWR.n3337 0.365
R9163 VPWR.n3219 VPWR 0.365
R9164 VPWR.n2378 VPWR 0.365
R9165 VPWR.n2369 VPWR 0.365
R9166 VPWR.n2359 VPWR 0.365
R9167 VPWR.n2350 VPWR 0.365
R9168 VPWR.n2340 VPWR 0.365
R9169 VPWR.n2998 VPWR 0.365
R9170 VPWR.n2988 VPWR 0.365
R9171 VPWR.n2979 VPWR 0.365
R9172 VPWR.n2969 VPWR 0.365
R9173 VPWR VPWR.n2471 0.365
R9174 VPWR.n2491 VPWR 0.365
R9175 VPWR VPWR.n2611 0.365
R9176 VPWR.n2633 VPWR 0.365
R9177 VPWR.n2624 VPWR 0.365
R9178 VPWR.n3828 VPWR 0.365
R9179 VPWR.n3819 VPWR 0.365
R9180 VPWR VPWR.n46 0.365
R9181 VPWR VPWR.n55 0.365
R9182 VPWR.n3768 VPWR 0.365
R9183 VPWR.n3759 VPWR 0.365
R9184 VPWR VPWR.n3692 0.365
R9185 VPWR VPWR.n1100 0.359
R9186 VPWR VPWR.n1682 0.3575
R9187 VPWR.n1419 VPWR.n1418 0.3545
R9188 VPWR.n973 VPWR.n972 0.35225
R9189 VPWR.n1587 VPWR.n1586 0.3515
R9190 VPWR.n1584 VPWR.n1583 0.3515
R9191 VPWR.n1532 VPWR.n1531 0.3515
R9192 VPWR.n1567 VPWR.n1566 0.3515
R9193 VPWR.n1564 VPWR.n1563 0.3515
R9194 VPWR.n1661 VPWR 0.3515
R9195 VPWR VPWR.n691 0.3515
R9196 VPWR.n1512 VPWR.n1511 0.3485
R9197 VPWR.n1678 VPWR 0.3485
R9198 VPWR.n2903 VPWR.n2902 0.3485
R9199 VPWR VPWR.n967 0.3425
R9200 VPWR.n1577 VPWR.n1576 0.34175
R9201 VPWR VPWR.n1422 0.341
R9202 VPWR VPWR.n1004 0.341
R9203 VPWR.n1449 VPWR.n1448 0.3395
R9204 VPWR.n1557 VPWR.n1556 0.33725
R9205 VPWR.n1551 VPWR.n1550 0.33725
R9206 VPWR.n3449 VPWR.n3444 0.3365
R9207 VPWR.n3456 VPWR.n3455 0.3365
R9208 VPWR.n3454 VPWR.n3453 0.3365
R9209 VPWR.n3453 VPWR.n3452 0.3365
R9210 VPWR.n3452 VPWR.n3451 0.3365
R9211 VPWR.n3464 VPWR.n3459 0.3365
R9212 VPWR.n3471 VPWR.n3470 0.3365
R9213 VPWR.n3469 VPWR.n3468 0.3365
R9214 VPWR.n3468 VPWR.n3467 0.3365
R9215 VPWR.n3467 VPWR.n3466 0.3365
R9216 VPWR.n3479 VPWR.n3474 0.3365
R9217 VPWR.n3486 VPWR.n3485 0.3365
R9218 VPWR.n3484 VPWR.n3483 0.3365
R9219 VPWR.n3483 VPWR.n3482 0.3365
R9220 VPWR.n3482 VPWR.n3481 0.3365
R9221 VPWR.n3494 VPWR.n3489 0.3365
R9222 VPWR.n3501 VPWR.n3500 0.3365
R9223 VPWR.n3499 VPWR.n3498 0.3365
R9224 VPWR.n3498 VPWR.n3497 0.3365
R9225 VPWR.n3497 VPWR.n3496 0.3365
R9226 VPWR.n3509 VPWR.n3504 0.3365
R9227 VPWR.n3516 VPWR.n3515 0.3365
R9228 VPWR.n3514 VPWR.n3513 0.3365
R9229 VPWR.n3513 VPWR.n3512 0.3365
R9230 VPWR.n3512 VPWR.n3511 0.3365
R9231 VPWR.n3524 VPWR.n3519 0.3365
R9232 VPWR.n3531 VPWR.n3530 0.3365
R9233 VPWR.n3529 VPWR.n3528 0.3365
R9234 VPWR.n3528 VPWR.n3527 0.3365
R9235 VPWR.n3527 VPWR.n3526 0.3365
R9236 VPWR.n3539 VPWR.n3534 0.3365
R9237 VPWR.n3546 VPWR.n3545 0.3365
R9238 VPWR.n3544 VPWR.n3543 0.3365
R9239 VPWR.n3543 VPWR.n3542 0.3365
R9240 VPWR.n3542 VPWR.n3541 0.3365
R9241 VPWR.n3554 VPWR.n3549 0.3365
R9242 VPWR.n3561 VPWR.n3560 0.3365
R9243 VPWR.n3559 VPWR.n3558 0.3365
R9244 VPWR.n3558 VPWR.n3557 0.3365
R9245 VPWR.n3557 VPWR.n3556 0.3365
R9246 VPWR.n3569 VPWR.n3564 0.3365
R9247 VPWR.n3576 VPWR.n3575 0.3365
R9248 VPWR.n3574 VPWR.n3573 0.3365
R9249 VPWR.n3573 VPWR.n3572 0.3365
R9250 VPWR.n3572 VPWR.n3571 0.3365
R9251 VPWR.n3584 VPWR.n3579 0.3365
R9252 VPWR.n3591 VPWR.n3590 0.3365
R9253 VPWR.n3589 VPWR.n3588 0.3365
R9254 VPWR.n3588 VPWR.n3587 0.3365
R9255 VPWR.n3587 VPWR.n3586 0.3365
R9256 VPWR.n3599 VPWR.n3594 0.3365
R9257 VPWR.n3606 VPWR.n3605 0.3365
R9258 VPWR.n3604 VPWR.n3603 0.3365
R9259 VPWR.n3603 VPWR.n3602 0.3365
R9260 VPWR.n3602 VPWR.n3601 0.3365
R9261 VPWR.n3614 VPWR.n3609 0.3365
R9262 VPWR.n3621 VPWR.n3620 0.3365
R9263 VPWR.n3619 VPWR.n3618 0.3365
R9264 VPWR.n3618 VPWR.n3617 0.3365
R9265 VPWR.n3617 VPWR.n3616 0.3365
R9266 VPWR.n3629 VPWR.n3624 0.3365
R9267 VPWR.n3636 VPWR.n3635 0.3365
R9268 VPWR.n3634 VPWR.n3633 0.3365
R9269 VPWR.n3633 VPWR.n3632 0.3365
R9270 VPWR.n3632 VPWR.n3631 0.3365
R9271 VPWR.n3644 VPWR.n3639 0.3365
R9272 VPWR.n3651 VPWR.n3650 0.3365
R9273 VPWR.n3649 VPWR.n3648 0.3365
R9274 VPWR.n3648 VPWR.n3647 0.3365
R9275 VPWR.n3647 VPWR.n3646 0.3365
R9276 VPWR.n3659 VPWR.n3654 0.3365
R9277 VPWR.n3666 VPWR.n3665 0.3365
R9278 VPWR.n3664 VPWR.n3663 0.3365
R9279 VPWR.n3663 VPWR.n3662 0.3365
R9280 VPWR.n3662 VPWR.n3661 0.3365
R9281 VPWR.n3674 VPWR.n3669 0.3365
R9282 VPWR.n3681 VPWR.n3680 0.3365
R9283 VPWR.n3679 VPWR.n3678 0.3365
R9284 VPWR.n3678 VPWR.n3677 0.3365
R9285 VPWR.n3677 VPWR.n3676 0.3365
R9286 VPWR.n1075 VPWR.n1074 0.3365
R9287 VPWR.n1479 VPWR.n1478 0.3365
R9288 VPWR.n1491 VPWR.n1490 0.3365
R9289 VPWR.n1492 VPWR.n1491 0.3365
R9290 VPWR.n1493 VPWR.n1492 0.3365
R9291 VPWR.n1495 VPWR.n1494 0.3365
R9292 VPWR.n1496 VPWR.n1495 0.3365
R9293 VPWR.n1497 VPWR.n1496 0.3365
R9294 VPWR.n1505 VPWR.n1504 0.3365
R9295 VPWR.n1504 VPWR.n1503 0.3365
R9296 VPWR.n1503 VPWR.n1502 0.3365
R9297 VPWR.n1501 VPWR.n1500 0.3365
R9298 VPWR.n1500 VPWR.n1499 0.3365
R9299 VPWR.n1499 VPWR.n1498 0.3365
R9300 VPWR VPWR.n1601 0.3365
R9301 VPWR.n1580 VPWR.n1579 0.3365
R9302 VPWR.n1578 VPWR.n1577 0.3365
R9303 VPWR.n1529 VPWR.n1528 0.3365
R9304 VPWR.n1531 VPWR.n1530 0.3365
R9305 VPWR.n1549 VPWR.n1548 0.3365
R9306 VPWR.n1547 VPWR.n1546 0.3365
R9307 VPWR.n1544 VPWR.n1543 0.3365
R9308 VPWR.n1537 VPWR.n1536 0.3365
R9309 VPWR.n1539 VPWR.n1538 0.3365
R9310 VPWR.n1540 VPWR.n1539 0.3365
R9311 VPWR.n1541 VPWR.n1540 0.3365
R9312 VPWR.n979 VPWR.n978 0.3365
R9313 VPWR.n3389 VPWR.n3388 0.3365
R9314 VPWR.n3390 VPWR.n3389 0.3365
R9315 VPWR.n3391 VPWR.n3390 0.3365
R9316 VPWR.n3393 VPWR.n3392 0.3365
R9317 VPWR.n3394 VPWR.n3393 0.3365
R9318 VPWR.n3395 VPWR.n3394 0.3365
R9319 VPWR.n3433 VPWR.n96 0.3365
R9320 VPWR.n3441 VPWR.n3440 0.3365
R9321 VPWR.n3439 VPWR.n3438 0.3365
R9322 VPWR.n3438 VPWR.n3437 0.3365
R9323 VPWR.n3437 VPWR.n3436 0.3365
R9324 VPWR.n1300 VPWR.n1299 0.3365
R9325 VPWR.n1299 VPWR.n1298 0.3365
R9326 VPWR.n3368 VPWR.n3367 0.3365
R9327 VPWR.n3362 VPWR.n3361 0.3365
R9328 VPWR.n3360 VPWR.n3359 0.3365
R9329 VPWR.n779 VPWR.n778 0.3365
R9330 VPWR.n766 VPWR.n765 0.3365
R9331 VPWR.n3284 VPWR.n3283 0.3365
R9332 VPWR.n3281 VPWR.n3280 0.3365
R9333 VPWR.n1724 VPWR.n1723 0.3365
R9334 VPWR.n1727 VPWR.n1726 0.3365
R9335 VPWR.n1775 VPWR.n1774 0.3365
R9336 VPWR.n1772 VPWR.n1771 0.3365
R9337 VPWR.n1807 VPWR 0.3365
R9338 VPWR.n1795 VPWR.n1794 0.3365
R9339 VPWR.n1792 VPWR.n1791 0.3365
R9340 VPWR.n3188 VPWR.n3187 0.3365
R9341 VPWR.n3185 VPWR.n3184 0.3365
R9342 VPWR.n164 VPWR.n163 0.3365
R9343 VPWR.n163 VPWR.n162 0.3365
R9344 VPWR.n162 VPWR.n161 0.3365
R9345 VPWR.n160 VPWR.n159 0.3365
R9346 VPWR.n159 VPWR.n158 0.3365
R9347 VPWR.n158 VPWR.n157 0.3365
R9348 VPWR.n1150 VPWR.n1149 0.3365
R9349 VPWR.n1149 VPWR.n1148 0.3365
R9350 VPWR.n1111 VPWR.n1110 0.3365
R9351 VPWR.n1826 VPWR.n1825 0.3365
R9352 VPWR.n1825 VPWR.n1824 0.3365
R9353 VPWR.n1822 VPWR.n1821 0.3365
R9354 VPWR.n3152 VPWR.n3151 0.3365
R9355 VPWR.n3151 VPWR.n3150 0.3365
R9356 VPWR.n3150 VPWR.n3149 0.3365
R9357 VPWR.n3148 VPWR.n3147 0.3365
R9358 VPWR.n3147 VPWR.n3146 0.3365
R9359 VPWR.n3146 VPWR.n3145 0.3365
R9360 VPWR.n2000 VPWR.n1999 0.3365
R9361 VPWR.n1999 VPWR.n1998 0.3365
R9362 VPWR.n1996 VPWR.n1995 0.3365
R9363 VPWR.n1995 VPWR.n1994 0.3365
R9364 VPWR.n1994 VPWR.n1993 0.3365
R9365 VPWR.n1941 VPWR.n1940 0.3365
R9366 VPWR.n2896 VPWR.n2895 0.3365
R9367 VPWR.n2888 VPWR.n2887 0.3365
R9368 VPWR.n2887 VPWR.n2886 0.3365
R9369 VPWR.n2886 VPWR.n2885 0.3365
R9370 VPWR.n2884 VPWR.n2883 0.3365
R9371 VPWR.n2883 VPWR.n2882 0.3365
R9372 VPWR.n2882 VPWR.n2881 0.3365
R9373 VPWR.n2128 VPWR.n2127 0.3365
R9374 VPWR.n2130 VPWR.n2129 0.3365
R9375 VPWR.n2131 VPWR.n2130 0.3365
R9376 VPWR.n2175 VPWR.n2174 0.3365
R9377 VPWR.n2174 VPWR.n2173 0.3365
R9378 VPWR.n2173 VPWR.n2172 0.3365
R9379 VPWR.n2171 VPWR.n2170 0.3365
R9380 VPWR.n2170 VPWR.n2169 0.3365
R9381 VPWR.n2169 VPWR.n2168 0.3365
R9382 VPWR.n339 VPWR.n338 0.3365
R9383 VPWR.n338 VPWR.n337 0.3365
R9384 VPWR.n337 VPWR.n336 0.3365
R9385 VPWR.n335 VPWR.n334 0.3365
R9386 VPWR.n334 VPWR.n333 0.3365
R9387 VPWR.n333 VPWR.n332 0.3365
R9388 VPWR.n2388 VPWR.n2387 0.3365
R9389 VPWR.n2387 VPWR.n2386 0.3365
R9390 VPWR.n2386 VPWR.n2384 0.3365
R9391 VPWR.n2392 VPWR.n2391 0.3365
R9392 VPWR.n2391 VPWR.n2390 0.3365
R9393 VPWR.n2390 VPWR.n2389 0.3365
R9394 VPWR.n2399 VPWR.n2398 0.3365
R9395 VPWR.n2398 VPWR.n2397 0.3365
R9396 VPWR.n2397 VPWR.n2395 0.3365
R9397 VPWR.n2403 VPWR.n2402 0.3365
R9398 VPWR.n2402 VPWR.n2401 0.3365
R9399 VPWR.n2401 VPWR.n2400 0.3365
R9400 VPWR.n2410 VPWR.n2409 0.3365
R9401 VPWR.n2409 VPWR.n2408 0.3365
R9402 VPWR.n2408 VPWR.n2406 0.3365
R9403 VPWR.n2414 VPWR.n2413 0.3365
R9404 VPWR.n2413 VPWR.n2412 0.3365
R9405 VPWR.n2412 VPWR.n2411 0.3365
R9406 VPWR.n2227 VPWR.n2226 0.3365
R9407 VPWR.n2226 VPWR.n2225 0.3365
R9408 VPWR.n2225 VPWR.n2224 0.3365
R9409 VPWR.n2223 VPWR.n2222 0.3365
R9410 VPWR.n2222 VPWR.n2221 0.3365
R9411 VPWR.n2221 VPWR.n2220 0.3365
R9412 VPWR.n2322 VPWR.n2321 0.3365
R9413 VPWR.n2321 VPWR.n2320 0.3365
R9414 VPWR.n2320 VPWR.n2317 0.3365
R9415 VPWR.n2381 VPWR.n2380 0.3365
R9416 VPWR.n2380 VPWR.n2379 0.3365
R9417 VPWR.n2379 VPWR.n2378 0.3365
R9418 VPWR.n2376 VPWR.n2375 0.3365
R9419 VPWR.n2375 VPWR.n2374 0.3365
R9420 VPWR.n2374 VPWR.n2373 0.3365
R9421 VPWR.n2372 VPWR.n2371 0.3365
R9422 VPWR.n2371 VPWR.n2370 0.3365
R9423 VPWR.n2370 VPWR.n2369 0.3365
R9424 VPWR.n2367 VPWR.n2366 0.3365
R9425 VPWR.n2366 VPWR.n2365 0.3365
R9426 VPWR.n2365 VPWR.n2364 0.3365
R9427 VPWR.n2361 VPWR.n2360 0.3365
R9428 VPWR.n2360 VPWR.n2359 0.3365
R9429 VPWR.n2357 VPWR.n2356 0.3365
R9430 VPWR.n2356 VPWR.n2355 0.3365
R9431 VPWR.n2355 VPWR.n2354 0.3365
R9432 VPWR.n2353 VPWR.n2352 0.3365
R9433 VPWR.n2352 VPWR.n2351 0.3365
R9434 VPWR.n2351 VPWR.n2350 0.3365
R9435 VPWR.n2348 VPWR.n2347 0.3365
R9436 VPWR.n2347 VPWR.n2346 0.3365
R9437 VPWR.n2346 VPWR.n2345 0.3365
R9438 VPWR.n2342 VPWR.n2341 0.3365
R9439 VPWR.n2341 VPWR.n2340 0.3365
R9440 VPWR.n2338 VPWR.n2337 0.3365
R9441 VPWR.n2337 VPWR.n2336 0.3365
R9442 VPWR.n2336 VPWR.n2335 0.3365
R9443 VPWR.n2334 VPWR.n2333 0.3365
R9444 VPWR.n2333 VPWR.n2332 0.3365
R9445 VPWR.n2332 VPWR.n2331 0.3365
R9446 VPWR.n2807 VPWR.n2806 0.3365
R9447 VPWR.n2805 VPWR.n2804 0.3365
R9448 VPWR.n2804 VPWR.n2803 0.3365
R9449 VPWR.n2792 VPWR.n2791 0.3365
R9450 VPWR.n2791 VPWR.n2790 0.3365
R9451 VPWR.n2758 VPWR.n2757 0.3365
R9452 VPWR.n2757 VPWR.n2756 0.3365
R9453 VPWR.n2756 VPWR.n2755 0.3365
R9454 VPWR.n2754 VPWR.n2753 0.3365
R9455 VPWR.n2753 VPWR.n2752 0.3365
R9456 VPWR.n2752 VPWR.n2751 0.3365
R9457 VPWR.n2091 VPWR.n2090 0.3365
R9458 VPWR.n2089 VPWR.n2088 0.3365
R9459 VPWR.n2087 VPWR.n2086 0.3365
R9460 VPWR.n2086 VPWR.n2085 0.3365
R9461 VPWR.n2663 VPWR.n2662 0.3365
R9462 VPWR.n2662 VPWR.n2661 0.3365
R9463 VPWR.n2661 VPWR.n2660 0.3365
R9464 VPWR.n2659 VPWR.n2658 0.3365
R9465 VPWR.n2658 VPWR.n2657 0.3365
R9466 VPWR.n2657 VPWR.n2656 0.3365
R9467 VPWR.n2652 VPWR.n2651 0.3365
R9468 VPWR.n2651 VPWR.n2650 0.3365
R9469 VPWR.n2650 VPWR.n2649 0.3365
R9470 VPWR.n2648 VPWR.n2647 0.3365
R9471 VPWR.n2647 VPWR.n2646 0.3365
R9472 VPWR.n215 VPWR.n214 0.3365
R9473 VPWR.n214 VPWR.n213 0.3365
R9474 VPWR.n213 VPWR.n212 0.3365
R9475 VPWR.n211 VPWR.n210 0.3365
R9476 VPWR.n210 VPWR.n209 0.3365
R9477 VPWR.n209 VPWR.n208 0.3365
R9478 VPWR.n1867 VPWR.n1866 0.3365
R9479 VPWR.n3063 VPWR.n3062 0.3365
R9480 VPWR.n3062 VPWR.n3061 0.3365
R9481 VPWR.n3061 VPWR.n3060 0.3365
R9482 VPWR.n3059 VPWR.n3058 0.3365
R9483 VPWR.n3058 VPWR.n3057 0.3365
R9484 VPWR.n3057 VPWR.n3056 0.3365
R9485 VPWR.n437 VPWR.n436 0.3365
R9486 VPWR.n2996 VPWR.n2995 0.3365
R9487 VPWR.n2995 VPWR.n2994 0.3365
R9488 VPWR.n2994 VPWR.n2993 0.3365
R9489 VPWR.n2992 VPWR.n2991 0.3365
R9490 VPWR.n2989 VPWR.n2988 0.3365
R9491 VPWR.n2986 VPWR.n2985 0.3365
R9492 VPWR.n2985 VPWR.n2984 0.3365
R9493 VPWR.n2984 VPWR.n2983 0.3365
R9494 VPWR.n2982 VPWR.n2981 0.3365
R9495 VPWR.n2981 VPWR.n2980 0.3365
R9496 VPWR.n2980 VPWR.n2979 0.3365
R9497 VPWR.n2977 VPWR.n2976 0.3365
R9498 VPWR.n2976 VPWR.n2975 0.3365
R9499 VPWR.n2975 VPWR.n2974 0.3365
R9500 VPWR.n2973 VPWR.n2972 0.3365
R9501 VPWR.n2970 VPWR.n2969 0.3365
R9502 VPWR.n2967 VPWR.n2966 0.3365
R9503 VPWR.n2966 VPWR.n2965 0.3365
R9504 VPWR.n2965 VPWR.n2964 0.3365
R9505 VPWR.n2963 VPWR.n2962 0.3365
R9506 VPWR.n2962 VPWR.n2961 0.3365
R9507 VPWR.n2961 VPWR.n2960 0.3365
R9508 VPWR.n270 VPWR.n269 0.3365
R9509 VPWR.n271 VPWR.n270 0.3365
R9510 VPWR.n2459 VPWR.n2458 0.3365
R9511 VPWR.n2469 VPWR.n2468 0.3365
R9512 VPWR.n2470 VPWR.n2469 0.3365
R9513 VPWR.n2471 VPWR.n2470 0.3365
R9514 VPWR.n2478 VPWR.n2477 0.3365
R9515 VPWR.n2477 VPWR.n2476 0.3365
R9516 VPWR.n2476 VPWR.n2475 0.3365
R9517 VPWR.n2474 VPWR.n2473 0.3365
R9518 VPWR.n2473 VPWR.n2472 0.3365
R9519 VPWR.n2472 VPWR.n265 0.3365
R9520 VPWR.n2500 VPWR 0.3365
R9521 VPWR.n2498 VPWR.n2497 0.3365
R9522 VPWR.n2497 VPWR.n2496 0.3365
R9523 VPWR.n2496 VPWR.n2495 0.3365
R9524 VPWR.n2494 VPWR.n2493 0.3365
R9525 VPWR.n2493 VPWR.n2492 0.3365
R9526 VPWR.n2492 VPWR.n2491 0.3365
R9527 VPWR.n2489 VPWR.n2488 0.3365
R9528 VPWR.n2488 VPWR.n2487 0.3365
R9529 VPWR.n2487 VPWR.n2486 0.3365
R9530 VPWR.n2485 VPWR.n2484 0.3365
R9531 VPWR.n2484 VPWR.n2483 0.3365
R9532 VPWR.n2483 VPWR.n258 0.3365
R9533 VPWR.n2605 VPWR.n2604 0.3365
R9534 VPWR.n2606 VPWR.n2605 0.3365
R9535 VPWR.n2607 VPWR.n2606 0.3365
R9536 VPWR.n2609 VPWR.n2608 0.3365
R9537 VPWR.n2610 VPWR.n2609 0.3365
R9538 VPWR.n2611 VPWR.n2610 0.3365
R9539 VPWR.n2618 VPWR.n2617 0.3365
R9540 VPWR.n2617 VPWR.n2616 0.3365
R9541 VPWR.n2616 VPWR.n2615 0.3365
R9542 VPWR.n2614 VPWR.n2613 0.3365
R9543 VPWR.n2613 VPWR.n2612 0.3365
R9544 VPWR.n2612 VPWR.n256 0.3365
R9545 VPWR.n2640 VPWR.n2639 0.3365
R9546 VPWR.n2639 VPWR.n2638 0.3365
R9547 VPWR.n2638 VPWR.n2637 0.3365
R9548 VPWR.n2636 VPWR.n2635 0.3365
R9549 VPWR.n2635 VPWR.n2634 0.3365
R9550 VPWR.n2634 VPWR.n2633 0.3365
R9551 VPWR.n2631 VPWR.n2630 0.3365
R9552 VPWR.n2630 VPWR.n2629 0.3365
R9553 VPWR.n2629 VPWR.n2628 0.3365
R9554 VPWR.n2627 VPWR.n2626 0.3365
R9555 VPWR.n2626 VPWR.n2625 0.3365
R9556 VPWR.n2625 VPWR.n2624 0.3365
R9557 VPWR.n3835 VPWR.n3834 0.3365
R9558 VPWR.n3834 VPWR.n3833 0.3365
R9559 VPWR.n3833 VPWR.n3832 0.3365
R9560 VPWR.n3831 VPWR.n3830 0.3365
R9561 VPWR.n3830 VPWR.n3829 0.3365
R9562 VPWR.n3829 VPWR.n3828 0.3365
R9563 VPWR.n3826 VPWR.n3825 0.3365
R9564 VPWR.n3825 VPWR.n3824 0.3365
R9565 VPWR.n3824 VPWR.n3823 0.3365
R9566 VPWR.n3822 VPWR.n3821 0.3365
R9567 VPWR.n3821 VPWR.n3820 0.3365
R9568 VPWR.n3820 VPWR.n3819 0.3365
R9569 VPWR.n40 VPWR.n7 0.3365
R9570 VPWR.n41 VPWR.n40 0.3365
R9571 VPWR.n42 VPWR.n41 0.3365
R9572 VPWR.n44 VPWR.n43 0.3365
R9573 VPWR.n45 VPWR.n44 0.3365
R9574 VPWR.n46 VPWR.n45 0.3365
R9575 VPWR.n49 VPWR.n48 0.3365
R9576 VPWR.n50 VPWR.n49 0.3365
R9577 VPWR.n51 VPWR.n50 0.3365
R9578 VPWR.n53 VPWR.n52 0.3365
R9579 VPWR.n54 VPWR.n53 0.3365
R9580 VPWR.n55 VPWR.n54 0.3365
R9581 VPWR.n3774 VPWR.n3773 0.3365
R9582 VPWR.n3773 VPWR.n3772 0.3365
R9583 VPWR.n3771 VPWR.n3770 0.3365
R9584 VPWR.n3770 VPWR.n3769 0.3365
R9585 VPWR.n3769 VPWR.n3768 0.3365
R9586 VPWR.n3766 VPWR.n3765 0.3365
R9587 VPWR.n3765 VPWR.n3764 0.3365
R9588 VPWR.n3764 VPWR.n3763 0.3365
R9589 VPWR.n3762 VPWR.n3761 0.3365
R9590 VPWR.n3761 VPWR.n3760 0.3365
R9591 VPWR.n3760 VPWR.n3759 0.3365
R9592 VPWR.n3687 VPWR.n60 0.3365
R9593 VPWR.n3688 VPWR.n3687 0.3365
R9594 VPWR.n3690 VPWR.n3689 0.3365
R9595 VPWR.n3691 VPWR.n3690 0.3365
R9596 VPWR.n3692 VPWR.n3691 0.3365
R9597 VPWR.n3695 VPWR.n3694 0.3365
R9598 VPWR.n3696 VPWR.n3695 0.3365
R9599 VPWR.n3697 VPWR.n3696 0.3365
R9600 VPWR.n3699 VPWR.n3698 0.3365
R9601 VPWR.n3705 VPWR.n3684 0.3365
R9602 VPWR.n3713 VPWR.n3712 0.3365
R9603 VPWR.n3711 VPWR.n3710 0.3365
R9604 VPWR.n3710 VPWR.n3709 0.3365
R9605 VPWR.n3709 VPWR.n3708 0.3365
R9606 VPWR.n2450 VPWR.n2449 0.3365
R9607 VPWR.n2449 VPWR.n2448 0.3365
R9608 VPWR.n2448 VPWR.n2447 0.3365
R9609 VPWR.n2436 VPWR.n2435 0.3365
R9610 VPWR.n2435 VPWR.n2434 0.3365
R9611 VPWR.n2434 VPWR.n2433 0.3365
R9612 VPWR.n2431 VPWR.n2430 0.3365
R9613 VPWR.n2430 VPWR.n263 0.3365
R9614 VPWR.n2518 VPWR.n2517 0.3365
R9615 VPWR.n2519 VPWR.n2518 0.3365
R9616 VPWR.n2596 VPWR.n2595 0.3365
R9617 VPWR.n2595 VPWR.n2594 0.3365
R9618 VPWR.n2594 VPWR.n2593 0.3365
R9619 VPWR.n2592 VPWR.n2591 0.3365
R9620 VPWR.n2583 VPWR.n2582 0.3365
R9621 VPWR.n2582 VPWR.n2581 0.3365
R9622 VPWR.n2581 VPWR.n2580 0.3365
R9623 VPWR.n2579 VPWR.n2578 0.3365
R9624 VPWR.n2577 VPWR.n2576 0.3365
R9625 VPWR.n2559 VPWR.n2558 0.3365
R9626 VPWR.n11 VPWR.n2 0.3365
R9627 VPWR.n12 VPWR.n11 0.3365
R9628 VPWR.n13 VPWR.n12 0.3365
R9629 VPWR.n15 VPWR.n14 0.3365
R9630 VPWR.n16 VPWR.n15 0.3365
R9631 VPWR.n29 VPWR.n28 0.3365
R9632 VPWR.n28 VPWR.n27 0.3365
R9633 VPWR.n27 VPWR.n26 0.3365
R9634 VPWR.n25 VPWR.n24 0.3365
R9635 VPWR.n24 VPWR.n23 0.3365
R9636 VPWR.n22 VPWR.n21 0.3365
R9637 VPWR.n65 VPWR.n36 0.3365
R9638 VPWR.n66 VPWR.n65 0.3365
R9639 VPWR.n68 VPWR.n67 0.3365
R9640 VPWR.n69 VPWR.n68 0.3365
R9641 VPWR.n70 VPWR.n69 0.3365
R9642 VPWR.n75 VPWR.n74 0.3365
R9643 VPWR.n76 VPWR.n75 0.3365
R9644 VPWR.n77 VPWR.n76 0.3365
R9645 VPWR.n79 VPWR.n78 0.3365
R9646 VPWR.n80 VPWR.n79 0.3365
R9647 VPWR.n81 VPWR.n80 0.3365
R9648 VPWR.n3719 VPWR.n3718 0.3365
R9649 VPWR.n94 VPWR.n93 0.3365
R9650 VPWR.n92 VPWR.n91 0.3365
R9651 VPWR.n91 VPWR.n90 0.3365
R9652 VPWR.n90 VPWR.n89 0.3365
R9653 VPWR.n1823 VPWR.n1822 0.335
R9654 VPWR.n887 VPWR 0.3335
R9655 VPWR.n798 VPWR.n797 0.3305
R9656 VPWR.n792 VPWR.n791 0.3275
R9657 VPWR VPWR.n1071 0.326
R9658 VPWR.n3376 VPWR.n3375 0.3245
R9659 VPWR.n1073 VPWR.n1072 0.3215
R9660 VPWR.n1481 VPWR.n1480 0.3215
R9661 VPWR.n1625 VPWR.n1624 0.3215
R9662 VPWR VPWR.n1660 0.3215
R9663 VPWR.n871 VPWR.n870 0.3215
R9664 VPWR.n3457 VPWR.n3456 0.3185
R9665 VPWR.n3472 VPWR.n3471 0.3185
R9666 VPWR.n3487 VPWR.n3486 0.3185
R9667 VPWR.n3502 VPWR.n3501 0.3185
R9668 VPWR.n3517 VPWR.n3516 0.3185
R9669 VPWR.n3532 VPWR.n3531 0.3185
R9670 VPWR.n3547 VPWR.n3546 0.3185
R9671 VPWR.n3562 VPWR.n3561 0.3185
R9672 VPWR.n3577 VPWR.n3576 0.3185
R9673 VPWR.n3592 VPWR.n3591 0.3185
R9674 VPWR.n3607 VPWR.n3606 0.3185
R9675 VPWR.n3622 VPWR.n3621 0.3185
R9676 VPWR.n3637 VPWR.n3636 0.3185
R9677 VPWR.n3652 VPWR.n3651 0.3185
R9678 VPWR.n3667 VPWR.n3666 0.3185
R9679 VPWR.n3682 VPWR.n3681 0.3185
R9680 VPWR.n1536 VPWR.n95 0.3185
R9681 VPWR.n3442 VPWR.n3441 0.3185
R9682 VPWR.n3714 VPWR.n3713 0.3185
R9683 VPWR.n3717 VPWR.n94 0.3185
R9684 VPWR.n1818 VPWR.n696 0.317
R9685 VPWR.n581 VPWR.n580 0.317
R9686 VPWR VPWR.n810 0.3155
R9687 VPWR.n401 VPWR.n400 0.314
R9688 VPWR.n1595 VPWR 0.31175
R9689 VPWR VPWR.n1808 0.31175
R9690 VPWR.n2862 VPWR.t325 0.31153
R9691 VPWR.n2864 VPWR.t3852 0.310074
R9692 VPWR.n2362 VPWR.n2361 0.308
R9693 VPWR.n1901 VPWR.n1900 0.308
R9694 VPWR.n2504 VPWR.n2503 0.308
R9695 VPWR VPWR.n1626 0.3065
R9696 VPWR VPWR.n1297 0.3065
R9697 VPWR.n1663 VPWR.n1662 0.3065
R9698 VPWR.n874 VPWR.n873 0.3065
R9699 VPWR.n861 VPWR.n860 0.3065
R9700 VPWR.n3323 VPWR.n3322 0.3065
R9701 VPWR.n3329 VPWR.n3328 0.3065
R9702 VPWR.n1767 VPWR.n699 0.3065
R9703 VPWR VPWR.n674 0.3065
R9704 VPWR VPWR.n645 0.3065
R9705 VPWR.n585 VPWR.n584 0.3065
R9706 VPWR.n579 VPWR.n578 0.3065
R9707 VPWR VPWR.n2831 0.302
R9708 VPWR.n969 VPWR.n968 0.30125
R9709 VPWR.n988 VPWR.n987 0.3005
R9710 VPWR.n1699 VPWR.n1698 0.3005
R9711 VPWR.n3186 VPWR.n3185 0.3005
R9712 VPWR.n417 VPWR 0.299
R9713 VPWR.n1942 VPWR.n1941 0.2975
R9714 VPWR.n1069 VPWR 0.2945
R9715 VPWR.n1648 VPWR.n1647 0.2945
R9716 VPWR.n865 VPWR 0.2945
R9717 VPWR VPWR.n3395 0.29225
R9718 VPWR.n254 VPWR 0.29225
R9719 VPWR.n2432 VPWR 0.29225
R9720 VPWR.n2578 VPWR 0.29225
R9721 VPWR.n23 VPWR 0.29225
R9722 VPWR VPWR.n81 0.29225
R9723 VPWR.n985 VPWR.n984 0.2915
R9724 VPWR.n3366 VPWR.n3365 0.2915
R9725 VPWR.n813 VPWR.n812 0.2915
R9726 VPWR.n3183 VPWR.n3182 0.2915
R9727 VPWR VPWR.n2917 0.2915
R9728 VPWR.n1381 VPWR.n1380 0.29
R9729 VPWR.n3181 VPWR 0.29
R9730 VPWR.n3327 VPWR.n3326 0.2885
R9731 VPWR.n3283 VPWR.n3282 0.2885
R9732 VPWR.n3024 VPWR.n3023 0.2885
R9733 VPWR.n3455 VPWR 0.28775
R9734 VPWR.n3470 VPWR 0.28775
R9735 VPWR.n3485 VPWR 0.28775
R9736 VPWR.n3500 VPWR 0.28775
R9737 VPWR.n3515 VPWR 0.28775
R9738 VPWR.n3530 VPWR 0.28775
R9739 VPWR.n3545 VPWR 0.28775
R9740 VPWR.n3560 VPWR 0.28775
R9741 VPWR.n3575 VPWR 0.28775
R9742 VPWR.n3590 VPWR 0.28775
R9743 VPWR.n3605 VPWR 0.28775
R9744 VPWR.n3620 VPWR 0.28775
R9745 VPWR.n3635 VPWR 0.28775
R9746 VPWR.n3650 VPWR 0.28775
R9747 VPWR.n3665 VPWR 0.28775
R9748 VPWR.n3680 VPWR 0.28775
R9749 VPWR VPWR.n1493 0.28775
R9750 VPWR.n1502 VPWR 0.28775
R9751 VPWR VPWR.n1537 0.28775
R9752 VPWR VPWR.n3391 0.28775
R9753 VPWR.n3440 VPWR 0.28775
R9754 VPWR.n161 VPWR 0.28775
R9755 VPWR.n3149 VPWR 0.28775
R9756 VPWR.n1998 VPWR 0.28775
R9757 VPWR.n1997 VPWR 0.28775
R9758 VPWR.n2885 VPWR 0.28775
R9759 VPWR.n2172 VPWR 0.28775
R9760 VPWR.n336 VPWR 0.28775
R9761 VPWR.n2224 VPWR 0.28775
R9762 VPWR.n2373 VPWR 0.28775
R9763 VPWR.n2364 VPWR 0.28775
R9764 VPWR.n2354 VPWR 0.28775
R9765 VPWR.n2345 VPWR 0.28775
R9766 VPWR.n2335 VPWR 0.28775
R9767 VPWR.n2755 VPWR 0.28775
R9768 VPWR.n2090 VPWR 0.28775
R9769 VPWR.n2088 VPWR 0.28775
R9770 VPWR.n2660 VPWR 0.28775
R9771 VPWR.n2649 VPWR 0.28775
R9772 VPWR.n212 VPWR 0.28775
R9773 VPWR.n3060 VPWR 0.28775
R9774 VPWR.n2993 VPWR 0.28775
R9775 VPWR.n2983 VPWR 0.28775
R9776 VPWR.n2974 VPWR 0.28775
R9777 VPWR.n2964 VPWR 0.28775
R9778 VPWR VPWR.n2467 0.28775
R9779 VPWR.n2475 VPWR 0.28775
R9780 VPWR.n2495 VPWR 0.28775
R9781 VPWR.n2486 VPWR 0.28775
R9782 VPWR VPWR.n2607 0.28775
R9783 VPWR.n2615 VPWR 0.28775
R9784 VPWR.n2637 VPWR 0.28775
R9785 VPWR.n2628 VPWR 0.28775
R9786 VPWR.n3832 VPWR 0.28775
R9787 VPWR.n3823 VPWR 0.28775
R9788 VPWR VPWR.n42 0.28775
R9789 VPWR VPWR.n51 0.28775
R9790 VPWR.n3772 VPWR 0.28775
R9791 VPWR.n3763 VPWR 0.28775
R9792 VPWR VPWR.n3688 0.28775
R9793 VPWR VPWR.n3697 0.28775
R9794 VPWR.n3712 VPWR 0.28775
R9795 VPWR.n2447 VPWR 0.28775
R9796 VPWR.n2433 VPWR 0.28775
R9797 VPWR.n2593 VPWR 0.28775
R9798 VPWR.n2580 VPWR 0.28775
R9799 VPWR VPWR.n13 0.28775
R9800 VPWR.n26 VPWR 0.28775
R9801 VPWR VPWR.n66 0.28775
R9802 VPWR VPWR.n77 0.28775
R9803 VPWR.n93 VPWR 0.28775
R9804 VPWR.n1517 VPWR 0.2825
R9805 VPWR.n1588 VPWR 0.2825
R9806 VPWR.n1585 VPWR 0.2825
R9807 VPWR.n1579 VPWR 0.2825
R9808 VPWR VPWR.n1529 0.2825
R9809 VPWR.n1568 VPWR 0.2825
R9810 VPWR.n1565 VPWR 0.2825
R9811 VPWR.n1558 VPWR 0.2825
R9812 VPWR.n1552 VPWR 0.2825
R9813 VPWR.n1548 VPWR 0.2825
R9814 VPWR.n1009 VPWR.n1008 0.2825
R9815 VPWR.n987 VPWR 0.2825
R9816 VPWR VPWR.n3383 0.2825
R9817 VPWR.n1329 VPWR 0.2825
R9818 VPWR.n1301 VPWR 0.2825
R9819 VPWR.n1654 VPWR 0.2825
R9820 VPWR.n1644 VPWR 0.2825
R9821 VPWR VPWR.n3320 0.2825
R9822 VPWR VPWR.n3330 0.2825
R9823 VPWR.n3361 VPWR 0.2825
R9824 VPWR.n1679 VPWR 0.2825
R9825 VPWR.n776 VPWR 0.2825
R9826 VPWR.n768 VPWR 0.2825
R9827 VPWR.n767 VPWR 0.2825
R9828 VPWR.n765 VPWR 0.2825
R9829 VPWR VPWR.n3235 0.2825
R9830 VPWR.n3246 VPWR 0.2825
R9831 VPWR.n3306 VPWR 0.2825
R9832 VPWR.n3275 VPWR 0.2825
R9833 VPWR VPWR.n1724 0.2825
R9834 VPWR VPWR.n1725 0.2825
R9835 VPWR.n1151 VPWR 0.2825
R9836 VPWR.n679 VPWR 0.2825
R9837 VPWR VPWR.n2128 0.2825
R9838 VPWR.n2806 VPWR 0.2825
R9839 VPWR VPWR.n2931 0.2825
R9840 VPWR VPWR.n2932 0.2825
R9841 VPWR VPWR.n2937 0.2825
R9842 VPWR VPWR.n271 0.2825
R9843 VPWR.n2837 VPWR.n2836 0.2795
R9844 VPWR.n2787 VPWR.n2786 0.2795
R9845 VPWR.n1356 VPWR 0.278
R9846 VPWR.n1014 VPWR.n1013 0.278
R9847 VPWR VPWR.n1131 0.278
R9848 VPWR VPWR.n2030 0.278
R9849 VPWR.n686 VPWR.n685 0.27725
R9850 VPWR.n549 VPWR.n548 0.2765
R9851 VPWR.n879 VPWR 0.275
R9852 VPWR.n1833 VPWR 0.275
R9853 VPWR.n1431 VPWR.n1430 0.27425
R9854 VPWR.n990 VPWR 0.27425
R9855 VPWR.n893 VPWR.n892 0.2735
R9856 VPWR.n3280 VPWR.n3279 0.2735
R9857 VPWR.n1774 VPWR.n1773 0.2735
R9858 VPWR.n1602 VPWR 0.272
R9859 VPWR VPWR.n1075 0.2705
R9860 VPWR VPWR.n669 0.2705
R9861 VPWR.n2913 VPWR.n2912 0.2705
R9862 VPWR.n1012 VPWR 0.2675
R9863 VPWR.n1001 VPWR.n1000 0.2675
R9864 VPWR VPWR.n859 0.2675
R9865 VPWR.n3311 VPWR 0.2675
R9866 VPWR.n3304 VPWR 0.2675
R9867 VPWR VPWR.n673 0.2675
R9868 VPWR.n2843 VPWR.n2842 0.2675
R9869 VPWR.n2946 VPWR 0.2675
R9870 VPWR.n1498 VPWR.n910 0.266
R9871 VPWR.n2642 VPWR.n256 0.266
R9872 VPWR.n2576 VPWR.n2575 0.266
R9873 VPWR.n3379 VPWR 0.2645
R9874 VPWR.n867 VPWR 0.2645
R9875 VPWR.n1737 VPWR.n1736 0.2645
R9876 VPWR.n1790 VPWR.n1789 0.2645
R9877 VPWR VPWR.n1787 0.2645
R9878 VPWR VPWR.n1838 0.2645
R9879 VPWR.n1850 VPWR.n1849 0.2645
R9880 VPWR VPWR.n1627 0.26375
R9881 VPWR.n1739 VPWR 0.263
R9882 VPWR VPWR.n1441 0.2615
R9883 VPWR.n1422 VPWR.n1421 0.2615
R9884 VPWR.n1420 VPWR.n1419 0.2615
R9885 VPWR.n1015 VPWR.n1014 0.2615
R9886 VPWR.n3333 VPWR.n3332 0.2615
R9887 VPWR.n796 VPWR.n795 0.2615
R9888 VPWR.n794 VPWR.n793 0.2615
R9889 VPWR.n3314 VPWR.n3313 0.2615
R9890 VPWR.n2908 VPWR.n2907 0.2615
R9891 VPWR.n2900 VPWR.n2899 0.2615
R9892 VPWR.n2789 VPWR.n2788 0.2615
R9893 VPWR.n2948 VPWR.n2947 0.2615
R9894 VPWR VPWR.n1614 0.2585
R9895 VPWR.n891 VPWR.n890 0.2585
R9896 VPWR VPWR.n2945 0.2585
R9897 VPWR.n1858 VPWR.n1857 0.25775
R9898 VPWR.n1700 VPWR 0.2555
R9899 VPWR.n2990 VPWR.n2989 0.254
R9900 VPWR.n1377 VPWR.n1376 0.2525
R9901 VPWR.n1455 VPWR.n1454 0.2525
R9902 VPWR.n1321 VPWR.n1320 0.2525
R9903 VPWR.n1242 VPWR.n1241 0.2525
R9904 VPWR.n3179 VPWR.n3178 0.2525
R9905 VPWR.n3177 VPWR.n3176 0.2525
R9906 VPWR.n3171 VPWR.n3170 0.2525
R9907 VPWR.n3169 VPWR.n3168 0.2525
R9908 VPWR.n3167 VPWR.n3166 0.2525
R9909 VPWR.n3165 VPWR.n3164 0.2525
R9910 VPWR.n3163 VPWR.n3162 0.2525
R9911 VPWR.n169 VPWR.n168 0.2525
R9912 VPWR.n167 VPWR.n166 0.2525
R9913 VPWR.n1118 VPWR.n1117 0.2525
R9914 VPWR.n672 VPWR.n671 0.2525
R9915 VPWR.n656 VPWR.n655 0.2525
R9916 VPWR.n654 VPWR.n653 0.2525
R9917 VPWR.n652 VPWR.n651 0.2525
R9918 VPWR.n650 VPWR.n649 0.2525
R9919 VPWR.n638 VPWR.n637 0.2525
R9920 VPWR.n636 VPWR.n172 0.2525
R9921 VPWR.n3113 VPWR.n3112 0.2525
R9922 VPWR.n3119 VPWR.n3118 0.2525
R9923 VPWR.n3121 VPWR.n3120 0.2525
R9924 VPWR.n3123 VPWR.n3122 0.2525
R9925 VPWR.n3125 VPWR.n3124 0.2525
R9926 VPWR.n3127 VPWR.n3126 0.2525
R9927 VPWR.n3129 VPWR.n3128 0.2525
R9928 VPWR.n3131 VPWR.n3130 0.2525
R9929 VPWR.n3140 VPWR.n3139 0.2525
R9930 VPWR.n3138 VPWR.n3137 0.2525
R9931 VPWR.n3136 VPWR.n3135 0.2525
R9932 VPWR.n3134 VPWR.n3133 0.2525
R9933 VPWR.n3132 VPWR.n171 0.2525
R9934 VPWR.n3157 VPWR.n3156 0.2525
R9935 VPWR.n3155 VPWR.n3154 0.2525
R9936 VPWR.n1932 VPWR.n1931 0.2525
R9937 VPWR.n1930 VPWR.n1929 0.2525
R9938 VPWR.n1944 VPWR.n1943 0.2525
R9939 VPWR.n352 VPWR.n351 0.2525
R9940 VPWR.n354 VPWR.n353 0.2525
R9941 VPWR.n356 VPWR.n355 0.2525
R9942 VPWR.n358 VPWR.n357 0.2525
R9943 VPWR.n2103 VPWR.n2102 0.2525
R9944 VPWR.n2105 VPWR.n2104 0.2525
R9945 VPWR.n2107 VPWR.n2106 0.2525
R9946 VPWR.n2113 VPWR.n2112 0.2525
R9947 VPWR.n2115 VPWR.n2114 0.2525
R9948 VPWR.n2117 VPWR.n2116 0.2525
R9949 VPWR.n2119 VPWR.n2118 0.2525
R9950 VPWR.n2121 VPWR.n2120 0.2525
R9951 VPWR.n2123 VPWR.n2122 0.2525
R9952 VPWR.n2125 VPWR.n2124 0.2525
R9953 VPWR.n2145 VPWR.n2144 0.2525
R9954 VPWR.n2147 VPWR.n2146 0.2525
R9955 VPWR.n2149 VPWR.n2148 0.2525
R9956 VPWR.n2151 VPWR.n2150 0.2525
R9957 VPWR.n2153 VPWR.n2152 0.2525
R9958 VPWR.n2155 VPWR.n2154 0.2525
R9959 VPWR.n2157 VPWR.n2156 0.2525
R9960 VPWR.n2163 VPWR.n2162 0.2525
R9961 VPWR.n2161 VPWR.n2160 0.2525
R9962 VPWR.n2159 VPWR.n2158 0.2525
R9963 VPWR.n2182 VPWR.n2181 0.2525
R9964 VPWR.n2180 VPWR.n2179 0.2525
R9965 VPWR.n2178 VPWR.n2177 0.2525
R9966 VPWR.n289 VPWR.n288 0.2525
R9967 VPWR.n291 VPWR.n290 0.2525
R9968 VPWR.n293 VPWR.n292 0.2525
R9969 VPWR.n295 VPWR.n294 0.2525
R9970 VPWR.n298 VPWR.n297 0.2525
R9971 VPWR.n300 VPWR.n299 0.2525
R9972 VPWR.n302 VPWR.n301 0.2525
R9973 VPWR.n308 VPWR.n307 0.2525
R9974 VPWR.n310 VPWR.n309 0.2525
R9975 VPWR.n312 VPWR.n311 0.2525
R9976 VPWR.n314 VPWR.n313 0.2525
R9977 VPWR.n316 VPWR.n315 0.2525
R9978 VPWR.n318 VPWR.n317 0.2525
R9979 VPWR.n320 VPWR.n319 0.2525
R9980 VPWR.n327 VPWR.n326 0.2525
R9981 VPWR.n325 VPWR.n324 0.2525
R9982 VPWR.n323 VPWR.n322 0.2525
R9983 VPWR.n321 VPWR.n285 0.2525
R9984 VPWR.n2274 VPWR.n2273 0.2525
R9985 VPWR.n2272 VPWR.n2271 0.2525
R9986 VPWR.n2270 VPWR.n2269 0.2525
R9987 VPWR.n2264 VPWR.n2263 0.2525
R9988 VPWR.n2262 VPWR.n2261 0.2525
R9989 VPWR.n2260 VPWR.n2259 0.2525
R9990 VPWR.n2258 VPWR.n2257 0.2525
R9991 VPWR.n2256 VPWR.n2255 0.2525
R9992 VPWR.n2254 VPWR.n2253 0.2525
R9993 VPWR.n2252 VPWR.n2251 0.2525
R9994 VPWR.n2246 VPWR.n2245 0.2525
R9995 VPWR.n2244 VPWR.n2243 0.2525
R9996 VPWR.n2242 VPWR.n2241 0.2525
R9997 VPWR.n346 VPWR.n345 0.2525
R9998 VPWR.n344 VPWR.n343 0.2525
R9999 VPWR.n342 VPWR.n341 0.2525
R10000 VPWR.n281 VPWR.n280 0.2525
R10001 VPWR.n279 VPWR.n278 0.2525
R10002 VPWR.n277 VPWR.n276 0.2525
R10003 VPWR.n275 VPWR.n274 0.2525
R10004 VPWR.n2314 VPWR.n2313 0.2525
R10005 VPWR.n2312 VPWR.n2311 0.2525
R10006 VPWR.n2310 VPWR.n2309 0.2525
R10007 VPWR.n2304 VPWR.n2303 0.2525
R10008 VPWR.n2302 VPWR.n2301 0.2525
R10009 VPWR.n2300 VPWR.n2299 0.2525
R10010 VPWR.n2298 VPWR.n2297 0.2525
R10011 VPWR.n2296 VPWR.n2295 0.2525
R10012 VPWR.n2294 VPWR.n2293 0.2525
R10013 VPWR.n2292 VPWR.n2291 0.2525
R10014 VPWR.n2286 VPWR.n2285 0.2525
R10015 VPWR.n2284 VPWR.n2283 0.2525
R10016 VPWR.n2282 VPWR.n2281 0.2525
R10017 VPWR.n2280 VPWR.n2279 0.2525
R10018 VPWR.n2187 VPWR.n284 0.2525
R10019 VPWR.n2189 VPWR.n2188 0.2525
R10020 VPWR.n2191 VPWR.n2190 0.2525
R10021 VPWR.n2197 VPWR.n2196 0.2525
R10022 VPWR.n2199 VPWR.n2198 0.2525
R10023 VPWR.n2201 VPWR.n2200 0.2525
R10024 VPWR.n2203 VPWR.n2202 0.2525
R10025 VPWR.n2205 VPWR.n2204 0.2525
R10026 VPWR.n2207 VPWR.n2206 0.2525
R10027 VPWR.n2209 VPWR.n2208 0.2525
R10028 VPWR.n2215 VPWR.n2214 0.2525
R10029 VPWR.n2213 VPWR.n2212 0.2525
R10030 VPWR.n2211 VPWR.n2210 0.2525
R10031 VPWR.n2234 VPWR.n2233 0.2525
R10032 VPWR.n2232 VPWR.n2231 0.2525
R10033 VPWR.n2230 VPWR.n2229 0.2525
R10034 VPWR.n2012 VPWR.n2011 0.2525
R10035 VPWR.n2010 VPWR.n2009 0.2525
R10036 VPWR.n2047 VPWR.n2046 0.2525
R10037 VPWR.n2045 VPWR.n2044 0.2525
R10038 VPWR.n2043 VPWR.n2042 0.2525
R10039 VPWR.n2041 VPWR.n2040 0.2525
R10040 VPWR.n2037 VPWR.n2036 0.2525
R10041 VPWR.n2035 VPWR.n2034 0.2525
R10042 VPWR.n2742 VPWR.n2741 0.2525
R10043 VPWR.n2740 VPWR.n2739 0.2525
R10044 VPWR.n2738 VPWR.n2737 0.2525
R10045 VPWR.n2736 VPWR.n2735 0.2525
R10046 VPWR.n2734 VPWR.n2733 0.2525
R10047 VPWR.n2732 VPWR.n2731 0.2525
R10048 VPWR.n2822 VPWR.n2821 0.2525
R10049 VPWR.n2820 VPWR.n2819 0.2525
R10050 VPWR.n2818 VPWR.n2817 0.2525
R10051 VPWR.n2816 VPWR.n2815 0.2525
R10052 VPWR.n2814 VPWR.n2813 0.2525
R10053 VPWR.n2812 VPWR.n2811 0.2525
R10054 VPWR.n2810 VPWR.n2809 0.2525
R10055 VPWR.n2775 VPWR.n2774 0.2525
R10056 VPWR.n2773 VPWR.n2772 0.2525
R10057 VPWR.n2771 VPWR.n2770 0.2525
R10058 VPWR.n2769 VPWR.n2768 0.2525
R10059 VPWR.n2767 VPWR.n2766 0.2525
R10060 VPWR.n2765 VPWR.n2764 0.2525
R10061 VPWR.n2761 VPWR.n2760 0.2525
R10062 VPWR.n595 VPWR.n594 0.2525
R10063 VPWR.n3036 VPWR.n3035 0.2525
R10064 VPWR.n3038 VPWR.n3037 0.2525
R10065 VPWR.n3040 VPWR.n3039 0.2525
R10066 VPWR.n3042 VPWR.n3041 0.2525
R10067 VPWR.n3051 VPWR.n3050 0.2525
R10068 VPWR.n3049 VPWR.n3048 0.2525
R10069 VPWR.n3047 VPWR.n3046 0.2525
R10070 VPWR.n3045 VPWR.n3044 0.2525
R10071 VPWR.n3043 VPWR.n173 0.2525
R10072 VPWR.n3105 VPWR.n3104 0.2525
R10073 VPWR.n3103 VPWR.n3102 0.2525
R10074 VPWR.n3097 VPWR.n3096 0.2525
R10075 VPWR.n3095 VPWR.n3094 0.2525
R10076 VPWR.n3093 VPWR.n3092 0.2525
R10077 VPWR.n3091 VPWR.n3090 0.2525
R10078 VPWR.n3089 VPWR.n3088 0.2525
R10079 VPWR.n3087 VPWR.n3086 0.2525
R10080 VPWR.n3085 VPWR.n3084 0.2525
R10081 VPWR.n3079 VPWR.n3078 0.2525
R10082 VPWR.n3077 VPWR.n3076 0.2525
R10083 VPWR.n3075 VPWR.n3074 0.2525
R10084 VPWR.n3073 VPWR.n3072 0.2525
R10085 VPWR.n3071 VPWR.n3070 0.2525
R10086 VPWR.n3068 VPWR.n3067 0.2525
R10087 VPWR.n3066 VPWR.n3065 0.2525
R10088 VPWR.n1903 VPWR.n1902 0.2525
R10089 VPWR.n435 VPWR.n434 0.2525
R10090 VPWR.n427 VPWR.n426 0.2525
R10091 VPWR.n3011 VPWR.n3010 0.2525
R10092 VPWR.n3009 VPWR.n3008 0.2525
R10093 VPWR.n3007 VPWR.n3006 0.2525
R10094 VPWR.n3003 VPWR.n3002 0.2525
R10095 VPWR.n3001 VPWR.n3000 0.2525
R10096 VPWR VPWR.n1835 0.2495
R10097 VPWR.n2857 VPWR.n2856 0.2495
R10098 VPWR VPWR.n2915 0.24875
R10099 VPWR.n3303 VPWR 0.248
R10100 VPWR.n2393 VPWR.n2384 0.2465
R10101 VPWR.n2404 VPWR.n2395 0.2465
R10102 VPWR.n2415 VPWR.n2406 0.2465
R10103 VPWR.n2382 VPWR.n2317 0.2465
R10104 VPWR.n2457 VPWR.n272 0.2465
R10105 VPWR.n666 VPWR 0.245
R10106 VPWR.n2920 VPWR.n184 0.245
R10107 VPWR.n1237 VPWR.n1236 0.2435
R10108 VPWR VPWR.n3198 0.2435
R10109 VPWR.n2796 VPWR 0.242
R10110 VPWR.n3364 VPWR 0.24125
R10111 VPWR VPWR.n2845 0.24125
R10112 VPWR.n1690 VPWR 0.2405
R10113 VPWR.n1756 VPWR.n1755 0.2405
R10114 VPWR.n1115 VPWR 0.2405
R10115 VPWR.n2645 VPWR.n254 0.239
R10116 VPWR.n2455 VPWR 0.237875
R10117 VPWR.n2502 VPWR 0.237875
R10118 VPWR.n2600 VPWR 0.237875
R10119 VPWR.n255 VPWR 0.237875
R10120 VPWR.n3838 VPWR 0.237875
R10121 VPWR.n3815 VPWR 0.237875
R10122 VPWR.n3777 VPWR 0.237875
R10123 VPWR.n3716 VPWR 0.237875
R10124 VPWR.n3754 VPWR 0.237875
R10125 VPWR.n1631 VPWR.n1630 0.2375
R10126 VPWR.n903 VPWR.n902 0.2375
R10127 VPWR VPWR.n3209 0.2375
R10128 VPWR.n3757 VPWR.n3756 0.236
R10129 VPWR.n1327 VPWR 0.23525
R10130 VPWR VPWR.n1735 0.2345
R10131 VPWR.n1758 VPWR 0.2345
R10132 VPWR.n3221 VPWR 0.2345
R10133 VPWR.n1863 VPWR.n1862 0.2345
R10134 VPWR.n1701 VPWR 0.233
R10135 VPWR VPWR.n1105 0.233
R10136 VPWR.n1743 VPWR.n1742 0.2315
R10137 VPWR.n2902 VPWR.n2901 0.2315
R10138 VPWR.n2184 VPWR.n348 0.2315
R10139 VPWR.n2240 VPWR.n2239 0.2315
R10140 VPWR.n2236 VPWR.n2186 0.2315
R10141 VPWR.n3030 VPWR.n3029 0.2315
R10142 VPWR.n399 VPWR 0.2315
R10143 VPWR.n583 VPWR.n582 0.23
R10144 VPWR.n1478 VPWR 0.2285
R10145 VPWR.n3296 VPWR.n3295 0.2285
R10146 VPWR.n3278 VPWR.n3277 0.2285
R10147 VPWR.n662 VPWR.n661 0.2285
R10148 VPWR VPWR.n2891 0.2285
R10149 VPWR.n884 VPWR.n883 0.2255
R10150 VPWR.n586 VPWR 0.2255
R10151 VPWR.n1828 VPWR 0.22475
R10152 VPWR VPWR.n1596 0.22325
R10153 VPWR VPWR.n1559 0.22325
R10154 VPWR VPWR.n1554 0.22325
R10155 VPWR VPWR.n1292 0.22325
R10156 VPWR.n426 VPWR 0.22325
R10157 VPWR.n1477 VPWR 0.2225
R10158 VPWR.n1594 VPWR 0.2225
R10159 VPWR VPWR.n1588 0.2225
R10160 VPWR VPWR.n1580 0.2225
R10161 VPWR.n1528 VPWR 0.2225
R10162 VPWR.n1457 VPWR 0.2225
R10163 VPWR.n1445 VPWR 0.2225
R10164 VPWR VPWR.n1436 0.2225
R10165 VPWR VPWR.n1416 0.2225
R10166 VPWR.n3383 VPWR 0.2225
R10167 VPWR VPWR.n1301 0.2225
R10168 VPWR VPWR.n1243 0.2225
R10169 VPWR VPWR.n1683 0.2225
R10170 VPWR VPWR.n3230 0.2225
R10171 VPWR.n1732 VPWR 0.2225
R10172 VPWR VPWR.n1795 0.2225
R10173 VPWR VPWR.n3203 0.2225
R10174 VPWR VPWR.n3188 0.2225
R10175 VPWR VPWR.n3172 0.2225
R10176 VPWR VPWR.n1151 0.2225
R10177 VPWR.n3117 VPWR 0.2225
R10178 VPWR VPWR.n3141 0.2225
R10179 VPWR VPWR.n2000 0.2225
R10180 VPWR VPWR.n1970 0.2225
R10181 VPWR VPWR.n1956 0.2225
R10182 VPWR VPWR.n1947 0.2225
R10183 VPWR.n2111 VPWR 0.2225
R10184 VPWR.n2137 VPWR 0.2225
R10185 VPWR.n2143 VPWR 0.2225
R10186 VPWR VPWR.n2164 0.2225
R10187 VPWR.n306 VPWR 0.2225
R10188 VPWR VPWR.n328 0.2225
R10189 VPWR VPWR.n2265 0.2225
R10190 VPWR VPWR.n2247 0.2225
R10191 VPWR VPWR.n2305 0.2225
R10192 VPWR VPWR.n2287 0.2225
R10193 VPWR.n2195 VPWR 0.2225
R10194 VPWR VPWR.n2216 0.2225
R10195 VPWR VPWR.n2743 0.2225
R10196 VPWR VPWR.n2823 0.2225
R10197 VPWR VPWR.n2782 0.2225
R10198 VPWR VPWR.n2780 0.2225
R10199 VPWR VPWR.n2776 0.2225
R10200 VPWR VPWR.n2683 0.2225
R10201 VPWR VPWR.n1867 0.2225
R10202 VPWR.n3028 VPWR 0.2225
R10203 VPWR VPWR.n3052 0.2225
R10204 VPWR VPWR.n3098 0.2225
R10205 VPWR VPWR.n3080 0.2225
R10206 VPWR VPWR.n440 0.2225
R10207 VPWR.n2931 VPWR 0.2225
R10208 VPWR.n2517 VPWR 0.2225
R10209 VPWR VPWR.n2559 0.2225
R10210 VPWR VPWR.n3798 0.2225
R10211 VPWR VPWR.n970 0.22025
R10212 VPWR VPWR.n683 0.22025
R10213 VPWR.n1017 VPWR.n1016 0.2195
R10214 VPWR.n1646 VPWR.n1645 0.2195
R10215 VPWR.n1753 VPWR.n1752 0.2195
R10216 VPWR.n690 VPWR.n689 0.2195
R10217 VPWR.n419 VPWR 0.2195
R10218 VPWR.n2999 VPWR.n2998 0.2195
R10219 VPWR.n3775 VPWR.n3774 0.2195
R10220 VPWR.n3778 VPWR.n36 0.2195
R10221 VPWR VPWR.n1488 0.218
R10222 VPWR VPWR.n2602 0.218
R10223 VPWR.n3242 VPWR.n3241 0.21725
R10224 VPWR VPWR.n3300 0.2165
R10225 VPWR.n2897 VPWR.n2896 0.2165
R10226 VPWR.n1820 VPWR.n1819 0.215
R10227 VPWR.n3249 VPWR 0.21425
R10228 VPWR.n1379 VPWR 0.2135
R10229 VPWR.n873 VPWR.n872 0.2135
R10230 VPWR.n552 VPWR 0.2135
R10231 VPWR.n563 VPWR.n562 0.21275
R10232 VPWR VPWR.n1366 0.212
R10233 VPWR.n1617 VPWR.n1616 0.212
R10234 VPWR.n1665 VPWR.n1664 0.2105
R10235 VPWR.n573 VPWR 0.2105
R10236 VPWR VPWR.n1073 0.209
R10237 VPWR.n1480 VPWR 0.209
R10238 VPWR VPWR.n811 0.209
R10239 VPWR.n3287 VPWR 0.209
R10240 VPWR.n1731 VPWR.n1730 0.209
R10241 VPWR.n567 VPWR.n566 0.20825
R10242 VPWR VPWR.n1634 0.2075
R10243 VPWR.n1688 VPWR.n1687 0.2075
R10244 VPWR.n1113 VPWR.n1112 0.2075
R10245 VPWR.n1230 VPWR 0.206
R10246 VPWR.n3276 VPWR 0.206
R10247 VPWR VPWR.n1515 0.2045
R10248 VPWR.n778 VPWR.n777 0.2045
R10249 VPWR.n547 VPWR.n546 0.2045
R10250 VPWR.n1116 VPWR 0.20375
R10251 VPWR.n1835 VPWR 0.20375
R10252 VPWR.n2039 VPWR 0.20375
R10253 VPWR.n3005 VPWR 0.20375
R10254 VPWR.n3211 VPWR.n3210 0.2015
R10255 VPWR.n1907 VPWR 0.2015
R10256 VPWR.n2927 VPWR.n2926 0.2015
R10257 VPWR.n2972 VPWR.n2971 0.2015
R10258 VPWR.n1007 VPWR 0.19925
R10259 VPWR VPWR.n3447 0.1985
R10260 VPWR VPWR.n3462 0.1985
R10261 VPWR VPWR.n3477 0.1985
R10262 VPWR VPWR.n3492 0.1985
R10263 VPWR VPWR.n3507 0.1985
R10264 VPWR VPWR.n3522 0.1985
R10265 VPWR VPWR.n3537 0.1985
R10266 VPWR VPWR.n3552 0.1985
R10267 VPWR VPWR.n3567 0.1985
R10268 VPWR VPWR.n3582 0.1985
R10269 VPWR VPWR.n3597 0.1985
R10270 VPWR VPWR.n3612 0.1985
R10271 VPWR VPWR.n3627 0.1985
R10272 VPWR VPWR.n3642 0.1985
R10273 VPWR VPWR.n3657 0.1985
R10274 VPWR VPWR.n3672 0.1985
R10275 VPWR.n1475 VPWR 0.1985
R10276 VPWR VPWR.n1520 0.1985
R10277 VPWR.n1519 VPWR 0.1985
R10278 VPWR VPWR.n1518 0.1985
R10279 VPWR.n1598 VPWR 0.1985
R10280 VPWR VPWR.n1594 0.1985
R10281 VPWR.n1574 VPWR 0.1985
R10282 VPWR.n1357 VPWR 0.1985
R10283 VPWR VPWR.n1364 0.1985
R10284 VPWR VPWR.n1610 0.1985
R10285 VPWR.n991 VPWR 0.1985
R10286 VPWR.n989 VPWR 0.1985
R10287 VPWR.n975 VPWR.n974 0.1985
R10288 VPWR.n1271 VPWR 0.1985
R10289 VPWR.n1333 VPWR 0.1985
R10290 VPWR.n1323 VPWR 0.1985
R10291 VPWR.n1289 VPWR 0.1985
R10292 VPWR.n880 VPWR 0.1985
R10293 VPWR VPWR.n3334 0.1985
R10294 VPWR.n3344 VPWR.n3343 0.1985
R10295 VPWR VPWR.n1261 0.1985
R10296 VPWR.n1248 VPWR 0.1985
R10297 VPWR VPWR.n1681 0.1985
R10298 VPWR.n808 VPWR 0.1985
R10299 VPWR.n3315 VPWR 0.1985
R10300 VPWR VPWR.n3307 0.1985
R10301 VPWR VPWR.n1200 0.1985
R10302 VPWR VPWR.n1197 0.1985
R10303 VPWR VPWR.n1194 0.1985
R10304 VPWR.n1185 VPWR 0.1985
R10305 VPWR.n1713 VPWR 0.1985
R10306 VPWR VPWR.n1085 0.1985
R10307 VPWR.n1084 VPWR 0.1985
R10308 VPWR.n1148 VPWR 0.1985
R10309 VPWR.n1103 VPWR.n1102 0.1985
R10310 VPWR.n687 VPWR 0.1985
R10311 VPWR.n674 VPWR 0.1985
R10312 VPWR.n667 VPWR 0.1985
R10313 VPWR.n640 VPWR 0.1985
R10314 VPWR VPWR.n3110 0.1985
R10315 VPWR.n1928 VPWR 0.1985
R10316 VPWR.n1955 VPWR 0.1985
R10317 VPWR VPWR.n2840 0.1985
R10318 VPWR VPWR.n2844 0.1985
R10319 VPWR VPWR.n2131 0.1985
R10320 VPWR VPWR.n2138 0.1985
R10321 VPWR.n2008 VPWR 0.1985
R10322 VPWR.n2049 VPWR 0.1985
R10323 VPWR.n2082 VPWR 0.1985
R10324 VPWR.n2695 VPWR 0.1985
R10325 VPWR VPWR.n1879 0.1985
R10326 VPWR.n597 VPWR 0.1985
R10327 VPWR.n1920 VPWR 0.1985
R10328 VPWR.n1909 VPWR 0.1985
R10329 VPWR.n444 VPWR 0.1985
R10330 VPWR.n439 VPWR 0.1985
R10331 VPWR.n2939 VPWR 0.1985
R10332 VPWR VPWR.n2465 0.1985
R10333 VPWR VPWR.n3413 0.197
R10334 VPWR VPWR.n3432 0.197
R10335 VPWR VPWR.n869 0.197
R10336 VPWR.n1142 VPWR 0.197
R10337 VPWR.n1973 VPWR 0.197
R10338 VPWR VPWR.n2711 0.197
R10339 VPWR.n2093 VPWR 0.197
R10340 VPWR.n2686 VPWR 0.197
R10341 VPWR.n2665 VPWR 0.197
R10342 VPWR.n237 VPWR 0.197
R10343 VPWR.n217 VPWR 0.197
R10344 VPWR.n1923 VPWR 0.197
R10345 VPWR VPWR.n3704 0.197
R10346 VPWR.n2452 VPWR 0.197
R10347 VPWR.n2438 VPWR 0.197
R10348 VPWR VPWR.n2514 0.197
R10349 VPWR.n2598 VPWR 0.197
R10350 VPWR.n2585 VPWR 0.197
R10351 VPWR.n2562 VPWR 0.197
R10352 VPWR VPWR.n0 0.197
R10353 VPWR VPWR.n20 0.197
R10354 VPWR.n3801 VPWR 0.197
R10355 VPWR.n3781 VPWR 0.197
R10356 VPWR.n3740 VPWR 0.197
R10357 VPWR.n3721 VPWR 0.197
R10358 VPWR.n1659 VPWR 0.1955
R10359 VPWR.n3224 VPWR.n131 0.1955
R10360 VPWR VPWR.n1806 0.1955
R10361 VPWR.n1831 VPWR.n1830 0.1955
R10362 VPWR.n1639 VPWR 0.194
R10363 VPWR VPWR.n1257 0.194
R10364 VPWR VPWR.n465 0.194
R10365 VPWR.n1078 VPWR 0.1925
R10366 VPWR VPWR.n3347 0.1925
R10367 VPWR.n1110 VPWR.n1109 0.1925
R10368 VPWR.n1013 VPWR.n1012 0.191
R10369 VPWR.n1642 VPWR.n909 0.191
R10370 VPWR.n1416 VPWR.n1415 0.1895
R10371 VPWR.n775 VPWR.n774 0.1895
R10372 VPWR.n3209 VPWR.n3208 0.1895
R10373 VPWR.n3202 VPWR 0.1895
R10374 VPWR.n2343 VPWR.n2342 0.1895
R10375 VPWR.n2828 VPWR.n2827 0.1895
R10376 VPWR VPWR.n3233 0.188
R10377 VPWR.n1183 VPWR.n1182 0.188
R10378 VPWR.n1855 VPWR.n1854 0.18725
R10379 VPWR.n1352 VPWR 0.1865
R10380 VPWR.n863 VPWR 0.1865
R10381 VPWR.n815 VPWR.n814 0.1865
R10382 VPWR.n3250 VPWR 0.1865
R10383 VPWR.n1729 VPWR.n1728 0.1865
R10384 VPWR.n3213 VPWR.n3212 0.1865
R10385 VPWR VPWR.n1086 0.1865
R10386 VPWR.n1805 VPWR 0.18575
R10387 VPWR.n592 VPWR 0.18575
R10388 VPWR VPWR.n432 0.18575
R10389 VPWR.n1003 VPWR.n1002 0.1835
R10390 VPWR.n886 VPWR.n885 0.1835
R10391 VPWR.n799 VPWR 0.1835
R10392 VPWR.n763 VPWR.n762 0.1835
R10393 VPWR.n3232 VPWR.n3231 0.1835
R10394 VPWR.n1740 VPWR.n1739 0.1835
R10395 VPWR.n1801 VPWR 0.1835
R10396 VPWR.n1841 VPWR.n1840 0.1835
R10397 VPWR.n1832 VPWR.n1831 0.1835
R10398 VPWR.n1236 VPWR.n1235 0.18275
R10399 VPWR VPWR.n1435 0.18125
R10400 VPWR.n803 VPWR 0.18125
R10401 VPWR VPWR.n1469 0.1805
R10402 VPWR.n3252 VPWR.n3251 0.1805
R10403 VPWR VPWR.n3303 0.1805
R10404 VPWR.n3197 VPWR.n3196 0.1805
R10405 VPWR VPWR.n2802 0.1805
R10406 VPWR.n2801 VPWR.n2800 0.1805
R10407 VPWR VPWR.n3014 0.1805
R10408 VPWR VPWR.n3226 0.1775
R10409 VPWR.n1949 VPWR.n1948 0.1775
R10410 VPWR.n2894 VPWR 0.1775
R10411 VPWR.n1866 VPWR.n1865 0.1775
R10412 VPWR.n550 VPWR 0.1775
R10413 VPWR VPWR.n1474 0.176
R10414 VPWR.n1573 VPWR 0.176
R10415 VPWR.n1562 VPWR 0.176
R10416 VPWR.n1624 VPWR.n1623 0.176
R10417 VPWR.n1613 VPWR.n1612 0.176
R10418 VPWR.n966 VPWR 0.176
R10419 VPWR.n1325 VPWR 0.176
R10420 VPWR.n3206 VPWR 0.176
R10421 VPWR.n1122 VPWR 0.176
R10422 VPWR.n1953 VPWR 0.176
R10423 VPWR.n2080 VPWR 0.176
R10424 VPWR.n1913 VPWR 0.176
R10425 VPWR.n454 VPWR 0.176
R10426 VPWR.n416 VPWR 0.176
R10427 VPWR.n1748 VPWR.n1747 0.1745
R10428 VPWR.n1750 VPWR.n1749 0.1745
R10429 VPWR VPWR.n564 0.1745
R10430 VPWR.n3025 VPWR 0.1745
R10431 VPWR VPWR.n415 0.173
R10432 VPWR.n1621 VPWR.n1620 0.1715
R10433 VPWR.n902 VPWR 0.1715
R10434 VPWR VPWR.n1753 0.1715
R10435 VPWR VPWR.n2911 0.1715
R10436 VPWR.n1510 VPWR 0.17075
R10437 VPWR.n1734 VPWR 0.17075
R10438 VPWR.n1430 VPWR 0.17
R10439 VPWR.n3316 VPWR.n3315 0.17
R10440 VPWR.n1601 VPWR 0.16925
R10441 VPWR.n3299 VPWR 0.16925
R10442 VPWR.n2910 VPWR 0.16925
R10443 VPWR.n3380 VPWR.n3379 0.1685
R10444 VPWR.n3381 VPWR.n3380 0.1685
R10445 VPWR.n3399 VPWR.n3398 0.1685
R10446 VPWR.n3402 VPWR.n3401 0.1685
R10447 VPWR.n3403 VPWR.n3402 0.1685
R10448 VPWR.n3404 VPWR.n3403 0.1685
R10449 VPWR.n3405 VPWR.n3404 0.1685
R10450 VPWR.n3406 VPWR.n3405 0.1685
R10451 VPWR.n3408 VPWR.n3407 0.1685
R10452 VPWR.n3409 VPWR.n3408 0.1685
R10453 VPWR.n3410 VPWR.n3409 0.1685
R10454 VPWR.n3411 VPWR.n3410 0.1685
R10455 VPWR.n3412 VPWR.n3411 0.1685
R10456 VPWR.n3413 VPWR.n3412 0.1685
R10457 VPWR.n3418 VPWR.n3417 0.1685
R10458 VPWR.n3419 VPWR.n3418 0.1685
R10459 VPWR.n3420 VPWR.n3419 0.1685
R10460 VPWR.n3421 VPWR.n3420 0.1685
R10461 VPWR.n3422 VPWR.n3421 0.1685
R10462 VPWR.n3423 VPWR.n3422 0.1685
R10463 VPWR.n3424 VPWR.n3423 0.1685
R10464 VPWR.n3426 VPWR.n3425 0.1685
R10465 VPWR.n3427 VPWR.n3426 0.1685
R10466 VPWR.n3428 VPWR.n3427 0.1685
R10467 VPWR.n3429 VPWR.n3428 0.1685
R10468 VPWR.n3430 VPWR.n3429 0.1685
R10469 VPWR.n3431 VPWR.n3430 0.1685
R10470 VPWR.n3432 VPWR.n3431 0.1685
R10471 VPWR.n1317 VPWR 0.1685
R10472 VPWR.n3346 VPWR.n3345 0.1685
R10473 VPWR.n1232 VPWR.n1231 0.1685
R10474 VPWR VPWR.n1715 0.1685
R10475 VPWR.n3198 VPWR.n3197 0.1685
R10476 VPWR.n1145 VPWR.n1144 0.1685
R10477 VPWR.n1143 VPWR.n1142 0.1685
R10478 VPWR.n2799 VPWR.n2798 0.1685
R10479 VPWR.n2062 VPWR.n2061 0.1685
R10480 VPWR.n2061 VPWR.n2060 0.1685
R10481 VPWR.n2059 VPWR.n2058 0.1685
R10482 VPWR.n2058 VPWR.n2057 0.1685
R10483 VPWR.n2056 VPWR.n2055 0.1685
R10484 VPWR.n2096 VPWR.n2095 0.1685
R10485 VPWR.n2095 VPWR.n2094 0.1685
R10486 VPWR.n2094 VPWR.n2093 0.1685
R10487 VPWR.n2690 VPWR.n2689 0.1685
R10488 VPWR.n2689 VPWR.n2688 0.1685
R10489 VPWR.n2687 VPWR.n2686 0.1685
R10490 VPWR.n2681 VPWR.n2680 0.1685
R10491 VPWR.n2680 VPWR.n2679 0.1685
R10492 VPWR.n2679 VPWR.n2678 0.1685
R10493 VPWR.n2678 VPWR.n2677 0.1685
R10494 VPWR.n2677 VPWR.n2676 0.1685
R10495 VPWR.n2676 VPWR.n2675 0.1685
R10496 VPWR.n2675 VPWR.n2674 0.1685
R10497 VPWR.n2673 VPWR.n2672 0.1685
R10498 VPWR.n2672 VPWR.n2671 0.1685
R10499 VPWR.n2671 VPWR.n2670 0.1685
R10500 VPWR.n2668 VPWR.n2667 0.1685
R10501 VPWR.n2667 VPWR.n2666 0.1685
R10502 VPWR.n251 VPWR.n250 0.1685
R10503 VPWR.n250 VPWR.n249 0.1685
R10504 VPWR.n249 VPWR.n248 0.1685
R10505 VPWR.n248 VPWR.n247 0.1685
R10506 VPWR.n247 VPWR.n246 0.1685
R10507 VPWR.n246 VPWR.n245 0.1685
R10508 VPWR.n245 VPWR.n244 0.1685
R10509 VPWR.n243 VPWR.n242 0.1685
R10510 VPWR.n242 VPWR.n241 0.1685
R10511 VPWR.n241 VPWR.n240 0.1685
R10512 VPWR.n240 VPWR.n239 0.1685
R10513 VPWR.n239 VPWR.n238 0.1685
R10514 VPWR.n238 VPWR.n237 0.1685
R10515 VPWR.n233 VPWR.n232 0.1685
R10516 VPWR.n232 VPWR.n231 0.1685
R10517 VPWR.n231 VPWR.n230 0.1685
R10518 VPWR.n230 VPWR.n229 0.1685
R10519 VPWR.n229 VPWR.n228 0.1685
R10520 VPWR.n228 VPWR.n227 0.1685
R10521 VPWR.n227 VPWR.n226 0.1685
R10522 VPWR.n225 VPWR.n224 0.1685
R10523 VPWR.n224 VPWR.n223 0.1685
R10524 VPWR.n223 VPWR.n222 0.1685
R10525 VPWR.n222 VPWR.n221 0.1685
R10526 VPWR.n221 VPWR.n220 0.1685
R10527 VPWR.n218 VPWR.n217 0.1685
R10528 VPWR.n366 VPWR.n365 0.1685
R10529 VPWR.n363 VPWR.n360 0.1685
R10530 VPWR.n415 VPWR.n414 0.1685
R10531 VPWR.n413 VPWR.n412 0.1685
R10532 VPWR.n411 VPWR.n410 0.1685
R10533 VPWR.n409 VPWR.n408 0.1685
R10534 VPWR.n2462 VPWR.n2461 0.1685
R10535 VPWR.n2463 VPWR.n2462 0.1685
R10536 VPWR.n2464 VPWR.n2463 0.1685
R10537 VPWR.n2465 VPWR.n2464 0.1685
R10538 VPWR.n3703 VPWR.n3702 0.1685
R10539 VPWR.n2423 VPWR.n2422 0.1685
R10540 VPWR.n2422 VPWR.n2421 0.1685
R10541 VPWR.n2421 VPWR.n2420 0.1685
R10542 VPWR.n2420 VPWR.n2419 0.1685
R10543 VPWR.n2418 VPWR.n2417 0.1685
R10544 VPWR.n2453 VPWR.n2452 0.1685
R10545 VPWR.n2443 VPWR.n2442 0.1685
R10546 VPWR.n2442 VPWR.n2441 0.1685
R10547 VPWR.n2441 VPWR.n2440 0.1685
R10548 VPWR.n2440 VPWR.n2439 0.1685
R10549 VPWR.n2439 VPWR.n2438 0.1685
R10550 VPWR.n2507 VPWR.n2506 0.1685
R10551 VPWR.n2508 VPWR.n2507 0.1685
R10552 VPWR.n2509 VPWR.n2508 0.1685
R10553 VPWR.n2510 VPWR.n2509 0.1685
R10554 VPWR.n2511 VPWR.n2510 0.1685
R10555 VPWR.n2512 VPWR.n2511 0.1685
R10556 VPWR.n2513 VPWR.n2512 0.1685
R10557 VPWR.n2533 VPWR.n2532 0.1685
R10558 VPWR.n2532 VPWR.n2531 0.1685
R10559 VPWR.n2531 VPWR.n2530 0.1685
R10560 VPWR.n2530 VPWR.n2529 0.1685
R10561 VPWR.n2529 VPWR.n2528 0.1685
R10562 VPWR.n2528 VPWR.n2527 0.1685
R10563 VPWR.n2527 VPWR.n2526 0.1685
R10564 VPWR.n2525 VPWR.n2524 0.1685
R10565 VPWR.n2524 VPWR.n2523 0.1685
R10566 VPWR.n2522 VPWR.n2521 0.1685
R10567 VPWR.n2521 VPWR.n2520 0.1685
R10568 VPWR.n2520 VPWR.n260 0.1685
R10569 VPWR.n2588 VPWR.n2587 0.1685
R10570 VPWR.n2587 VPWR.n2586 0.1685
R10571 VPWR.n2586 VPWR.n2585 0.1685
R10572 VPWR.n2572 VPWR.n2571 0.1685
R10573 VPWR.n2571 VPWR.n2570 0.1685
R10574 VPWR.n2570 VPWR.n2569 0.1685
R10575 VPWR.n2569 VPWR.n2568 0.1685
R10576 VPWR.n2568 VPWR.n2567 0.1685
R10577 VPWR.n2567 VPWR.n2566 0.1685
R10578 VPWR.n2566 VPWR.n2565 0.1685
R10579 VPWR.n2564 VPWR.n2563 0.1685
R10580 VPWR.n2563 VPWR.n2562 0.1685
R10581 VPWR.n2556 VPWR.n2555 0.1685
R10582 VPWR.n2555 VPWR.n2554 0.1685
R10583 VPWR.n2554 VPWR.n2553 0.1685
R10584 VPWR.n2553 VPWR.n2552 0.1685
R10585 VPWR.n2552 VPWR.n2551 0.1685
R10586 VPWR.n2551 VPWR.n2550 0.1685
R10587 VPWR.n2550 VPWR.n2549 0.1685
R10588 VPWR.n2548 VPWR.n2547 0.1685
R10589 VPWR.n2547 VPWR.n2546 0.1685
R10590 VPWR.n2546 VPWR.n2545 0.1685
R10591 VPWR.n2545 VPWR.n2544 0.1685
R10592 VPWR.n2543 VPWR.n2542 0.1685
R10593 VPWR.n2542 VPWR.n0 0.1685
R10594 VPWR.n20 VPWR.n19 0.1685
R10595 VPWR.n3813 VPWR.n3812 0.1685
R10596 VPWR.n3812 VPWR.n3811 0.1685
R10597 VPWR.n3811 VPWR.n3810 0.1685
R10598 VPWR.n3810 VPWR.n3809 0.1685
R10599 VPWR.n3809 VPWR.n3808 0.1685
R10600 VPWR.n3808 VPWR.n3807 0.1685
R10601 VPWR.n3807 VPWR.n3806 0.1685
R10602 VPWR.n3805 VPWR.n3804 0.1685
R10603 VPWR.n3804 VPWR.n3803 0.1685
R10604 VPWR.n3803 VPWR.n3802 0.1685
R10605 VPWR.n3802 VPWR.n3801 0.1685
R10606 VPWR.n3796 VPWR.n3795 0.1685
R10607 VPWR.n3795 VPWR.n3794 0.1685
R10608 VPWR.n3794 VPWR.n3793 0.1685
R10609 VPWR.n3793 VPWR.n3792 0.1685
R10610 VPWR.n3792 VPWR.n3791 0.1685
R10611 VPWR.n3791 VPWR.n3790 0.1685
R10612 VPWR.n3790 VPWR.n3789 0.1685
R10613 VPWR.n3788 VPWR.n3787 0.1685
R10614 VPWR.n3787 VPWR.n3786 0.1685
R10615 VPWR.n3786 VPWR.n3785 0.1685
R10616 VPWR.n3785 VPWR.n3784 0.1685
R10617 VPWR.n3784 VPWR.n3783 0.1685
R10618 VPWR.n3783 VPWR.n3782 0.1685
R10619 VPWR.n83 VPWR.n62 0.1685
R10620 VPWR.n3752 VPWR.n3751 0.1685
R10621 VPWR.n3751 VPWR.n3750 0.1685
R10622 VPWR.n3750 VPWR.n3749 0.1685
R10623 VPWR.n3749 VPWR.n3748 0.1685
R10624 VPWR.n3748 VPWR.n3747 0.1685
R10625 VPWR.n3746 VPWR.n3745 0.1685
R10626 VPWR.n3745 VPWR.n3744 0.1685
R10627 VPWR.n3744 VPWR.n3743 0.1685
R10628 VPWR.n3743 VPWR.n3742 0.1685
R10629 VPWR.n3742 VPWR.n3741 0.1685
R10630 VPWR.n3741 VPWR.n3740 0.1685
R10631 VPWR.n3736 VPWR.n3735 0.1685
R10632 VPWR.n3735 VPWR.n3734 0.1685
R10633 VPWR.n3734 VPWR.n3733 0.1685
R10634 VPWR.n3733 VPWR.n3732 0.1685
R10635 VPWR.n3732 VPWR.n3731 0.1685
R10636 VPWR.n3731 VPWR.n3730 0.1685
R10637 VPWR.n3730 VPWR.n3729 0.1685
R10638 VPWR.n3728 VPWR.n3727 0.1685
R10639 VPWR.n3727 VPWR.n3726 0.1685
R10640 VPWR.n3726 VPWR.n3725 0.1685
R10641 VPWR.n3725 VPWR.n3724 0.1685
R10642 VPWR.n3724 VPWR.n3723 0.1685
R10643 VPWR.n3723 VPWR.n3722 0.1685
R10644 VPWR.n3722 VPWR.n3721 0.1685
R10645 VPWR.n3316 VPWR.n122 0.167
R10646 VPWR.n977 VPWR 0.1655
R10647 VPWR.n2911 VPWR.n2910 0.1655
R10648 VPWR.n869 VPWR 0.16475
R10649 VPWR.n1768 VPWR.n1767 0.16475
R10650 VPWR.n1220 VPWR.n1219 0.164
R10651 VPWR.n1246 VPWR.n1245 0.164
R10652 VPWR.n1695 VPWR.n1694 0.164
R10653 VPWR.n1180 VPWR.n1179 0.164
R10654 VPWR.n1146 VPWR.n1145 0.164
R10655 VPWR.n1967 VPWR.n1966 0.164
R10656 VPWR.n1918 VPWR.n1917 0.164
R10657 VPWR VPWR.n1604 0.16325
R10658 VPWR VPWR.n3336 0.1625
R10659 VPWR.n1697 VPWR 0.1625
R10660 VPWR.n1747 VPWR.n1746 0.1625
R10661 VPWR.n1751 VPWR.n1750 0.1625
R10662 VPWR.n1793 VPWR 0.1625
R10663 VPWR.n3216 VPWR 0.1625
R10664 VPWR.n1098 VPWR 0.1625
R10665 VPWR.n1837 VPWR.n1836 0.1625
R10666 VPWR.n2004 VPWR.n1926 0.1625
R10667 VPWR.n2053 VPWR.n2006 0.1625
R10668 VPWR VPWR.n2793 0.1625
R10669 VPWR.n1924 VPWR.n360 0.1625
R10670 VPWR VPWR.n1486 0.161
R10671 VPWR.n997 VPWR.n996 0.161
R10672 VPWR.n1815 VPWR.n699 0.161
R10673 VPWR.n578 VPWR.n577 0.161
R10674 VPWR VPWR.n131 0.1595
R10675 VPWR.n3226 VPWR.n3225 0.1595
R10676 VPWR VPWR.n3239 0.1595
R10677 VPWR VPWR.n3297 0.1595
R10678 VPWR.n1187 VPWR.n1186 0.1595
R10679 VPWR.n1746 VPWR.n1745 0.1595
R10680 VPWR.n1752 VPWR.n1751 0.1595
R10681 VPWR.n1109 VPWR.n1108 0.1595
R10682 VPWR.n693 VPWR 0.1595
R10683 VPWR VPWR.n663 0.1595
R10684 VPWR.n1950 VPWR.n1949 0.1595
R10685 VPWR.n2912 VPWR 0.1595
R10686 VPWR.n1871 VPWR 0.1595
R10687 VPWR VPWR.n419 0.1595
R10688 VPWR.n1814 VPWR.n1813 0.15875
R10689 VPWR.n1687 VPWR 0.158
R10690 VPWR.n1297 VPWR 0.15725
R10691 VPWR.n3294 VPWR 0.15725
R10692 VPWR.n1771 VPWR.n1770 0.15725
R10693 VPWR.n660 VPWR 0.15725
R10694 VPWR VPWR.n1477 0.1565
R10695 VPWR VPWR.n1483 0.1565
R10696 VPWR.n1443 VPWR 0.1565
R10697 VPWR.n1436 VPWR 0.1565
R10698 VPWR VPWR.n1316 0.1565
R10699 VPWR.n1315 VPWR 0.1565
R10700 VPWR.n1313 VPWR 0.1565
R10701 VPWR.n1281 VPWR 0.1565
R10702 VPWR VPWR.n818 0.1565
R10703 VPWR.n1650 VPWR 0.1565
R10704 VPWR.n898 VPWR 0.1565
R10705 VPWR.n3348 VPWR 0.1565
R10706 VPWR.n3343 VPWR.n3342 0.1565
R10707 VPWR.n3371 VPWR 0.1565
R10708 VPWR.n1683 VPWR 0.1565
R10709 VPWR.n3288 VPWR.n3287 0.1565
R10710 VPWR.n2835 VPWR 0.1565
R10711 VPWR.n2803 VPWR 0.1565
R10712 VPWR.n2802 VPWR.n2801 0.1565
R10713 VPWR.n2800 VPWR 0.1565
R10714 VPWR VPWR.n1848 0.1565
R10715 VPWR VPWR.n593 0.1565
R10716 VPWR VPWR.n406 0.1565
R10717 VPWR VPWR.n2927 0.1565
R10718 VPWR.n1596 VPWR 0.15575
R10719 VPWR VPWR.n1575 0.15575
R10720 VPWR.n1435 VPWR 0.15575
R10721 VPWR VPWR.n1425 0.15575
R10722 VPWR.n1319 VPWR 0.15575
R10723 VPWR.n1287 VPWR 0.15575
R10724 VPWR.n1657 VPWR 0.15575
R10725 VPWR VPWR.n888 0.15575
R10726 VPWR VPWR.n1842 0.15575
R10727 VPWR.n1859 VPWR 0.15575
R10728 VPWR VPWR.n590 0.15575
R10729 VPWR VPWR.n431 0.15575
R10730 VPWR.n403 VPWR 0.15575
R10731 VPWR.n398 VPWR 0.15575
R10732 VPWR.n2935 VPWR 0.15575
R10733 VPWR.n1074 VPWR 0.155
R10734 VPWR VPWR.n1479 0.155
R10735 VPWR VPWR.n1632 0.155
R10736 VPWR VPWR.n1622 0.155
R10737 VPWR.n812 VPWR 0.155
R10738 VPWR.n3192 VPWR 0.155
R10739 VPWR VPWR.n1446 0.1535
R10740 VPWR.n1607 VPWR.n1017 0.1535
R10741 VPWR.n1295 VPWR.n1294 0.1535
R10742 VPWR.n764 VPWR.n763 0.1535
R10743 VPWR.n1777 VPWR.n1776 0.1535
R10744 VPWR.n689 VPWR 0.1535
R10745 VPWR.n1465 VPWR 0.15275
R10746 VPWR.n1270 VPWR 0.15275
R10747 VPWR.n1693 VPWR 0.15275
R10748 VPWR.n1083 VPWR 0.15275
R10749 VPWR.n1977 VPWR 0.15275
R10750 VPWR VPWR.n2134 0.15275
R10751 VPWR VPWR.n2729 0.15275
R10752 VPWR.n2693 VPWR 0.15275
R10753 VPWR.n1870 VPWR 0.15275
R10754 VPWR.n1885 VPWR 0.15275
R10755 VPWR.n443 VPWR 0.15275
R10756 VPWR VPWR.n1010 0.152
R10757 VPWR.n866 VPWR 0.152
R10758 VPWR VPWR.n1196 0.152
R10759 VPWR.n1100 VPWR.n1099 0.152
R10760 VPWR.n574 VPWR 0.152
R10761 VPWR VPWR.n1595 0.15125
R10762 VPWR.n1576 VPWR 0.15125
R10763 VPWR VPWR.n1318 0.15125
R10764 VPWR VPWR.n1290 0.15125
R10765 VPWR.n1672 VPWR 0.15125
R10766 VPWR.n889 VPWR 0.15125
R10767 VPWR.n790 VPWR 0.15125
R10768 VPWR.n784 VPWR 0.15125
R10769 VPWR VPWR.n1768 0.15125
R10770 VPWR.n591 VPWR 0.15125
R10771 VPWR VPWR.n567 0.15125
R10772 VPWR.n432 VPWR 0.15125
R10773 VPWR VPWR.n402 0.15125
R10774 VPWR VPWR.n2934 0.15125
R10775 VPWR.n816 VPWR 0.1505
R10776 VPWR.n1760 VPWR 0.1505
R10777 VPWR.n1609 VPWR 0.14975
R10778 VPWR.n1366 VPWR.n1365 0.149
R10779 VPWR.n1415 VPWR.n1414 0.1475
R10780 VPWR.n1620 VPWR.n1619 0.1475
R10781 VPWR.n780 VPWR 0.1475
R10782 VPWR.n774 VPWR.n773 0.1475
R10783 VPWR.n3292 VPWR.n3291 0.1475
R10784 VPWR VPWR.n692 0.1475
R10785 VPWR.n2344 VPWR.n2343 0.1475
R10786 VPWR.n2670 VPWR.n2669 0.1475
R10787 VPWR VPWR.n1852 0.1475
R10788 VPWR.n420 VPWR 0.1475
R10789 VPWR.n2602 VPWR.n258 0.1475
R10790 VPWR.n2599 VPWR.n260 0.1475
R10791 VPWR.n791 VPWR.n790 0.14675
R10792 VPWR.n1072 VPWR 0.146
R10793 VPWR VPWR.n1475 0.146
R10794 VPWR.n1337 VPWR 0.146
R10795 VPWR.n875 VPWR.n874 0.146
R10796 VPWR VPWR.n3349 0.146
R10797 VPWR VPWR.n1705 0.146
R10798 VPWR VPWR.n3311 0.146
R10799 VPWR.n3302 VPWR 0.146
R10800 VPWR.n1815 VPWR.n1814 0.146
R10801 VPWR VPWR.n600 0.146
R10802 VPWR.n577 VPWR.n576 0.146
R10803 VPWR VPWR.n2946 0.146
R10804 VPWR.n1619 VPWR 0.14525
R10805 VPWR.n1332 VPWR.n1331 0.14525
R10806 VPWR.n695 VPWR 0.14525
R10807 VPWR.n1414 VPWR.n1413 0.1445
R10808 VPWR.n905 VPWR.n904 0.1445
R10809 VPWR.n773 VPWR.n772 0.1445
R10810 VPWR.n771 VPWR.n770 0.1445
R10811 VPWR.n3237 VPWR.n3236 0.1445
R10812 VPWR.n3289 VPWR 0.1445
R10813 VPWR.n1138 VPWR.n1137 0.1445
R10814 VPWR.n678 VPWR.n677 0.1445
R10815 VPWR.n643 VPWR.n642 0.1445
R10816 VPWR.n1947 VPWR.n1946 0.1445
R10817 VPWR.n2718 VPWR.n2717 0.1445
R10818 VPWR.n1874 VPWR.n1873 0.1445
R10819 VPWR.n555 VPWR.n554 0.1445
R10820 VPWR.n1890 VPWR.n1889 0.1445
R10821 VPWR.n3016 VPWR.n3015 0.1445
R10822 VPWR.n1946 VPWR 0.14375
R10823 VPWR VPWR.n1078 0.143
R10824 VPWR VPWR.n1356 0.143
R10825 VPWR.n1362 VPWR 0.143
R10826 VPWR.n1365 VPWR 0.143
R10827 VPWR VPWR.n1465 0.143
R10828 VPWR.n1274 VPWR 0.143
R10829 VPWR VPWR.n1273 0.143
R10830 VPWR VPWR.n1270 0.143
R10831 VPWR VPWR.n1342 0.143
R10832 VPWR.n1339 VPWR 0.143
R10833 VPWR VPWR.n1338 0.143
R10834 VPWR VPWR.n1332 0.143
R10835 VPWR.n1228 VPWR 0.143
R10836 VPWR.n1227 VPWR 0.143
R10837 VPWR VPWR.n1222 0.143
R10838 VPWR VPWR.n1218 0.143
R10839 VPWR VPWR.n1693 0.143
R10840 VPWR.n800 VPWR.n799 0.143
R10841 VPWR.n785 VPWR 0.143
R10842 VPWR.n1167 VPWR 0.143
R10843 VPWR VPWR.n1166 0.143
R10844 VPWR.n1163 VPWR 0.143
R10845 VPWR VPWR.n1162 0.143
R10846 VPWR VPWR.n1214 0.143
R10847 VPWR VPWR.n1209 0.143
R10848 VPWR VPWR.n1208 0.143
R10849 VPWR.n1207 VPWR 0.143
R10850 VPWR.n1206 VPWR 0.143
R10851 VPWR.n1198 VPWR 0.143
R10852 VPWR.n1188 VPWR 0.143
R10853 VPWR VPWR.n1184 0.143
R10854 VPWR.n1179 VPWR 0.143
R10855 VPWR.n1086 VPWR 0.143
R10856 VPWR VPWR.n1083 0.143
R10857 VPWR.n1139 VPWR 0.143
R10858 VPWR VPWR.n1125 0.143
R10859 VPWR.n1969 VPWR 0.143
R10860 VPWR.n1966 VPWR 0.143
R10861 VPWR.n1965 VPWR 0.143
R10862 VPWR VPWR.n2716 0.143
R10863 VPWR VPWR.n2697 0.143
R10864 VPWR.n508 VPWR 0.143
R10865 VPWR.n507 VPWR 0.143
R10866 VPWR VPWR.n502 0.143
R10867 VPWR VPWR.n501 0.143
R10868 VPWR VPWR.n499 0.143
R10869 VPWR.n1880 VPWR 0.143
R10870 VPWR.n1875 VPWR 0.143
R10871 VPWR VPWR.n1870 0.143
R10872 VPWR VPWR.n1915 0.143
R10873 VPWR.n453 VPWR 0.143
R10874 VPWR.n452 VPWR 0.143
R10875 VPWR VPWR.n447 0.143
R10876 VPWR VPWR.n446 0.143
R10877 VPWR VPWR.n443 0.143
R10878 VPWR.n1664 VPWR 0.1415
R10879 VPWR.n3229 VPWR.n3228 0.1415
R10880 VPWR VPWR.n1812 0.1415
R10881 VPWR.n1844 VPWR.n603 0.1415
R10882 VPWR.n584 VPWR.n583 0.1415
R10883 VPWR.n1082 VPWR.n1081 0.14
R10884 VPWR.n1140 VPWR.n1139 0.14
R10885 VPWR.n1987 VPWR.n1986 0.14
R10886 VPWR.n1985 VPWR.n1984 0.14
R10887 VPWR.n2716 VPWR.n2715 0.14
R10888 VPWR.n2720 VPWR.n2719 0.14
R10889 VPWR.n2722 VPWR.n2721 0.14
R10890 VPWR.n2075 VPWR.n2074 0.14
R10891 VPWR.n2073 VPWR.n2072 0.14
R10892 VPWR.n2071 VPWR.n2070 0.14
R10893 VPWR.n2069 VPWR.n2068 0.14
R10894 VPWR.n2067 VPWR.n197 0.14
R10895 VPWR.n2706 VPWR.n2705 0.14
R10896 VPWR.n493 VPWR.n492 0.14
R10897 VPWR.n495 VPWR.n494 0.14
R10898 VPWR.n1077 VPWR.n1076 0.1385
R10899 VPWR.n1483 VPWR.n1482 0.1385
R10900 VPWR.n1490 VPWR.n1489 0.1385
R10901 VPWR.n1506 VPWR.n1505 0.1385
R10902 VPWR.n1599 VPWR.n1598 0.1385
R10903 VPWR.n1593 VPWR.n1592 0.1385
R10904 VPWR.n1545 VPWR.n1544 0.1385
R10905 VPWR.n1360 VPWR.n1359 0.1385
R10906 VPWR.n1637 VPWR.n1636 0.1385
R10907 VPWR VPWR.n1625 0.1385
R10908 VPWR.n976 VPWR.n975 0.1385
R10909 VPWR.n974 VPWR.n973 0.1385
R10910 VPWR.n3386 VPWR.n3385 0.1385
R10911 VPWR.n3388 VPWR.n3387 0.1385
R10912 VPWR.n3398 VPWR.n3397 0.1385
R10913 VPWR.n3415 VPWR.n3414 0.1385
R10914 VPWR.n1341 VPWR.n1340 0.1385
R10915 VPWR.n1655 VPWR.n1654 0.1385
R10916 VPWR VPWR.n875 0.1385
R10917 VPWR.n3325 VPWR.n3324 0.1385
R10918 VPWR VPWR.n1221 0.1385
R10919 VPWR VPWR.n1696 0.1385
R10920 VPWR.n3290 VPWR.n3289 0.1385
R10921 VPWR.n1211 VPWR.n1210 0.1385
R10922 VPWR.n1203 VPWR 0.1385
R10923 VPWR.n1745 VPWR.n1744 0.1385
R10924 VPWR.n3175 VPWR.n3174 0.1385
R10925 VPWR VPWR.n1119 0.1385
R10926 VPWR.n1102 VPWR.n1101 0.1385
R10927 VPWR.n665 VPWR.n664 0.1385
R10928 VPWR VPWR.n657 0.1385
R10929 VPWR.n648 VPWR.n647 0.1385
R10930 VPWR VPWR.n643 0.1385
R10931 VPWR.n3115 VPWR.n3114 0.1385
R10932 VPWR.n3144 VPWR.n3143 0.1385
R10933 VPWR.n1972 VPWR.n1971 0.1385
R10934 VPWR.n1962 VPWR 0.1385
R10935 VPWR VPWR.n1950 0.1385
R10936 VPWR.n2845 VPWR 0.1385
R10937 VPWR.n2860 VPWR.n2859 0.1385
R10938 VPWR.n2109 VPWR.n2108 0.1385
R10939 VPWR.n2141 VPWR.n2140 0.1385
R10940 VPWR.n2167 VPWR.n2166 0.1385
R10941 VPWR.n304 VPWR.n303 0.1385
R10942 VPWR.n331 VPWR.n330 0.1385
R10943 VPWR.n2268 VPWR.n2267 0.1385
R10944 VPWR.n2250 VPWR.n2249 0.1385
R10945 VPWR.n2308 VPWR.n2307 0.1385
R10946 VPWR.n2290 VPWR.n2289 0.1385
R10947 VPWR.n2193 VPWR.n2192 0.1385
R10948 VPWR.n2219 VPWR.n2218 0.1385
R10949 VPWR.n2368 VPWR.n2367 0.1385
R10950 VPWR.n2358 VPWR.n2357 0.1385
R10951 VPWR.n2349 VPWR.n2348 0.1385
R10952 VPWR.n2339 VPWR.n2338 0.1385
R10953 VPWR.n2051 VPWR.n2050 0.1385
R10954 VPWR.n2033 VPWR.n2032 0.1385
R10955 VPWR.n2728 VPWR 0.1385
R10956 VPWR.n2746 VPWR.n2745 0.1385
R10957 VPWR.n2826 VPWR.n2825 0.1385
R10958 VPWR.n2795 VPWR.n2794 0.1385
R10959 VPWR.n2779 VPWR.n2778 0.1385
R10960 VPWR.n2092 VPWR.n2091 0.1385
R10961 VPWR.n2685 VPWR.n2684 0.1385
R10962 VPWR.n2682 VPWR.n2681 0.1385
R10963 VPWR.n2664 VPWR.n2663 0.1385
R10964 VPWR.n2655 VPWR.n2654 0.1385
R10965 VPWR.n2653 VPWR.n2652 0.1385
R10966 VPWR.n252 VPWR.n251 0.1385
R10967 VPWR.n236 VPWR.n235 0.1385
R10968 VPWR.n468 VPWR 0.1385
R10969 VPWR VPWR.n469 0.1385
R10970 VPWR.n492 VPWR 0.1385
R10971 VPWR.n568 VPWR 0.1385
R10972 VPWR.n554 VPWR 0.1385
R10973 VPWR.n3027 VPWR.n3026 0.1385
R10974 VPWR.n3034 VPWR 0.1385
R10975 VPWR.n3055 VPWR.n3054 0.1385
R10976 VPWR.n3101 VPWR.n3100 0.1385
R10977 VPWR.n3083 VPWR.n3082 0.1385
R10978 VPWR.n361 VPWR 0.1385
R10979 VPWR.n369 VPWR.n368 0.1385
R10980 VPWR VPWR.n1910 0.1385
R10981 VPWR VPWR.n1904 0.1385
R10982 VPWR.n445 VPWR.n444 0.1385
R10983 VPWR VPWR.n399 0.1385
R10984 VPWR.n3013 VPWR.n3012 0.1385
R10985 VPWR.n2997 VPWR.n2996 0.1385
R10986 VPWR.n2987 VPWR.n2986 0.1385
R10987 VPWR.n2978 VPWR.n2977 0.1385
R10988 VPWR.n2968 VPWR.n2967 0.1385
R10989 VPWR.n2461 VPWR.n2460 0.1385
R10990 VPWR.n2479 VPWR.n2478 0.1385
R10991 VPWR.n2499 VPWR.n2498 0.1385
R10992 VPWR.n2490 VPWR.n2489 0.1385
R10993 VPWR.n2604 VPWR.n2603 0.1385
R10994 VPWR.n2619 VPWR.n2618 0.1385
R10995 VPWR.n2641 VPWR.n2640 0.1385
R10996 VPWR.n2632 VPWR.n2631 0.1385
R10997 VPWR.n3827 VPWR.n3826 0.1385
R10998 VPWR.n48 VPWR.n47 0.1385
R10999 VPWR.n56 VPWR.n38 0.1385
R11000 VPWR.n3767 VPWR.n3766 0.1385
R11001 VPWR.n3758 VPWR.n3757 0.1385
R11002 VPWR.n3694 VPWR.n3693 0.1385
R11003 VPWR.n3706 VPWR.n3705 0.1385
R11004 VPWR.n2445 VPWR.n2444 0.1385
R11005 VPWR.n2437 VPWR.n2436 0.1385
R11006 VPWR.n2506 VPWR.n2505 0.1385
R11007 VPWR.n2516 VPWR.n2515 0.1385
R11008 VPWR.n2534 VPWR.n2533 0.1385
R11009 VPWR.n2597 VPWR.n2596 0.1385
R11010 VPWR.n2590 VPWR.n2589 0.1385
R11011 VPWR.n2584 VPWR.n2583 0.1385
R11012 VPWR.n2573 VPWR.n2572 0.1385
R11013 VPWR.n2561 VPWR.n2560 0.1385
R11014 VPWR.n2557 VPWR.n2556 0.1385
R11015 VPWR.n18 VPWR.n17 0.1385
R11016 VPWR.n30 VPWR.n29 0.1385
R11017 VPWR.n3800 VPWR.n3799 0.1385
R11018 VPWR.n3797 VPWR.n3796 0.1385
R11019 VPWR.n3780 VPWR.n3779 0.1385
R11020 VPWR.n72 VPWR.n71 0.1385
R11021 VPWR.n74 VPWR.n73 0.1385
R11022 VPWR.n84 VPWR.n83 0.1385
R11023 VPWR.n3739 VPWR.n3738 0.1385
R11024 VPWR.n1425 VPWR 0.13775
R11025 VPWR VPWR.n574 0.13775
R11026 VPWR VPWR.n1481 0.137
R11027 VPWR.n1513 VPWR.n1512 0.137
R11028 VPWR.n1591 VPWR.n1590 0.137
R11029 VPWR.n1461 VPWR 0.137
R11030 VPWR.n1704 VPWR 0.137
R11031 VPWR.n1710 VPWR.n726 0.137
R11032 VPWR.n1842 VPWR 0.137
R11033 VPWR.n1881 VPWR.n457 0.137
R11034 VPWR.n599 VPWR 0.137
R11035 VPWR.n3818 VPWR.n3817 0.137
R11036 VPWR.n3814 VPWR.n9 0.137
R11037 VPWR VPWR.n1427 0.13625
R11038 VPWR.n1044 VPWR.n1043 0.1355
R11039 VPWR.n3341 VPWR.n107 0.1355
R11040 VPWR.n3372 VPWR.n3371 0.1355
R11041 VPWR.n781 VPWR.n780 0.1355
R11042 VPWR.n1716 VPWR 0.1355
R11043 VPWR.n2905 VPWR.n2904 0.1355
R11044 VPWR.n2377 VPWR.n2376 0.1355
R11045 VPWR.n477 VPWR.n476 0.1355
R11046 VPWR.n481 VPWR.n480 0.1355
R11047 VPWR.n485 VPWR.n484 0.1355
R11048 VPWR.n1876 VPWR.n1875 0.1355
R11049 VPWR.n2971 VPWR.n2970 0.1355
R11050 VPWR.n2467 VPWR.n2466 0.1355
R11051 VPWR.n589 VPWR 0.134
R11052 VPWR VPWR.n1834 0.13325
R11053 VPWR.n777 VPWR.n776 0.1325
R11054 VPWR.n1200 VPWR.n1199 0.1325
R11055 VPWR.n1189 VPWR.n1188 0.1325
R11056 VPWR.n3200 VPWR.n3199 0.1325
R11057 VPWR VPWR.n690 0.1325
R11058 VPWR.n1433 VPWR.n1432 0.13175
R11059 VPWR.n3446 VPWR 0.131
R11060 VPWR.n3461 VPWR 0.131
R11061 VPWR.n3476 VPWR 0.131
R11062 VPWR.n3491 VPWR 0.131
R11063 VPWR.n3506 VPWR 0.131
R11064 VPWR.n3521 VPWR 0.131
R11065 VPWR.n3536 VPWR 0.131
R11066 VPWR.n3551 VPWR 0.131
R11067 VPWR.n3566 VPWR 0.131
R11068 VPWR.n3581 VPWR 0.131
R11069 VPWR.n3596 VPWR 0.131
R11070 VPWR.n3611 VPWR 0.131
R11071 VPWR.n3626 VPWR 0.131
R11072 VPWR.n3641 VPWR 0.131
R11073 VPWR.n3656 VPWR 0.131
R11074 VPWR.n3671 VPWR 0.131
R11075 VPWR VPWR.n1054 0.131
R11076 VPWR.n1476 VPWR 0.131
R11077 VPWR VPWR.n1597 0.131
R11078 VPWR.n1533 VPWR 0.131
R11079 VPWR VPWR.n1561 0.131
R11080 VPWR VPWR.n1552 0.131
R11081 VPWR VPWR.n1443 0.131
R11082 VPWR VPWR.n1417 0.131
R11083 VPWR.n996 VPWR.n995 0.131
R11084 VPWR VPWR.n989 0.131
R11085 VPWR VPWR.n1275 0.131
R11086 VPWR VPWR.n1330 0.131
R11087 VPWR VPWR.n1302 0.131
R11088 VPWR VPWR.n905 0.131
R11089 VPWR VPWR.n893 0.131
R11090 VPWR VPWR.n861 0.131
R11091 VPWR VPWR.n1238 0.131
R11092 VPWR VPWR.n728 0.131
R11093 VPWR VPWR.n1685 0.131
R11094 VPWR VPWR.n769 0.131
R11095 VPWR VPWR.n3246 0.131
R11096 VPWR VPWR.n3309 0.131
R11097 VPWR VPWR.n3275 0.131
R11098 VPWR VPWR.n1178 0.131
R11099 VPWR.n1722 VPWR 0.131
R11100 VPWR VPWR.n1152 0.131
R11101 VPWR VPWR.n1975 0.131
R11102 VPWR.n2833 VPWR 0.131
R11103 VPWR.n2839 VPWR 0.131
R11104 VPWR VPWR.n2889 0.131
R11105 VPWR.n350 VPWR 0.131
R11106 VPWR.n287 VPWR 0.131
R11107 VPWR VPWR.n282 0.131
R11108 VPWR VPWR.n2017 0.131
R11109 VPWR VPWR.n2784 0.131
R11110 VPWR VPWR.n2063 0.131
R11111 VPWR VPWR.n2691 0.131
R11112 VPWR VPWR.n500 0.131
R11113 VPWR VPWR.n597 0.131
R11114 VPWR.n576 VPWR.n575 0.131
R11115 VPWR VPWR.n367 0.131
R11116 VPWR VPWR.n424 0.131
R11117 VPWR.n3702 VPWR 0.131
R11118 VPWR VPWR.n2425 0.131
R11119 VPWR.n1434 VPWR.n1433 0.13025
R11120 VPWR.n1351 VPWR.n1350 0.1295
R11121 VPWR.n3227 VPWR 0.1295
R11122 VPWR.n1112 VPWR.n1111 0.1295
R11123 VPWR.n562 VPWR.n561 0.1295
R11124 VPWR.n1730 VPWR.n1729 0.128
R11125 VPWR.n3450 VPWR 0.12725
R11126 VPWR.n3465 VPWR 0.12725
R11127 VPWR.n3480 VPWR 0.12725
R11128 VPWR.n3495 VPWR 0.12725
R11129 VPWR.n3510 VPWR 0.12725
R11130 VPWR.n3525 VPWR 0.12725
R11131 VPWR.n3540 VPWR 0.12725
R11132 VPWR.n3555 VPWR 0.12725
R11133 VPWR.n3570 VPWR 0.12725
R11134 VPWR.n3585 VPWR 0.12725
R11135 VPWR.n3600 VPWR 0.12725
R11136 VPWR.n3615 VPWR 0.12725
R11137 VPWR.n3630 VPWR 0.12725
R11138 VPWR.n3645 VPWR 0.12725
R11139 VPWR.n3660 VPWR 0.12725
R11140 VPWR.n3675 VPWR 0.12725
R11141 VPWR VPWR.n1509 0.12725
R11142 VPWR.n1521 VPWR 0.12725
R11143 VPWR.n1582 VPWR 0.12725
R11144 VPWR.n1570 VPWR 0.12725
R11145 VPWR.n1553 VPWR 0.12725
R11146 VPWR.n1468 VPWR 0.12725
R11147 VPWR.n1460 VPWR 0.12725
R11148 VPWR.n1439 VPWR 0.12725
R11149 VPWR.n1424 VPWR 0.12725
R11150 VPWR.n1005 VPWR 0.12725
R11151 VPWR.n907 VPWR 0.12725
R11152 VPWR.n3369 VPWR 0.12725
R11153 VPWR.n1240 VPWR 0.12725
R11154 VPWR.n1686 VPWR 0.12725
R11155 VPWR.n3312 VPWR 0.12725
R11156 VPWR.n3301 VPWR 0.12725
R11157 VPWR.n3218 VPWR 0.12725
R11158 VPWR.n165 VPWR 0.12725
R11159 VPWR.n1141 VPWR 0.12725
R11160 VPWR.n1107 VPWR 0.12725
R11161 VPWR.n1829 VPWR 0.12725
R11162 VPWR.n3153 VPWR 0.12725
R11163 VPWR.n2002 VPWR 0.12725
R11164 VPWR.n1992 VPWR 0.12725
R11165 VPWR VPWR.n2832 0.12725
R11166 VPWR.n2916 VPWR 0.12725
R11167 VPWR VPWR.n2126 0.12725
R11168 VPWR.n2176 VPWR 0.12725
R11169 VPWR.n340 VPWR 0.12725
R11170 VPWR.n2228 VPWR 0.12725
R11171 VPWR VPWR.n2712 0.12725
R11172 VPWR.n2808 VPWR 0.12725
R11173 VPWR.n2759 VPWR 0.12725
R11174 VPWR.n2084 VPWR 0.12725
R11175 VPWR.n1877 VPWR 0.12725
R11176 VPWR.n1861 VPWR 0.12725
R11177 VPWR.n564 VPWR.n563 0.12725
R11178 VPWR.n3064 VPWR 0.12725
R11179 VPWR.n2950 VPWR 0.12725
R11180 VPWR.n1421 VPWR.n1420 0.1265
R11181 VPWR.n1634 VPWR.n1633 0.1265
R11182 VPWR.n1668 VPWR 0.1265
R11183 VPWR.n3342 VPWR 0.1265
R11184 VPWR.n782 VPWR.n781 0.1265
R11185 VPWR.n3254 VPWR 0.1265
R11186 VPWR.n1099 VPWR.n1098 0.1265
R11187 VPWR.n645 VPWR.n644 0.1265
R11188 VPWR.n2924 VPWR.n2923 0.12575
R11189 VPWR.n3240 VPWR 0.12425
R11190 VPWR.n2666 VPWR 0.12425
R11191 VPWR.n2523 VPWR 0.12425
R11192 VPWR.n2544 VPWR 0.12425
R11193 VPWR.n3782 VPWR 0.12425
R11194 VPWR.n1463 VPWR.n1462 0.1235
R11195 VPWR.n885 VPWR.n884 0.1235
R11196 VPWR.n877 VPWR.n876 0.1235
R11197 VPWR VPWR.n868 0.1235
R11198 VPWR.n1703 VPWR.n1702 0.1235
R11199 VPWR.n408 VPWR.n407 0.1235
R11200 VPWR.n789 VPWR.n788 0.12275
R11201 VPWR VPWR.n3445 0.122
R11202 VPWR VPWR.n3460 0.122
R11203 VPWR VPWR.n3475 0.122
R11204 VPWR VPWR.n3490 0.122
R11205 VPWR VPWR.n3505 0.122
R11206 VPWR VPWR.n3520 0.122
R11207 VPWR VPWR.n3535 0.122
R11208 VPWR VPWR.n3550 0.122
R11209 VPWR VPWR.n3565 0.122
R11210 VPWR VPWR.n3580 0.122
R11211 VPWR VPWR.n3595 0.122
R11212 VPWR VPWR.n3610 0.122
R11213 VPWR VPWR.n3625 0.122
R11214 VPWR VPWR.n3640 0.122
R11215 VPWR VPWR.n3655 0.122
R11216 VPWR VPWR.n3670 0.122
R11217 VPWR.n1428 VPWR 0.122
R11218 VPWR.n1821 VPWR.n1820 0.122
R11219 VPWR.n1979 VPWR 0.122
R11220 VPWR VPWR.n2838 0.122
R11221 VPWR.n2890 VPWR 0.122
R11222 VPWR VPWR.n349 0.122
R11223 VPWR VPWR.n286 0.122
R11224 VPWR.n283 VPWR 0.122
R11225 VPWR.n2785 VPWR 0.122
R11226 VPWR VPWR.n489 0.122
R11227 VPWR.n425 VPWR 0.122
R11228 VPWR.n894 VPWR 0.12125
R11229 VPWR VPWR.n1804 0.12125
R11230 VPWR.n402 VPWR.n401 0.12125
R11231 VPWR.n2945 VPWR 0.12125
R11232 VPWR.n1079 VPWR 0.1205
R11233 VPWR VPWR.n1347 0.1205
R11234 VPWR VPWR.n1663 0.1205
R11235 VPWR.n3336 VPWR.n3335 0.1205
R11236 VPWR VPWR.n3227 0.1205
R11237 VPWR.n3300 VPWR.n3299 0.1205
R11238 VPWR.n1215 VPWR 0.1205
R11239 VPWR.n1794 VPWR.n1793 0.1205
R11240 VPWR.n3217 VPWR.n3216 0.1205
R11241 VPWR.n219 VPWR.n218 0.1205
R11242 VPWR.n3836 VPWR.n3835 0.1205
R11243 VPWR.n3839 VPWR.n2 0.1205
R11244 VPWR VPWR.n1423 0.11975
R11245 VPWR VPWR.n3406 0.11975
R11246 VPWR VPWR.n3424 0.11975
R11247 VPWR.n2674 VPWR 0.11975
R11248 VPWR.n244 VPWR 0.11975
R11249 VPWR.n226 VPWR 0.11975
R11250 VPWR.n1856 VPWR.n1855 0.11975
R11251 VPWR VPWR.n2513 0.11975
R11252 VPWR.n2526 VPWR 0.11975
R11253 VPWR.n2565 VPWR 0.11975
R11254 VPWR.n2549 VPWR 0.11975
R11255 VPWR.n3806 VPWR 0.11975
R11256 VPWR.n3789 VPWR 0.11975
R11257 VPWR.n3747 VPWR 0.11975
R11258 VPWR.n3729 VPWR 0.11975
R11259 VPWR.n1285 VPWR.n1284 0.119
R11260 VPWR.n1426 VPWR 0.1175
R11261 VPWR.n1645 VPWR.n1644 0.1175
R11262 VPWR.n1217 VPWR 0.1175
R11263 VPWR.n1202 VPWR.n1201 0.1175
R11264 VPWR.n1961 VPWR.n1960 0.1175
R11265 VPWR.n467 VPWR.n466 0.1175
R11266 VPWR.n433 VPWR 0.1175
R11267 VPWR.n3775 VPWR.n38 0.1175
R11268 VPWR.n3779 VPWR.n3778 0.1175
R11269 VPWR VPWR.n906 0.11675
R11270 VPWR.n807 VPWR.n806 0.11675
R11271 VPWR.n3243 VPWR.n3242 0.11675
R11272 VPWR VPWR.n2909 0.11675
R11273 VPWR VPWR.n1311 0.116
R11274 VPWR.n1798 VPWR 0.11525
R11275 VPWR.n1076 VPWR 0.1145
R11276 VPWR VPWR.n1476 0.1145
R11277 VPWR.n1600 VPWR 0.1145
R11278 VPWR.n1597 VPWR 0.1145
R11279 VPWR.n1589 VPWR 0.1145
R11280 VPWR.n1581 VPWR 0.1145
R11281 VPWR VPWR.n1527 0.1145
R11282 VPWR VPWR.n1533 0.1145
R11283 VPWR.n1555 VPWR 0.1145
R11284 VPWR VPWR.n1041 0.1145
R11285 VPWR.n1042 VPWR 0.1145
R11286 VPWR.n1046 VPWR 0.1145
R11287 VPWR.n1050 VPWR 0.1145
R11288 VPWR.n1466 VPWR 0.1145
R11289 VPWR.n1464 VPWR 0.1145
R11290 VPWR.n1417 VPWR 0.1145
R11291 VPWR.n978 VPWR 0.1145
R11292 VPWR.n3378 VPWR 0.1145
R11293 VPWR VPWR.n3382 0.1145
R11294 VPWR VPWR.n3386 0.1145
R11295 VPWR.n1268 VPWR 0.1145
R11296 VPWR.n1343 VPWR 0.1145
R11297 VPWR VPWR.n1334 0.1145
R11298 VPWR.n1330 VPWR 0.1145
R11299 VPWR.n1309 VPWR.n1308 0.1145
R11300 VPWR.n1302 VPWR 0.1145
R11301 VPWR.n1283 VPWR 0.1145
R11302 VPWR.n1670 VPWR.n1669 0.1145
R11303 VPWR VPWR.n1658 0.1145
R11304 VPWR VPWR.n901 0.1145
R11305 VPWR.n899 VPWR 0.1145
R11306 VPWR VPWR.n3325 0.1145
R11307 VPWR.n3350 VPWR 0.1145
R11308 VPWR.n3345 VPWR 0.1145
R11309 VPWR.n3363 VPWR 0.1145
R11310 VPWR.n1262 VPWR 0.1145
R11311 VPWR VPWR.n1255 0.1145
R11312 VPWR.n1252 VPWR 0.1145
R11313 VPWR.n1238 VPWR 0.1145
R11314 VPWR.n1233 VPWR 0.1145
R11315 VPWR.n1231 VPWR 0.1145
R11316 VPWR.n1691 VPWR 0.1145
R11317 VPWR VPWR.n3238 0.1145
R11318 VPWR.n3247 VPWR 0.1145
R11319 VPWR.n3298 VPWR 0.1145
R11320 VPWR.n3293 VPWR 0.1145
R11321 VPWR VPWR.n1169 0.1145
R11322 VPWR VPWR.n1722 0.1145
R11323 VPWR VPWR.n1759 0.1145
R11324 VPWR.n1809 VPWR 0.1145
R11325 VPWR.n3210 VPWR 0.1145
R11326 VPWR.n3207 VPWR 0.1145
R11327 VPWR.n3205 VPWR.n3204 0.1145
R11328 VPWR.n3199 VPWR 0.1145
R11329 VPWR.n3189 VPWR 0.1145
R11330 VPWR.n1152 VPWR 0.1145
R11331 VPWR.n1144 VPWR 0.1145
R11332 VPWR.n1132 VPWR 0.1145
R11333 VPWR.n1120 VPWR 0.1145
R11334 VPWR VPWR.n1843 0.1145
R11335 VPWR.n1838 VPWR 0.1145
R11336 VPWR.n664 VPWR 0.1145
R11337 VPWR.n658 VPWR 0.1145
R11338 VPWR.n1934 VPWR 0.1145
R11339 VPWR.n2001 VPWR 0.1145
R11340 VPWR VPWR.n1989 0.1145
R11341 VPWR.n1982 VPWR 0.1145
R11342 VPWR.n1971 VPWR 0.1145
R11343 VPWR.n1951 VPWR 0.1145
R11344 VPWR.n1948 VPWR 0.1145
R11345 VPWR.n2859 VPWR 0.1145
R11346 VPWR.n2898 VPWR 0.1145
R11347 VPWR.n2014 VPWR 0.1145
R11348 VPWR VPWR.n2028 0.1145
R11349 VPWR.n2025 VPWR 0.1145
R11350 VPWR.n2021 VPWR 0.1145
R11351 VPWR.n2017 VPWR 0.1145
R11352 VPWR.n2016 VPWR 0.1145
R11353 VPWR VPWR.n2714 0.1145
R11354 VPWR VPWR.n2724 0.1145
R11355 VPWR VPWR.n2727 0.1145
R11356 VPWR.n2794 VPWR 0.1145
R11357 VPWR.n2781 VPWR 0.1145
R11358 VPWR.n2063 VPWR 0.1145
R11359 VPWR.n2060 VPWR 0.1145
R11360 VPWR.n2057 VPWR 0.1145
R11361 VPWR.n2097 VPWR 0.1145
R11362 VPWR.n2078 VPWR 0.1145
R11363 VPWR VPWR.n2077 0.1145
R11364 VPWR.n2703 VPWR 0.1145
R11365 VPWR.n2698 VPWR 0.1145
R11366 VPWR.n2691 VPWR 0.1145
R11367 VPWR.n2688 VPWR 0.1145
R11368 VPWR.n2684 VPWR 0.1145
R11369 VPWR.n2654 VPWR 0.1145
R11370 VPWR VPWR.n460 0.1145
R11371 VPWR VPWR.n478 0.1145
R11372 VPWR.n479 VPWR 0.1145
R11373 VPWR VPWR.n482 0.1145
R11374 VPWR.n483 VPWR 0.1145
R11375 VPWR VPWR.n486 0.1145
R11376 VPWR.n487 VPWR 0.1145
R11377 VPWR.n500 VPWR 0.1145
R11378 VPWR VPWR.n457 0.1145
R11379 VPWR.n1851 VPWR 0.1145
R11380 VPWR VPWR.n572 0.1145
R11381 VPWR.n558 VPWR.n557 0.1145
R11382 VPWR.n556 VPWR 0.1145
R11383 VPWR VPWR.n3024 0.1145
R11384 VPWR VPWR.n3027 0.1145
R11385 VPWR VPWR.n3033 0.1145
R11386 VPWR VPWR.n362 0.1145
R11387 VPWR.n367 VPWR 0.1145
R11388 VPWR.n365 VPWR 0.1145
R11389 VPWR.n364 VPWR 0.1145
R11390 VPWR.n1916 VPWR 0.1145
R11391 VPWR.n1911 VPWR 0.1145
R11392 VPWR.n1905 VPWR 0.1145
R11393 VPWR VPWR.n1898 0.1145
R11394 VPWR VPWR.n2930 0.1145
R11395 VPWR VPWR.n2938 0.1145
R11396 VPWR VPWR.n2940 0.1145
R11397 VPWR.n3019 VPWR 0.1145
R11398 VPWR.n3000 VPWR 0.1145
R11399 VPWR VPWR.n268 0.1145
R11400 VPWR VPWR.n3703 0.1145
R11401 VPWR.n2425 VPWR 0.1145
R11402 VPWR.n2424 VPWR 0.1145
R11403 VPWR.n2419 VPWR 0.1145
R11404 VPWR.n2444 VPWR 0.1145
R11405 VPWR VPWR.n2516 0.1145
R11406 VPWR.n2589 VPWR 0.1145
R11407 VPWR.n2560 VPWR 0.1145
R11408 VPWR VPWR.n18 0.1145
R11409 VPWR.n3799 VPWR 0.1145
R11410 VPWR VPWR.n72 0.1145
R11411 VPWR.n1559 VPWR 0.11375
R11412 VPWR.n1556 VPWR 0.11375
R11413 VPWR.n1554 VPWR 0.11375
R11414 VPWR.n1550 VPWR 0.11375
R11415 VPWR VPWR.n3448 0.113
R11416 VPWR VPWR.n3463 0.113
R11417 VPWR VPWR.n3478 0.113
R11418 VPWR VPWR.n3493 0.113
R11419 VPWR VPWR.n3508 0.113
R11420 VPWR VPWR.n3523 0.113
R11421 VPWR VPWR.n3538 0.113
R11422 VPWR VPWR.n3553 0.113
R11423 VPWR VPWR.n3568 0.113
R11424 VPWR VPWR.n3583 0.113
R11425 VPWR VPWR.n3598 0.113
R11426 VPWR VPWR.n3613 0.113
R11427 VPWR VPWR.n3628 0.113
R11428 VPWR VPWR.n3643 0.113
R11429 VPWR VPWR.n3658 0.113
R11430 VPWR VPWR.n3673 0.113
R11431 VPWR.n1363 VPWR.n1362 0.113
R11432 VPWR.n1336 VPWR.n1335 0.113
R11433 VPWR.n1326 VPWR 0.113
R11434 VPWR.n1296 VPWR 0.113
R11435 VPWR.n1241 VPWR 0.113
R11436 VPWR.n769 VPWR 0.113
R11437 VPWR.n1171 VPWR.n1170 0.113
R11438 VPWR.n1182 VPWR.n1181 0.113
R11439 VPWR.n1718 VPWR.n1717 0.113
R11440 VPWR.n3176 VPWR 0.113
R11441 VPWR.n166 VPWR 0.113
R11442 VPWR.n1123 VPWR 0.113
R11443 VPWR.n649 VPWR 0.113
R11444 VPWR VPWR.n3113 0.113
R11445 VPWR VPWR.n3131 0.113
R11446 VPWR.n3154 VPWR 0.113
R11447 VPWR.n2003 VPWR 0.113
R11448 VPWR.n1975 VPWR.n1974 0.113
R11449 VPWR.n1954 VPWR 0.113
R11450 VPWR.n2889 VPWR 0.113
R11451 VPWR VPWR.n2107 0.113
R11452 VPWR VPWR.n2125 0.113
R11453 VPWR VPWR.n2139 0.113
R11454 VPWR VPWR.n2157 0.113
R11455 VPWR.n2177 VPWR 0.113
R11456 VPWR VPWR.n302 0.113
R11457 VPWR VPWR.n320 0.113
R11458 VPWR.n2269 VPWR 0.113
R11459 VPWR.n2251 VPWR 0.113
R11460 VPWR.n341 VPWR 0.113
R11461 VPWR VPWR.n2385 0.113
R11462 VPWR VPWR.n2396 0.113
R11463 VPWR VPWR.n2407 0.113
R11464 VPWR.n2309 VPWR 0.113
R11465 VPWR.n2291 VPWR 0.113
R11466 VPWR VPWR.n2191 0.113
R11467 VPWR VPWR.n2209 0.113
R11468 VPWR.n2229 VPWR 0.113
R11469 VPWR.n2052 VPWR 0.113
R11470 VPWR.n2034 VPWR 0.113
R11471 VPWR.n2710 VPWR.n194 0.113
R11472 VPWR VPWR.n2730 0.113
R11473 VPWR.n2827 VPWR 0.113
R11474 VPWR.n2809 VPWR 0.113
R11475 VPWR.n2780 VPWR 0.113
R11476 VPWR.n2760 VPWR 0.113
R11477 VPWR.n2081 VPWR 0.113
R11478 VPWR.n462 VPWR.n461 0.113
R11479 VPWR VPWR.n474 0.113
R11480 VPWR VPWR.n496 0.113
R11481 VPWR.n498 VPWR.n497 0.113
R11482 VPWR.n1862 VPWR 0.113
R11483 VPWR VPWR.n3042 0.113
R11484 VPWR.n3102 VPWR 0.113
R11485 VPWR.n3084 VPWR 0.113
R11486 VPWR.n3065 VPWR 0.113
R11487 VPWR.n1914 VPWR 0.113
R11488 VPWR.n1896 VPWR 0.113
R11489 VPWR.n3014 VPWR 0.113
R11490 VPWR.n1812 VPWR 0.11225
R11491 VPWR.n596 VPWR.n595 0.11225
R11492 VPWR VPWR.n2928 0.11225
R11493 VPWR.n1636 VPWR.n1635 0.1115
R11494 VPWR.n3700 VPWR.n3699 0.1115
R11495 VPWR VPWR.n1569 0.11075
R11496 VPWR VPWR.n2949 0.11075
R11497 VPWR.n1304 VPWR 0.11
R11498 VPWR.n2797 VPWR.n2796 0.11
R11499 VPWR.n461 VPWR 0.11
R11500 VPWR VPWR.n1894 0.11
R11501 VPWR.n1893 VPWR 0.11
R11502 VPWR VPWR.n1892 0.11
R11503 VPWR.n1887 VPWR 0.11
R11504 VPWR.n1605 VPWR 0.10925
R11505 VPWR.n1575 VPWR.n1574 0.10925
R11506 VPWR.n1373 VPWR.n1033 0.10925
R11507 VPWR.n1282 VPWR.n1281 0.10925
R11508 VPWR.n1658 VPWR.n1657 0.10925
R11509 VPWR.n1235 VPWR 0.10925
R11510 VPWR VPWR.n1733 0.10925
R11511 VPWR VPWR.n1858 0.10925
R11512 VPWR.n1520 VPWR.n1519 0.1085
R11513 VPWR.n1518 VPWR.n1517 0.1085
R11514 VPWR.n1438 VPWR.n1437 0.1085
R11515 VPWR.n1272 VPWR.n1271 0.1085
R11516 VPWR.n1334 VPWR.n1333 0.1085
R11517 VPWR.n1226 VPWR.n1225 0.1085
R11518 VPWR.n1224 VPWR.n1223 0.1085
R11519 VPWR.n1685 VPWR.n1684 0.1085
R11520 VPWR.n3235 VPWR.n3234 0.1085
R11521 VPWR.n1169 VPWR.n1168 0.1085
R11522 VPWR.n1165 VPWR.n1164 0.1085
R11523 VPWR.n1161 VPWR.n1160 0.1085
R11524 VPWR.n1213 VPWR.n1212 0.1085
R11525 VPWR.n1205 VPWR.n1204 0.1085
R11526 VPWR.n1714 VPWR.n1713 0.1085
R11527 VPWR.n1085 VPWR.n1084 0.1085
R11528 VPWR.n1130 VPWR.n1129 0.1085
R11529 VPWR.n1128 VPWR.n1127 0.1085
R11530 VPWR.n1105 VPWR.n1104 0.1085
R11531 VPWR.n688 VPWR.n687 0.1085
R11532 VPWR.n677 VPWR.n676 0.1085
R11533 VPWR.n668 VPWR.n667 0.1085
R11534 VPWR.n642 VPWR.n641 0.1085
R11535 VPWR.n1964 VPWR.n1963 0.1085
R11536 VPWR.n2719 VPWR.n2718 0.1085
R11537 VPWR.n2701 VPWR 0.1085
R11538 VPWR.n464 VPWR.n463 0.1085
R11539 VPWR.n506 VPWR.n505 0.1085
R11540 VPWR.n504 VPWR.n503 0.1085
R11541 VPWR.n1879 VPWR.n1878 0.1085
R11542 VPWR.n1873 VPWR.n1872 0.1085
R11543 VPWR.n1869 VPWR.n1868 0.1085
R11544 VPWR.n451 VPWR.n450 0.1085
R11545 VPWR.n449 VPWR.n448 0.1085
R11546 VPWR.n2940 VPWR.n2939 0.1085
R11547 VPWR VPWR.n119 0.107
R11548 VPWR VPWR.n3351 0.107
R11549 VPWR VPWR.n807 0.107
R11550 VPWR VPWR.n800 0.107
R11551 VPWR VPWR.n1190 0.107
R11552 VPWR VPWR.n1134 0.107
R11553 VPWR VPWR.n1103 0.107
R11554 VPWR VPWR.n1667 0.10625
R11555 VPWR.n692 VPWR 0.10625
R11556 VPWR.n560 VPWR 0.10625
R11557 VPWR VPWR.n398 0.10625
R11558 VPWR.n1361 VPWR.n1360 0.1055
R11559 VPWR.n1612 VPWR.n1611 0.1055
R11560 VPWR.n3377 VPWR.n3376 0.1055
R11561 VPWR.n3286 VPWR.n3285 0.1055
R11562 VPWR.n1791 VPWR.n1790 0.1055
R11563 VPWR.n3214 VPWR.n3213 0.1055
R11564 VPWR.n3191 VPWR.n3190 0.1055
R11565 VPWR VPWR.n2834 0.1055
R11566 VPWR.n2895 VPWR.n2894 0.1055
R11567 VPWR.n1865 VPWR 0.1055
R11568 VPWR VPWR.n560 0.1055
R11569 VPWR.n551 VPWR.n550 0.1055
R11570 VPWR.n3029 VPWR.n3028 0.1055
R11571 VPWR VPWR.n1106 0.10475
R11572 VPWR VPWR.n1374 0.104
R11573 VPWR.n1452 VPWR 0.104
R11574 VPWR VPWR.n1609 0.104
R11575 VPWR.n1196 VPWR.n1195 0.104
R11576 VPWR.n1348 VPWR 0.1025
R11577 VPWR.n1290 VPWR 0.1025
R11578 VPWR VPWR.n889 0.1025
R11579 VPWR.n1736 VPWR 0.1025
R11580 VPWR VPWR.n1757 0.1025
R11581 VPWR VPWR.n1991 0.1025
R11582 VPWR VPWR.n2079 0.1025
R11583 VPWR.n1864 VPWR.n1863 0.1025
R11584 VPWR.n3023 VPWR 0.1025
R11585 VPWR VPWR.n2924 0.1025
R11586 VPWR.n1310 VPWR 0.10175
R11587 VPWR VPWR.n1656 0.10175
R11588 VPWR.n1135 VPWR 0.10175
R11589 VPWR.n3401 VPWR.n3400 0.101
R11590 VPWR VPWR.n1760 0.101
R11591 VPWR.n3756 VPWR.n60 0.101
R11592 VPWR.n3753 VPWR.n3752 0.101
R11593 VPWR VPWR.n1303 0.10025
R11594 VPWR VPWR.n1136 0.10025
R11595 VPWR VPWR.n509 0.10025
R11596 VPWR.n1486 VPWR 0.0995
R11597 VPWR VPWR.n910 0.0995
R11598 VPWR VPWR.n1593 0.0995
R11599 VPWR.n1592 VPWR 0.0995
R11600 VPWR.n1586 VPWR 0.0995
R11601 VPWR.n1583 VPWR 0.0995
R11602 VPWR VPWR.n1532 0.0995
R11603 VPWR.n1569 VPWR 0.0995
R11604 VPWR.n1566 VPWR 0.0995
R11605 VPWR.n1563 VPWR 0.0995
R11606 VPWR.n1462 VPWR 0.0995
R11607 VPWR.n1632 VPWR.n1631 0.0995
R11608 VPWR.n1630 VPWR.n1629 0.0995
R11609 VPWR VPWR.n1288 0.0995
R11610 VPWR VPWR.n1286 0.0995
R11611 VPWR.n810 VPWR.n809 0.0995
R11612 VPWR.n3305 VPWR.n3304 0.0995
R11613 VPWR.n1802 VPWR.n1801 0.0995
R11614 VPWR.n1108 VPWR 0.0995
R11615 VPWR VPWR.n2914 0.0995
R11616 VPWR.n2642 VPWR 0.0995
R11617 VPWR.n968 VPWR 0.09875
R11618 VPWR.n802 VPWR.n801 0.09875
R11619 VPWR VPWR.n3253 0.09875
R11620 VPWR.n1754 VPWR 0.09875
R11621 VPWR VPWR.n596 0.09875
R11622 VPWR.n566 VPWR.n565 0.09875
R11623 VPWR.n1643 VPWR.n1642 0.098
R11624 VPWR.n788 VPWR 0.098
R11625 VPWR VPWR.n3202 0.098
R11626 VPWR.n2646 VPWR.n2645 0.098
R11627 VPWR VPWR.n3237 0.09725
R11628 VPWR VPWR.n1719 0.09725
R11629 VPWR.n1843 VPWR 0.09725
R11630 VPWR.n572 VPWR 0.09725
R11631 VPWR.n1349 VPWR.n1348 0.0965
R11632 VPWR VPWR.n1450 0.0965
R11633 VPWR VPWR.n1015 0.0965
R11634 VPWR.n994 VPWR.n993 0.0965
R11635 VPWR VPWR.n1329 0.0965
R11636 VPWR VPWR.n1315 0.0965
R11637 VPWR.n1666 VPWR.n1665 0.0965
R11638 VPWR.n3330 VPWR 0.0965
R11639 VPWR VPWR.n1233 0.0965
R11640 VPWR VPWR.n3276 0.0965
R11641 VPWR.n1186 VPWR 0.0965
R11642 VPWR.n1757 VPWR.n1756 0.0965
R11643 VPWR.n1101 VPWR 0.0965
R11644 VPWR VPWR.n660 0.0965
R11645 VPWR.n2854 VPWR.n2853 0.0965
R11646 VPWR VPWR.n403 0.0965
R11647 VPWR VPWR.n2948 0.0965
R11648 VPWR VPWR.n3449 0.09575
R11649 VPWR VPWR.n3464 0.09575
R11650 VPWR VPWR.n3479 0.09575
R11651 VPWR VPWR.n3494 0.09575
R11652 VPWR VPWR.n3509 0.09575
R11653 VPWR VPWR.n3524 0.09575
R11654 VPWR VPWR.n3539 0.09575
R11655 VPWR VPWR.n3554 0.09575
R11656 VPWR VPWR.n3569 0.09575
R11657 VPWR VPWR.n3584 0.09575
R11658 VPWR VPWR.n3599 0.09575
R11659 VPWR VPWR.n3614 0.09575
R11660 VPWR VPWR.n3629 0.09575
R11661 VPWR VPWR.n3644 0.09575
R11662 VPWR VPWR.n3659 0.09575
R11663 VPWR VPWR.n3674 0.09575
R11664 VPWR VPWR.n1600 0.09575
R11665 VPWR VPWR.n1585 0.09575
R11666 VPWR VPWR.n1581 0.09575
R11667 VPWR VPWR.n1568 0.09575
R11668 VPWR VPWR.n1565 0.09575
R11669 VPWR VPWR.n1558 0.09575
R11670 VPWR VPWR.n1555 0.09575
R11671 VPWR VPWR.n1549 0.09575
R11672 VPWR.n1354 VPWR 0.09575
R11673 VPWR VPWR.n1467 0.09575
R11674 VPWR VPWR.n1464 0.09575
R11675 VPWR VPWR.n1438 0.09575
R11676 VPWR VPWR.n1314 0.09575
R11677 VPWR VPWR.n1313 0.09575
R11678 VPWR.n3335 VPWR 0.09575
R11679 VPWR VPWR.n3368 0.09575
R11680 VPWR VPWR.n3363 0.09575
R11681 VPWR VPWR.n768 0.09575
R11682 VPWR.n3238 VPWR 0.09575
R11683 VPWR VPWR.n3298 0.09575
R11684 VPWR VPWR.n3293 0.09575
R11685 VPWR VPWR.n3284 0.09575
R11686 VPWR.n1770 VPWR 0.09575
R11687 VPWR VPWR.n1797 0.09575
R11688 VPWR VPWR.n3217 0.09575
R11689 VPWR VPWR.n2001 0.09575
R11690 VPWR VPWR.n1976 0.09575
R11691 VPWR.n2846 VPWR 0.09575
R11692 VPWR VPWR.n2898 0.09575
R11693 VPWR VPWR.n2888 0.09575
R11694 VPWR.n2135 VPWR 0.09575
R11695 VPWR VPWR.n2388 0.09575
R11696 VPWR VPWR.n2399 0.09575
R11697 VPWR VPWR.n2410 0.09575
R11698 VPWR VPWR.n2322 0.09575
R11699 VPWR VPWR.n2018 0.09575
R11700 VPWR.n2727 VPWR 0.09575
R11701 VPWR VPWR.n2064 0.09575
R11702 VPWR VPWR.n2083 0.09575
R11703 VPWR VPWR.n2692 0.09575
R11704 VPWR.n459 VPWR 0.09575
R11705 VPWR VPWR.n1869 0.09575
R11706 VPWR VPWR.n1851 0.09575
R11707 VPWR VPWR.n570 0.09575
R11708 VPWR.n2930 VPWR 0.09575
R11709 VPWR VPWR.n3016 0.09575
R11710 VPWR.n268 VPWR 0.09575
R11711 VPWR.n3701 VPWR 0.09575
R11712 VPWR VPWR.n2426 0.09575
R11713 VPWR.n472 VPWR.n471 0.095
R11714 VPWR VPWR.n2942 0.095
R11715 VPWR.n1382 VPWR.n1381 0.09425
R11716 VPWR.n3434 VPWR 0.09425
R11717 VPWR.n216 VPWR 0.09425
R11718 VPWR.n1860 VPWR.n1859 0.09425
R11719 VPWR.n3720 VPWR 0.09425
R11720 VPWR VPWR.n1361 0.0935
R11721 VPWR.n1611 VPWR 0.0935
R11722 VPWR.n1312 VPWR 0.0935
R11723 VPWR.n3239 VPWR 0.0935
R11724 VPWR.n3308 VPWR 0.0935
R11725 VPWR VPWR.n1740 0.0935
R11726 VPWR.n414 VPWR.n413 0.0935
R11727 VPWR VPWR.n3248 0.09275
R11728 VPWR.n516 VPWR.t5174 0.0922506
R11729 VPWR.n1053 VPWR.n1052 0.092
R11730 VPWR VPWR.n983 0.092
R11731 VPWR.n1260 VPWR 0.092
R11732 VPWR VPWR.n2929 0.092
R11733 VPWR.n681 VPWR.n680 0.09125
R11734 VPWR.n1344 VPWR.n1343 0.0905
R11735 VPWR.n1742 VPWR.n1741 0.0905
R11736 VPWR VPWR.n666 0.0905
R11737 VPWR.n2004 VPWR.n2003 0.0905
R11738 VPWR.n2053 VPWR.n2052 0.0905
R11739 VPWR.n2098 VPWR.n2097 0.0905
R11740 VPWR.n588 VPWR.n587 0.0905
R11741 VPWR.n2454 VPWR.n2453 0.0905
R11742 VPWR.n1376 VPWR.n1375 0.08975
R11743 VPWR.n2451 VPWR 0.08975
R11744 VPWR.n1353 VPWR.n1352 0.089
R11745 VPWR VPWR.n997 0.089
R11746 VPWR.n1305 VPWR.n1304 0.089
R11747 VPWR.n1247 VPWR.n1246 0.089
R11748 VPWR.n806 VPWR.n805 0.089
R11749 VPWR.n804 VPWR.n803 0.089
R11750 VPWR.n1978 VPWR.n1977 0.089
R11751 VPWR.n2694 VPWR.n2693 0.089
R11752 VPWR.n491 VPWR.n490 0.089
R11753 VPWR.n1919 VPWR.n1918 0.089
R11754 VPWR.n1908 VPWR.n1907 0.089
R11755 VPWR.n1892 VPWR.n1891 0.089
R11756 VPWR.n1888 VPWR.n1887 0.089
R11757 VPWR.n1886 VPWR.n1885 0.089
R11758 VPWR.n430 VPWR 0.089
R11759 VPWR.n1488 VPWR.n1487 0.0875
R11760 VPWR.n1193 VPWR.n1192 0.0875
R11761 VPWR.n998 VPWR 0.08675
R11762 VPWR VPWR.n1651 0.08675
R11763 VPWR VPWR.n862 0.08675
R11764 VPWR.n801 VPWR 0.08675
R11765 VPWR VPWR.n3240 0.08675
R11766 VPWR VPWR.n1853 0.08675
R11767 VPWR.n1470 VPWR 0.086
R11768 VPWR.n1638 VPWR 0.086
R11769 VPWR.n1320 VPWR.n1319 0.08525
R11770 VPWR.n1803 VPWR 0.08525
R11771 VPWR.n404 VPWR 0.08525
R11772 VPWR.n1045 VPWR.n1044 0.0845
R11773 VPWR.n1047 VPWR.n1046 0.0845
R11774 VPWR.n1049 VPWR.n1048 0.0845
R11775 VPWR.n1051 VPWR.n1050 0.0845
R11776 VPWR.n1358 VPWR.n1357 0.0845
R11777 VPWR.n1384 VPWR 0.0845
R11778 VPWR.n1459 VPWR.n1458 0.0845
R11779 VPWR.n1458 VPWR.n1457 0.0845
R11780 VPWR.n1454 VPWR.n1453 0.0845
R11781 VPWR.n981 VPWR 0.0845
R11782 VPWR.n980 VPWR.n979 0.0845
R11783 VPWR.n971 VPWR 0.0845
R11784 VPWR VPWR.n3416 0.0845
R11785 VPWR.n1269 VPWR.n1268 0.0845
R11786 VPWR.n1267 VPWR.n1266 0.0845
R11787 VPWR.n1324 VPWR.n1323 0.0845
R11788 VPWR.n1307 VPWR.n1306 0.0845
R11789 VPWR.n1259 VPWR.n1258 0.0845
R11790 VPWR.n1257 VPWR.n1256 0.0845
R11791 VPWR.n1255 VPWR.n1254 0.0845
R11792 VPWR.n1253 VPWR.n1252 0.0845
R11793 VPWR.n1251 VPWR.n1250 0.0845
R11794 VPWR.n1249 VPWR.n1248 0.0845
R11795 VPWR.n1243 VPWR.n1242 0.0845
R11796 VPWR.n1692 VPWR.n1691 0.0845
R11797 VPWR.n1689 VPWR.n1688 0.0845
R11798 VPWR.n1191 VPWR 0.0845
R11799 VPWR.n1810 VPWR.n1809 0.0845
R11800 VPWR.n3180 VPWR.n3179 0.0845
R11801 VPWR.n3172 VPWR.n3171 0.0845
R11802 VPWR.n3170 VPWR.n3169 0.0845
R11803 VPWR.n3168 VPWR.n3167 0.0845
R11804 VPWR.n3166 VPWR.n3165 0.0845
R11805 VPWR.n3164 VPWR.n3163 0.0845
R11806 VPWR.n168 VPWR.n167 0.0845
R11807 VPWR.n1155 VPWR.n1154 0.0845
R11808 VPWR.n1121 VPWR.n1120 0.0845
R11809 VPWR.n1119 VPWR.n1118 0.0845
R11810 VPWR.n1114 VPWR.n1113 0.0845
R11811 VPWR.n659 VPWR.n658 0.0845
R11812 VPWR.n657 VPWR.n656 0.0845
R11813 VPWR.n655 VPWR.n654 0.0845
R11814 VPWR.n651 VPWR.n650 0.0845
R11815 VPWR.n641 VPWR.n640 0.0845
R11816 VPWR.n639 VPWR.n638 0.0845
R11817 VPWR.n637 VPWR.n636 0.0845
R11818 VPWR.n3112 VPWR.n3111 0.0845
R11819 VPWR.n3116 VPWR.n3115 0.0845
R11820 VPWR.n3118 VPWR.n3117 0.0845
R11821 VPWR.n3120 VPWR.n3119 0.0845
R11822 VPWR.n3122 VPWR.n3121 0.0845
R11823 VPWR.n3126 VPWR.n3125 0.0845
R11824 VPWR.n3128 VPWR.n3127 0.0845
R11825 VPWR.n3130 VPWR.n3129 0.0845
R11826 VPWR.n3141 VPWR.n3140 0.0845
R11827 VPWR.n3139 VPWR.n3138 0.0845
R11828 VPWR.n3137 VPWR.n3136 0.0845
R11829 VPWR.n3135 VPWR.n3134 0.0845
R11830 VPWR.n3133 VPWR.n3132 0.0845
R11831 VPWR.n3156 VPWR.n3155 0.0845
R11832 VPWR.n1935 VPWR.n1934 0.0845
R11833 VPWR.n1933 VPWR.n1932 0.0845
R11834 VPWR.n1931 VPWR.n1930 0.0845
R11835 VPWR.n1927 VPWR.n1926 0.0845
R11836 VPWR.n1991 VPWR.n1990 0.0845
R11837 VPWR.n1989 VPWR.n1988 0.0845
R11838 VPWR.n1983 VPWR.n1982 0.0845
R11839 VPWR.n1981 VPWR.n1980 0.0845
R11840 VPWR.n1958 VPWR.n1957 0.0845
R11841 VPWR.n1952 VPWR.n1951 0.0845
R11842 VPWR.n2840 VPWR.n2839 0.0845
R11843 VPWR.n2842 VPWR.n2841 0.0845
R11844 VPWR.n351 VPWR.n350 0.0845
R11845 VPWR.n353 VPWR.n352 0.0845
R11846 VPWR.n355 VPWR.n354 0.0845
R11847 VPWR.n2104 VPWR.n2103 0.0845
R11848 VPWR.n2106 VPWR.n2105 0.0845
R11849 VPWR.n2112 VPWR.n2111 0.0845
R11850 VPWR.n2114 VPWR.n2113 0.0845
R11851 VPWR.n2116 VPWR.n2115 0.0845
R11852 VPWR.n2118 VPWR.n2117 0.0845
R11853 VPWR.n2120 VPWR.n2119 0.0845
R11854 VPWR.n2122 VPWR.n2121 0.0845
R11855 VPWR.n2124 VPWR.n2123 0.0845
R11856 VPWR.n2136 VPWR.n2135 0.0845
R11857 VPWR.n2138 VPWR.n2137 0.0845
R11858 VPWR.n2142 VPWR.n2141 0.0845
R11859 VPWR.n2144 VPWR.n2143 0.0845
R11860 VPWR.n2146 VPWR.n2145 0.0845
R11861 VPWR.n2148 VPWR.n2147 0.0845
R11862 VPWR.n2152 VPWR.n2151 0.0845
R11863 VPWR.n2154 VPWR.n2153 0.0845
R11864 VPWR.n2156 VPWR.n2155 0.0845
R11865 VPWR.n2164 VPWR.n2163 0.0845
R11866 VPWR.n2162 VPWR.n2161 0.0845
R11867 VPWR.n2160 VPWR.n2159 0.0845
R11868 VPWR.n2158 VPWR.n348 0.0845
R11869 VPWR.n2183 VPWR.n2182 0.0845
R11870 VPWR.n2181 VPWR.n2180 0.0845
R11871 VPWR.n2179 VPWR.n2178 0.0845
R11872 VPWR.n288 VPWR.n287 0.0845
R11873 VPWR.n290 VPWR.n289 0.0845
R11874 VPWR.n292 VPWR.n291 0.0845
R11875 VPWR.n299 VPWR.n298 0.0845
R11876 VPWR.n301 VPWR.n300 0.0845
R11877 VPWR.n307 VPWR.n306 0.0845
R11878 VPWR.n309 VPWR.n308 0.0845
R11879 VPWR.n311 VPWR.n310 0.0845
R11880 VPWR.n313 VPWR.n312 0.0845
R11881 VPWR.n315 VPWR.n314 0.0845
R11882 VPWR.n317 VPWR.n316 0.0845
R11883 VPWR.n319 VPWR.n318 0.0845
R11884 VPWR.n328 VPWR.n327 0.0845
R11885 VPWR.n326 VPWR.n325 0.0845
R11886 VPWR.n324 VPWR.n323 0.0845
R11887 VPWR.n322 VPWR.n321 0.0845
R11888 VPWR.n2273 VPWR.n2272 0.0845
R11889 VPWR.n2271 VPWR.n2270 0.0845
R11890 VPWR.n2265 VPWR.n2264 0.0845
R11891 VPWR.n2263 VPWR.n2262 0.0845
R11892 VPWR.n2261 VPWR.n2260 0.0845
R11893 VPWR.n2259 VPWR.n2258 0.0845
R11894 VPWR.n2257 VPWR.n2256 0.0845
R11895 VPWR.n2255 VPWR.n2254 0.0845
R11896 VPWR.n2253 VPWR.n2252 0.0845
R11897 VPWR.n2247 VPWR.n2246 0.0845
R11898 VPWR.n2245 VPWR.n2244 0.0845
R11899 VPWR.n2243 VPWR.n2242 0.0845
R11900 VPWR.n2241 VPWR.n2240 0.0845
R11901 VPWR.n347 VPWR.n346 0.0845
R11902 VPWR.n345 VPWR.n344 0.0845
R11903 VPWR.n343 VPWR.n342 0.0845
R11904 VPWR.n282 VPWR.n281 0.0845
R11905 VPWR.n280 VPWR.n279 0.0845
R11906 VPWR.n278 VPWR.n277 0.0845
R11907 VPWR.n2313 VPWR.n2312 0.0845
R11908 VPWR.n2311 VPWR.n2310 0.0845
R11909 VPWR.n2305 VPWR.n2304 0.0845
R11910 VPWR.n2303 VPWR.n2302 0.0845
R11911 VPWR.n2301 VPWR.n2300 0.0845
R11912 VPWR.n2299 VPWR.n2298 0.0845
R11913 VPWR.n2297 VPWR.n2296 0.0845
R11914 VPWR.n2295 VPWR.n2294 0.0845
R11915 VPWR.n2293 VPWR.n2292 0.0845
R11916 VPWR.n2287 VPWR.n2286 0.0845
R11917 VPWR.n2285 VPWR.n2284 0.0845
R11918 VPWR.n2283 VPWR.n2282 0.0845
R11919 VPWR.n2281 VPWR.n2280 0.0845
R11920 VPWR.n2188 VPWR.n2187 0.0845
R11921 VPWR.n2190 VPWR.n2189 0.0845
R11922 VPWR.n2196 VPWR.n2195 0.0845
R11923 VPWR.n2198 VPWR.n2197 0.0845
R11924 VPWR.n2200 VPWR.n2199 0.0845
R11925 VPWR.n2202 VPWR.n2201 0.0845
R11926 VPWR.n2204 VPWR.n2203 0.0845
R11927 VPWR.n2206 VPWR.n2205 0.0845
R11928 VPWR.n2208 VPWR.n2207 0.0845
R11929 VPWR.n2216 VPWR.n2215 0.0845
R11930 VPWR.n2214 VPWR.n2213 0.0845
R11931 VPWR.n2212 VPWR.n2211 0.0845
R11932 VPWR.n2210 VPWR.n2186 0.0845
R11933 VPWR.n2235 VPWR.n2234 0.0845
R11934 VPWR.n2233 VPWR.n2232 0.0845
R11935 VPWR.n2231 VPWR.n2230 0.0845
R11936 VPWR.n2015 VPWR.n2014 0.0845
R11937 VPWR.n2013 VPWR.n2012 0.0845
R11938 VPWR.n2011 VPWR.n2010 0.0845
R11939 VPWR.n2007 VPWR.n2006 0.0845
R11940 VPWR.n2050 VPWR.n2049 0.0845
R11941 VPWR.n2048 VPWR.n2047 0.0845
R11942 VPWR.n2046 VPWR.n2045 0.0845
R11943 VPWR.n2044 VPWR.n2043 0.0845
R11944 VPWR.n2040 VPWR.n2039 0.0845
R11945 VPWR.n2038 VPWR.n2037 0.0845
R11946 VPWR.n2036 VPWR.n2035 0.0845
R11947 VPWR.n2032 VPWR.n2031 0.0845
R11948 VPWR.n2030 VPWR.n2029 0.0845
R11949 VPWR.n2028 VPWR.n2027 0.0845
R11950 VPWR.n2026 VPWR.n2025 0.0845
R11951 VPWR.n2024 VPWR.n2023 0.0845
R11952 VPWR.n2022 VPWR.n2021 0.0845
R11953 VPWR.n2020 VPWR.n2019 0.0845
R11954 VPWR.n2714 VPWR.n2713 0.0845
R11955 VPWR.n2724 VPWR.n2723 0.0845
R11956 VPWR.n2726 VPWR.n2725 0.0845
R11957 VPWR.n2745 VPWR.n2744 0.0845
R11958 VPWR.n2743 VPWR.n2742 0.0845
R11959 VPWR.n2741 VPWR.n2740 0.0845
R11960 VPWR.n2739 VPWR.n2738 0.0845
R11961 VPWR.n2735 VPWR.n2734 0.0845
R11962 VPWR.n2733 VPWR.n2732 0.0845
R11963 VPWR.n2731 VPWR.n192 0.0845
R11964 VPWR.n2823 VPWR.n2822 0.0845
R11965 VPWR.n2821 VPWR.n2820 0.0845
R11966 VPWR.n2819 VPWR.n2818 0.0845
R11967 VPWR.n2817 VPWR.n2816 0.0845
R11968 VPWR.n2815 VPWR.n2814 0.0845
R11969 VPWR.n2813 VPWR.n2812 0.0845
R11970 VPWR.n2811 VPWR.n2810 0.0845
R11971 VPWR.n2784 VPWR.n2783 0.0845
R11972 VPWR.n2782 VPWR.n2781 0.0845
R11973 VPWR.n2776 VPWR.n2775 0.0845
R11974 VPWR.n2774 VPWR.n2773 0.0845
R11975 VPWR.n2772 VPWR.n2771 0.0845
R11976 VPWR.n2770 VPWR.n2769 0.0845
R11977 VPWR.n2768 VPWR.n2767 0.0845
R11978 VPWR.n2766 VPWR.n2765 0.0845
R11979 VPWR.n2083 VPWR.n2082 0.0845
R11980 VPWR.n2704 VPWR.n2703 0.0845
R11981 VPWR.n2702 VPWR.n2701 0.0845
R11982 VPWR.n2699 VPWR.n2698 0.0845
R11983 VPWR.n2696 VPWR.n2695 0.0845
R11984 VPWR.n234 VPWR 0.0845
R11985 VPWR VPWR.n475 0.0845
R11986 VPWR.n510 VPWR 0.0845
R11987 VPWR.n598 VPWR 0.0845
R11988 VPWR.n594 VPWR 0.0845
R11989 VPWR.n3033 VPWR.n3032 0.0845
R11990 VPWR.n3035 VPWR.n3034 0.0845
R11991 VPWR.n3037 VPWR.n3036 0.0845
R11992 VPWR.n3041 VPWR.n3040 0.0845
R11993 VPWR.n3052 VPWR.n3051 0.0845
R11994 VPWR.n3050 VPWR.n3049 0.0845
R11995 VPWR.n3048 VPWR.n3047 0.0845
R11996 VPWR.n3046 VPWR.n3045 0.0845
R11997 VPWR.n3044 VPWR.n3043 0.0845
R11998 VPWR.n3104 VPWR.n3103 0.0845
R11999 VPWR.n3098 VPWR.n3097 0.0845
R12000 VPWR.n3096 VPWR.n3095 0.0845
R12001 VPWR.n3094 VPWR.n3093 0.0845
R12002 VPWR.n3092 VPWR.n3091 0.0845
R12003 VPWR.n3090 VPWR.n3089 0.0845
R12004 VPWR.n3088 VPWR.n3087 0.0845
R12005 VPWR.n3086 VPWR.n3085 0.0845
R12006 VPWR.n3080 VPWR.n3079 0.0845
R12007 VPWR.n3078 VPWR.n3077 0.0845
R12008 VPWR.n3076 VPWR.n3075 0.0845
R12009 VPWR.n3074 VPWR.n3073 0.0845
R12010 VPWR.n3072 VPWR.n3071 0.0845
R12011 VPWR.n3067 VPWR.n3066 0.0845
R12012 VPWR.n1921 VPWR.n1920 0.0845
R12013 VPWR.n1917 VPWR.n1916 0.0845
R12014 VPWR.n1912 VPWR.n1911 0.0845
R12015 VPWR.n1910 VPWR.n1909 0.0845
R12016 VPWR.n1906 VPWR.n1905 0.0845
R12017 VPWR.n1904 VPWR.n1903 0.0845
R12018 VPWR.n1900 VPWR.n1899 0.0845
R12019 VPWR.n1898 VPWR.n1897 0.0845
R12020 VPWR.n1895 VPWR 0.0845
R12021 VPWR.n442 VPWR.n441 0.0845
R12022 VPWR.n440 VPWR.n439 0.0845
R12023 VPWR.n2937 VPWR.n2936 0.0845
R12024 VPWR.n3012 VPWR.n3011 0.0845
R12025 VPWR.n3010 VPWR.n3009 0.0845
R12026 VPWR.n3006 VPWR.n3005 0.0845
R12027 VPWR.n3004 VPWR.n3003 0.0845
R12028 VPWR.n3002 VPWR.n3001 0.0845
R12029 VPWR.n3737 VPWR 0.0845
R12030 VPWR.n1633 VPWR 0.083
R12031 VPWR VPWR.n1312 0.083
R12032 VPWR VPWR.n3370 0.083
R12033 VPWR.n3109 VPWR.n172 0.083
R12034 VPWR.n2132 VPWR 0.083
R12035 VPWR VPWR.n2319 0.083
R12036 VPWR.n3106 VPWR.n173 0.083
R12037 VPWR.n2991 VPWR.n2990 0.083
R12038 VPWR.n1806 VPWR.n1805 0.08225
R12039 VPWR VPWR.n1671 0.0815
R12040 VPWR VPWR.n1700 0.0815
R12041 VPWR.n1776 VPWR.n1775 0.0815
R12042 VPWR.n673 VPWR.n672 0.0815
R12043 VPWR.n1849 VPWR 0.0815
R12044 VPWR VPWR.n104 0.08
R12045 VPWR.n1048 VPWR.n1047 0.08
R12046 VPWR.n3375 VPWR 0.08
R12047 VPWR.n1250 VPWR.n1249 0.08
R12048 VPWR.n1721 VPWR.n1720 0.08
R12049 VPWR VPWR.n1743 0.08
R12050 VPWR.n1124 VPWR.n1123 0.08
R12051 VPWR.n1980 VPWR.n1979 0.08
R12052 VPWR.n2023 VPWR.n2022 0.08
R12053 VPWR.n2076 VPWR.n2075 0.08
R12054 VPWR.n2697 VPWR.n2696 0.08
R12055 VPWR.n489 VPWR.n488 0.08
R12056 VPWR.n1922 VPWR.n1921 0.08
R12057 VPWR.n1915 VPWR.n1914 0.08
R12058 VPWR.n593 VPWR.n592 0.07925
R12059 VPWR.n1079 VPWR.n1054 0.0785
R12060 VPWR.n1004 VPWR.n1003 0.0785
R12061 VPWR.n3208 VPWR 0.0785
R12062 VPWR.n2101 VPWR.n358 0.0785
R12063 VPWR.n296 VPWR.n295 0.0785
R12064 VPWR.n2315 VPWR.n274 0.0785
R12065 VPWR.n2098 VPWR.n2055 0.0785
R12066 VPWR.n2454 VPWR.n2417 0.0785
R12067 VPWR.n1383 VPWR 0.07775
R12068 VPWR.n967 VPWR 0.077
R12069 VPWR.n3349 VPWR.n3348 0.077
R12070 VPWR.n3370 VPWR 0.077
R12071 VPWR.n1194 VPWR.n1193 0.077
R12072 VPWR.n2904 VPWR 0.077
R12073 VPWR.n571 VPWR 0.077
R12074 VPWR VPWR.n3025 0.077
R12075 VPWR VPWR.n1378 0.0755
R12076 VPWR.n3353 VPWR.n3352 0.0755
R12077 VPWR VPWR.n3206 0.0755
R12078 VPWR.n3018 VPWR.n3017 0.0755
R12079 VPWR VPWR.n1440 0.07475
R12080 VPWR.n1671 VPWR.n1670 0.07475
R12081 VPWR VPWR.n1738 0.074
R12082 VPWR.n1157 VPWR.n1080 0.074
R12083 VPWR.n1827 VPWR.n1826 0.074
R12084 VPWR.n982 VPWR 0.07325
R12085 VPWR.n1314 VPWR 0.07325
R12086 VPWR VPWR.n1721 0.07325
R12087 VPWR.n1153 VPWR 0.07325
R12088 VPWR.n1133 VPWR 0.07325
R12089 VPWR.n1052 VPWR.n1051 0.0725
R12090 VPWR.n1467 VPWR 0.0725
R12091 VPWR VPWR.n986 0.0725
R12092 VPWR VPWR.n3377 0.0725
R12093 VPWR.n1291 VPWR 0.0725
R12094 VPWR VPWR.n897 0.0725
R12095 VPWR.n882 VPWR.n881 0.0725
R12096 VPWR.n3331 VPWR 0.0725
R12097 VPWR VPWR.n1678 0.0725
R12098 VPWR VPWR.n1677 0.0725
R12099 VPWR.n3234 VPWR 0.0725
R12100 VPWR.n1738 VPWR.n1737 0.0725
R12101 VPWR.n1759 VPWR.n1758 0.0725
R12102 VPWR VPWR.n1800 0.0725
R12103 VPWR.n1104 VPWR 0.0725
R12104 VPWR.n1836 VPWR 0.0725
R12105 VPWR.n644 VPWR 0.0725
R12106 VPWR.n1945 VPWR 0.0725
R12107 VPWR VPWR.n549 0.0725
R12108 VPWR.n436 VPWR 0.0725
R12109 VPWR.n422 VPWR 0.0725
R12110 VPWR VPWR.n418 0.0725
R12111 VPWR VPWR.n1459 0.07175
R12112 VPWR.n1432 VPWR.n1431 0.07175
R12113 VPWR VPWR.n787 0.07175
R12114 VPWR VPWR.n1959 0.07175
R12115 VPWR.n473 VPWR 0.07175
R12116 VPWR VPWR.n559 0.07175
R12117 VPWR.n1311 VPWR.n1310 0.071
R12118 VPWR.n900 VPWR.n899 0.071
R12119 VPWR.n2947 VPWR 0.071
R12120 VPWR.n2575 VPWR.n2574 0.071
R12121 VPWR.n1294 VPWR.n1293 0.0695
R12122 VPWR.n3251 VPWR.n3250 0.0695
R12123 VPWR.n691 VPWR 0.0695
R12124 VPWR.n553 VPWR.n552 0.0695
R12125 VPWR.n1266 VPWR 0.06875
R12126 VPWR.n2019 VPWR 0.06875
R12127 VPWR VPWR.n2726 0.06875
R12128 VPWR.n1561 VPWR.n1560 0.068
R12129 VPWR.n3400 VPWR.n3399 0.068
R12130 VPWR.n3753 VPWR.n62 0.068
R12131 VPWR.n1040 VPWR 0.06725
R12132 VPWR.n1375 VPWR 0.06725
R12133 VPWR.n858 VPWR 0.06725
R12134 VPWR.n805 VPWR 0.06725
R12135 VPWR VPWR.n804 0.06725
R12136 VPWR.n1808 VPWR.n1807 0.06725
R12137 VPWR.n3372 VPWR.n107 0.0665
R12138 VPWR.n1680 VPWR.n1679 0.0665
R12139 VPWR VPWR.n1731 0.0665
R12140 VPWR.n1157 VPWR.n1156 0.0665
R12141 VPWR.n2836 VPWR.n2835 0.0665
R12142 VPWR.n2907 VPWR.n2906 0.0665
R12143 VPWR.n2788 VPWR.n2787 0.0665
R12144 VPWR.n1628 VPWR 0.06575
R12145 VPWR.n1653 VPWR.n1652 0.06575
R12146 VPWR.n3201 VPWR.n3200 0.06575
R12147 VPWR.n1629 VPWR.n1628 0.065
R12148 VPWR.n3233 VPWR.n3232 0.065
R12149 VPWR.n1852 VPWR 0.06425
R12150 VPWR.n1378 VPWR.n1377 0.0635
R12151 VPWR.n1450 VPWR.n1449 0.0635
R12152 VPWR VPWR.n871 0.0635
R12153 VPWR.n3297 VPWR.n3296 0.0635
R12154 VPWR.n1773 VPWR.n1772 0.0635
R12155 VPWR.n1796 VPWR 0.0635
R12156 VPWR VPWR.n3211 0.0635
R12157 VPWR.n670 VPWR 0.0635
R12158 VPWR.n663 VPWR.n662 0.0635
R12159 VPWR.n2828 VPWR.n192 0.0635
R12160 VPWR.n587 VPWR.n586 0.0635
R12161 VPWR.n546 VPWR 0.0635
R12162 VPWR VPWR.n428 0.0635
R12163 VPWR.n421 VPWR.n420 0.0635
R12164 VPWR VPWR.n1006 0.06275
R12165 VPWR.n1380 VPWR.n1379 0.062
R12166 VPWR.n1006 VPWR 0.062
R12167 VPWR.n1264 VPWR.n1263 0.062
R12168 VPWR.n3313 VPWR 0.062
R12169 VPWR.n3195 VPWR.n3194 0.062
R12170 VPWR.n1959 VPWR 0.062
R12171 VPWR.n2068 VPWR 0.062
R12172 VPWR.n559 VPWR 0.062
R12173 VPWR.n557 VPWR 0.062
R12174 VPWR.n1355 VPWR.n1354 0.0605
R12175 VPWR VPWR.n879 0.0605
R12176 VPWR.n860 VPWR 0.0605
R12177 VPWR.n1225 VPWR.n1224 0.0605
R12178 VPWR.n1204 VPWR.n1203 0.0605
R12179 VPWR.n1178 VPWR.n726 0.0605
R12180 VPWR.n1741 VPWR 0.0605
R12181 VPWR.n1129 VPWR.n1128 0.0605
R12182 VPWR VPWR.n1837 0.0605
R12183 VPWR.n1968 VPWR.n1967 0.0605
R12184 VPWR.n1963 VPWR.n1962 0.0605
R12185 VPWR.n2914 VPWR.n2913 0.0605
R12186 VPWR.n2893 VPWR.n2892 0.0605
R12187 VPWR.n2793 VPWR.n2792 0.0605
R12188 VPWR.n469 VPWR.n468 0.0605
R12189 VPWR.n505 VPWR.n504 0.0605
R12190 VPWR.n569 VPWR.n568 0.0605
R12191 VPWR.n3031 VPWR.n3030 0.0605
R12192 VPWR.n450 VPWR.n449 0.0605
R12193 VPWR VPWR.n1672 0.05975
R12194 VPWR.n684 VPWR 0.05975
R12195 VPWR.n3020 VPWR 0.05975
R12196 VPWR VPWR.n1045 0.059
R12197 VPWR VPWR.n1049 0.059
R12198 VPWR VPWR.n1349 0.059
R12199 VPWR.n1440 VPWR 0.059
R12200 VPWR VPWR.n1267 0.059
R12201 VPWR.n1256 VPWR 0.059
R12202 VPWR VPWR.n1251 0.059
R12203 VPWR.n1706 VPWR 0.059
R12204 VPWR VPWR.n1711 0.059
R12205 VPWR.n1081 VPWR 0.059
R12206 VPWR VPWR.n1080 0.059
R12207 VPWR VPWR.n1828 0.059
R12208 VPWR.n1990 VPWR 0.059
R12209 VPWR.n1986 VPWR 0.059
R12210 VPWR VPWR.n1985 0.059
R12211 VPWR VPWR.n1981 0.059
R12212 VPWR.n2029 VPWR 0.059
R12213 VPWR VPWR.n2024 0.059
R12214 VPWR VPWR.n2020 0.059
R12215 VPWR VPWR.n2720 0.059
R12216 VPWR.n2721 VPWR 0.059
R12217 VPWR.n2725 VPWR 0.059
R12218 VPWR.n2074 VPWR 0.059
R12219 VPWR VPWR.n2073 0.059
R12220 VPWR.n2070 VPWR 0.059
R12221 VPWR VPWR.n2069 0.059
R12222 VPWR VPWR.n2706 0.059
R12223 VPWR VPWR.n2702 0.059
R12224 VPWR VPWR.n493 0.059
R12225 VPWR.n494 VPWR 0.059
R12226 VPWR.n1899 VPWR 0.059
R12227 VPWR.n1656 VPWR 0.05825
R12228 VPWR.n3230 VPWR.n3229 0.0575
R12229 VPWR.n3253 VPWR.n3252 0.0575
R12230 VPWR.n1192 VPWR 0.0575
R12231 VPWR.n1735 VPWR.n1734 0.0575
R12232 VPWR.n3193 VPWR.n3192 0.0575
R12233 VPWR.n2838 VPWR.n2837 0.0575
R12234 VPWR.n2786 VPWR.n2785 0.0575
R12235 VPWR.n2707 VPWR.n197 0.0575
R12236 VPWR.n548 VPWR.n547 0.0575
R12237 VPWR VPWR.n1382 0.05675
R12238 VPWR VPWR.n571 0.05675
R12239 VPWR VPWR.n1383 0.056
R12240 VPWR.n1275 VPWR.n1274 0.056
R12241 VPWR.n1273 VPWR.n1272 0.056
R12242 VPWR.n1340 VPWR.n1339 0.056
R12243 VPWR.n1338 VPWR.n1337 0.056
R12244 VPWR.n1168 VPWR.n1167 0.056
R12245 VPWR.n1166 VPWR.n1165 0.056
R12246 VPWR.n1164 VPWR.n1163 0.056
R12247 VPWR.n1162 VPWR.n1161 0.056
R12248 VPWR.n1160 VPWR.n1159 0.056
R12249 VPWR.n1214 VPWR.n1213 0.056
R12250 VPWR.n1970 VPWR.n1969 0.056
R12251 VPWR.n2133 VPWR.n2132 0.056
R12252 VPWR.n2275 VPWR.n2274 0.056
R12253 VPWR.n2278 VPWR.n284 0.056
R12254 VPWR.n2711 VPWR.n2710 0.056
R12255 VPWR.n1328 VPWR.n1327 0.05525
R12256 VPWR.n3447 VPWR 0.0545
R12257 VPWR.n3448 VPWR 0.0545
R12258 VPWR.n3462 VPWR 0.0545
R12259 VPWR.n3463 VPWR 0.0545
R12260 VPWR.n3477 VPWR 0.0545
R12261 VPWR.n3478 VPWR 0.0545
R12262 VPWR.n3492 VPWR 0.0545
R12263 VPWR.n3493 VPWR 0.0545
R12264 VPWR.n3507 VPWR 0.0545
R12265 VPWR.n3508 VPWR 0.0545
R12266 VPWR.n3522 VPWR 0.0545
R12267 VPWR.n3523 VPWR 0.0545
R12268 VPWR.n3537 VPWR 0.0545
R12269 VPWR.n3538 VPWR 0.0545
R12270 VPWR.n3552 VPWR 0.0545
R12271 VPWR.n3553 VPWR 0.0545
R12272 VPWR.n3567 VPWR 0.0545
R12273 VPWR.n3568 VPWR 0.0545
R12274 VPWR.n3582 VPWR 0.0545
R12275 VPWR.n3583 VPWR 0.0545
R12276 VPWR.n3597 VPWR 0.0545
R12277 VPWR.n3598 VPWR 0.0545
R12278 VPWR.n3612 VPWR 0.0545
R12279 VPWR.n3613 VPWR 0.0545
R12280 VPWR.n3627 VPWR 0.0545
R12281 VPWR.n3628 VPWR 0.0545
R12282 VPWR.n3642 VPWR 0.0545
R12283 VPWR.n3643 VPWR 0.0545
R12284 VPWR.n3657 VPWR 0.0545
R12285 VPWR.n3658 VPWR 0.0545
R12286 VPWR.n3672 VPWR 0.0545
R12287 VPWR.n3673 VPWR 0.0545
R12288 VPWR VPWR.n1516 0.0545
R12289 VPWR VPWR.n1587 0.0545
R12290 VPWR VPWR.n1584 0.0545
R12291 VPWR VPWR.n1578 0.0545
R12292 VPWR.n1530 VPWR 0.0545
R12293 VPWR VPWR.n1567 0.0545
R12294 VPWR VPWR.n1564 0.0545
R12295 VPWR VPWR.n1557 0.0545
R12296 VPWR VPWR.n1551 0.0545
R12297 VPWR VPWR.n1547 0.0545
R12298 VPWR VPWR.n1353 0.0545
R12299 VPWR VPWR.n1355 0.0545
R12300 VPWR.n1456 VPWR 0.0545
R12301 VPWR VPWR.n1007 0.0545
R12302 VPWR VPWR.n976 0.0545
R12303 VPWR.n3382 VPWR 0.0545
R12304 VPWR.n3384 VPWR 0.0545
R12305 VPWR.n3417 VPWR 0.0545
R12306 VPWR VPWR.n1328 0.0545
R12307 VPWR VPWR.n1322 0.0545
R12308 VPWR VPWR.n1321 0.0545
R12309 VPWR VPWR.n1305 0.0545
R12310 VPWR VPWR.n1300 0.0545
R12311 VPWR VPWR.n1291 0.0545
R12312 VPWR VPWR.n1653 0.0545
R12313 VPWR VPWR.n1643 0.0545
R12314 VPWR VPWR.n903 0.0545
R12315 VPWR.n870 VPWR 0.0545
R12316 VPWR.n3337 VPWR 0.0545
R12317 VPWR VPWR.n3341 0.0545
R12318 VPWR VPWR.n3360 0.0545
R12319 VPWR VPWR.n1247 0.0545
R12320 VPWR VPWR.n1244 0.0545
R12321 VPWR VPWR.n1239 0.0545
R12322 VPWR VPWR.n1237 0.0545
R12323 VPWR VPWR.n1232 0.0545
R12324 VPWR VPWR.n1690 0.0545
R12325 VPWR VPWR.n779 0.0545
R12326 VPWR VPWR.n775 0.0545
R12327 VPWR VPWR.n771 0.0545
R12328 VPWR.n770 VPWR 0.0545
R12329 VPWR VPWR.n767 0.0545
R12330 VPWR VPWR.n766 0.0545
R12331 VPWR VPWR.n764 0.0545
R12332 VPWR.n3236 VPWR 0.0545
R12333 VPWR VPWR.n122 0.0545
R12334 VPWR VPWR.n3294 0.0545
R12335 VPWR VPWR.n3288 0.0545
R12336 VPWR VPWR.n3274 0.0545
R12337 VPWR.n1712 VPWR 0.0545
R12338 VPWR.n1723 VPWR 0.0545
R12339 VPWR.n1725 VPWR 0.0545
R12340 VPWR.n1726 VPWR 0.0545
R12341 VPWR VPWR.n1769 0.0545
R12342 VPWR.n1811 VPWR.n1810 0.0545
R12343 VPWR VPWR.n1792 0.0545
R12344 VPWR VPWR.n3215 0.0545
R12345 VPWR VPWR.n3177 0.0545
R12346 VPWR VPWR.n1153 0.0545
R12347 VPWR VPWR.n1150 0.0545
R12348 VPWR VPWR.n1143 0.0545
R12349 VPWR VPWR.n1138 0.0545
R12350 VPWR.n1137 VPWR 0.0545
R12351 VPWR VPWR.n1132 0.0545
R12352 VPWR VPWR.n1116 0.0545
R12353 VPWR VPWR.n678 0.0545
R12354 VPWR VPWR.n675 0.0545
R12355 VPWR VPWR.n652 0.0545
R12356 VPWR VPWR.n639 0.0545
R12357 VPWR.n3111 VPWR 0.0545
R12358 VPWR VPWR.n1933 0.0545
R12359 VPWR VPWR.n1928 0.0545
R12360 VPWR VPWR.n1927 0.0545
R12361 VPWR VPWR.n1978 0.0545
R12362 VPWR VPWR.n1973 0.0545
R12363 VPWR VPWR.n1968 0.0545
R12364 VPWR VPWR.n1955 0.0545
R12365 VPWR VPWR.n1954 0.0545
R12366 VPWR.n2841 VPWR 0.0545
R12367 VPWR VPWR.n2893 0.0545
R12368 VPWR.n2129 VPWR 0.0545
R12369 VPWR.n2139 VPWR 0.0545
R12370 VPWR VPWR.n2013 0.0545
R12371 VPWR VPWR.n2008 0.0545
R12372 VPWR VPWR.n2007 0.0545
R12373 VPWR VPWR.n2048 0.0545
R12374 VPWR VPWR.n2016 0.0545
R12375 VPWR VPWR.n194 0.0545
R12376 VPWR.n2715 VPWR 0.0545
R12377 VPWR.n2717 VPWR 0.0545
R12378 VPWR VPWR.n2805 0.0545
R12379 VPWR VPWR.n2062 0.0545
R12380 VPWR VPWR.n2059 0.0545
R12381 VPWR VPWR.n2056 0.0545
R12382 VPWR VPWR.n2096 0.0545
R12383 VPWR VPWR.n2081 0.0545
R12384 VPWR.n2700 VPWR.n2699 0.0545
R12385 VPWR VPWR.n2694 0.0545
R12386 VPWR VPWR.n2687 0.0545
R12387 VPWR VPWR.n233 0.0545
R12388 VPWR.n460 VPWR 0.0545
R12389 VPWR.n490 VPWR 0.0545
R12390 VPWR VPWR.n1864 0.0545
R12391 VPWR VPWR.n581 0.0545
R12392 VPWR VPWR.n569 0.0545
R12393 VPWR VPWR.n555 0.0545
R12394 VPWR VPWR.n553 0.0545
R12395 VPWR VPWR.n551 0.0545
R12396 VPWR.n3039 VPWR 0.0545
R12397 VPWR.n362 VPWR 0.0545
R12398 VPWR VPWR.n366 0.0545
R12399 VPWR VPWR.n364 0.0545
R12400 VPWR VPWR.n363 0.0545
R12401 VPWR VPWR.n1919 0.0545
R12402 VPWR VPWR.n1901 0.0545
R12403 VPWR.n1891 VPWR 0.0545
R12404 VPWR VPWR.n1890 0.0545
R12405 VPWR.n1889 VPWR 0.0545
R12406 VPWR VPWR.n1888 0.0545
R12407 VPWR VPWR.n1886 0.0545
R12408 VPWR VPWR.n455 0.0545
R12409 VPWR VPWR.n438 0.0545
R12410 VPWR VPWR.n437 0.0545
R12411 VPWR.n2932 VPWR 0.0545
R12412 VPWR.n2933 VPWR 0.0545
R12413 VPWR.n2938 VPWR 0.0545
R12414 VPWR.n269 VPWR 0.0545
R12415 VPWR.n272 VPWR 0.0545
R12416 VPWR.n3704 VPWR 0.0545
R12417 VPWR VPWR.n2424 0.0545
R12418 VPWR VPWR.n2423 0.0545
R12419 VPWR VPWR.n2418 0.0545
R12420 VPWR VPWR.n2443 0.0545
R12421 VPWR VPWR.n2588 0.0545
R12422 VPWR.n19 VPWR 0.0545
R12423 VPWR VPWR.n3736 0.0545
R12424 VPWR VPWR.n1618 0.05375
R12425 VPWR.n1261 VPWR 0.053
R12426 VPWR.n1705 VPWR.n1704 0.053
R12427 VPWR.n1374 VPWR.n1373 0.05225
R12428 VPWR.n3352 VPWR 0.05225
R12429 VPWR.n1755 VPWR.n1754 0.05225
R12430 VPWR.n3017 VPWR 0.05225
R12431 VPWR.n1527 VPWR.n104 0.0515
R12432 VPWR.n1364 VPWR.n1363 0.0515
R12433 VPWR.n1673 VPWR 0.0515
R12434 VPWR.n3291 VPWR.n3290 0.0515
R12435 VPWR.n1717 VPWR.n1716 0.0515
R12436 VPWR.n1797 VPWR.n1796 0.0515
R12437 VPWR.n3161 VPWR.n169 0.0515
R12438 VPWR.n1136 VPWR.n1135 0.0515
R12439 VPWR.n1844 VPWR 0.0515
R12440 VPWR.n694 VPWR.n693 0.0515
R12441 VPWR.n3158 VPWR.n3157 0.0515
R12442 VPWR.n476 VPWR 0.0515
R12443 VPWR.n499 VPWR.n498 0.0515
R12444 VPWR VPWR.n1876 0.0515
R12445 VPWR.n1847 VPWR 0.0515
R12446 VPWR.n3069 VPWR.n3068 0.0515
R12447 VPWR.n1618 VPWR.n1617 0.05
R12448 VPWR VPWR.n3243 0.05
R12449 VPWR.n3196 VPWR.n3195 0.05
R12450 VPWR VPWR.n3454 0.04925
R12451 VPWR VPWR.n3469 0.04925
R12452 VPWR VPWR.n3484 0.04925
R12453 VPWR VPWR.n3499 0.04925
R12454 VPWR VPWR.n3514 0.04925
R12455 VPWR VPWR.n3529 0.04925
R12456 VPWR VPWR.n3544 0.04925
R12457 VPWR VPWR.n3559 0.04925
R12458 VPWR VPWR.n3574 0.04925
R12459 VPWR VPWR.n3589 0.04925
R12460 VPWR VPWR.n3604 0.04925
R12461 VPWR VPWR.n3619 0.04925
R12462 VPWR VPWR.n3634 0.04925
R12463 VPWR VPWR.n3649 0.04925
R12464 VPWR VPWR.n3664 0.04925
R12465 VPWR VPWR.n3679 0.04925
R12466 VPWR.n1494 VPWR 0.04925
R12467 VPWR VPWR.n1501 0.04925
R12468 VPWR.n1538 VPWR 0.04925
R12469 VPWR.n3392 VPWR 0.04925
R12470 VPWR.n3407 VPWR 0.04925
R12471 VPWR.n3425 VPWR 0.04925
R12472 VPWR VPWR.n3439 0.04925
R12473 VPWR VPWR.n3362 0.04925
R12474 VPWR VPWR.n3278 0.04925
R12475 VPWR VPWR.n160 0.04925
R12476 VPWR VPWR.n1147 0.04925
R12477 VPWR VPWR.n1115 0.04925
R12478 VPWR.n3124 VPWR 0.04925
R12479 VPWR VPWR.n3148 0.04925
R12480 VPWR VPWR.n1997 0.04925
R12481 VPWR VPWR.n1996 0.04925
R12482 VPWR VPWR.n1945 0.04925
R12483 VPWR.n2844 VPWR 0.04925
R12484 VPWR VPWR.n2884 0.04925
R12485 VPWR.n357 VPWR 0.04925
R12486 VPWR.n2150 VPWR 0.04925
R12487 VPWR VPWR.n2171 0.04925
R12488 VPWR.n294 VPWR 0.04925
R12489 VPWR VPWR.n335 0.04925
R12490 VPWR VPWR.n2392 0.04925
R12491 VPWR VPWR.n2403 0.04925
R12492 VPWR VPWR.n2414 0.04925
R12493 VPWR VPWR.n275 0.04925
R12494 VPWR VPWR.n2223 0.04925
R12495 VPWR VPWR.n2381 0.04925
R12496 VPWR VPWR.n2372 0.04925
R12497 VPWR VPWR.n2363 0.04925
R12498 VPWR VPWR.n2353 0.04925
R12499 VPWR VPWR.n2344 0.04925
R12500 VPWR VPWR.n2334 0.04925
R12501 VPWR VPWR.n2041 0.04925
R12502 VPWR VPWR.n2038 0.04925
R12503 VPWR VPWR.n2736 0.04925
R12504 VPWR VPWR.n2754 0.04925
R12505 VPWR VPWR.n2089 0.04925
R12506 VPWR VPWR.n2087 0.04925
R12507 VPWR VPWR.n2690 0.04925
R12508 VPWR VPWR.n2673 0.04925
R12509 VPWR VPWR.n2659 0.04925
R12510 VPWR VPWR.n2648 0.04925
R12511 VPWR VPWR.n243 0.04925
R12512 VPWR VPWR.n225 0.04925
R12513 VPWR VPWR.n211 0.04925
R12514 VPWR VPWR.n3059 0.04925
R12515 VPWR VPWR.n1908 0.04925
R12516 VPWR.n431 VPWR.n430 0.04925
R12517 VPWR VPWR.n3007 0.04925
R12518 VPWR VPWR.n3004 0.04925
R12519 VPWR VPWR.n2992 0.04925
R12520 VPWR VPWR.n2982 0.04925
R12521 VPWR VPWR.n2973 0.04925
R12522 VPWR VPWR.n2963 0.04925
R12523 VPWR.n2458 VPWR 0.04925
R12524 VPWR.n2468 VPWR 0.04925
R12525 VPWR VPWR.n2474 0.04925
R12526 VPWR VPWR.n2494 0.04925
R12527 VPWR VPWR.n2485 0.04925
R12528 VPWR.n2608 VPWR 0.04925
R12529 VPWR VPWR.n2614 0.04925
R12530 VPWR VPWR.n2636 0.04925
R12531 VPWR VPWR.n2627 0.04925
R12532 VPWR VPWR.n3831 0.04925
R12533 VPWR VPWR.n3822 0.04925
R12534 VPWR.n43 VPWR 0.04925
R12535 VPWR.n52 VPWR 0.04925
R12536 VPWR VPWR.n3771 0.04925
R12537 VPWR VPWR.n3762 0.04925
R12538 VPWR.n3689 VPWR 0.04925
R12539 VPWR.n3698 VPWR 0.04925
R12540 VPWR VPWR.n3711 0.04925
R12541 VPWR VPWR.n2450 0.04925
R12542 VPWR VPWR.n2446 0.04925
R12543 VPWR VPWR.n2432 0.04925
R12544 VPWR.n2514 VPWR 0.04925
R12545 VPWR VPWR.n2525 0.04925
R12546 VPWR VPWR.n2592 0.04925
R12547 VPWR VPWR.n2579 0.04925
R12548 VPWR VPWR.n2564 0.04925
R12549 VPWR VPWR.n2548 0.04925
R12550 VPWR.n14 VPWR 0.04925
R12551 VPWR VPWR.n25 0.04925
R12552 VPWR VPWR.n3805 0.04925
R12553 VPWR VPWR.n3788 0.04925
R12554 VPWR.n67 VPWR 0.04925
R12555 VPWR.n78 VPWR 0.04925
R12556 VPWR VPWR.n3746 0.04925
R12557 VPWR VPWR.n3728 0.04925
R12558 VPWR VPWR.n92 0.04925
R12559 VPWR.n1448 VPWR 0.0485
R12560 VPWR.n909 VPWR.n908 0.0485
R12561 VPWR.n881 VPWR.n880 0.0485
R12562 VPWR VPWR.n1699 0.0485
R12563 VPWR.n3282 VPWR.n3281 0.0485
R12564 VPWR.n1733 VPWR.n1732 0.0485
R12565 VPWR VPWR.n1803 0.0485
R12566 VPWR.n2764 VPWR.n2763 0.0485
R12567 VPWR.n220 VPWR.n219 0.0485
R12568 VPWR.n418 VPWR.n417 0.0485
R12569 VPWR.n680 VPWR.n679 0.04775
R12570 VPWR.n1560 VPWR 0.047
R12571 VPWR VPWR.n1351 0.047
R12572 VPWR VPWR.n1326 0.047
R12573 VPWR VPWR.n1324 0.047
R12574 VPWR.n862 VPWR 0.047
R12575 VPWR VPWR.n3323 0.047
R12576 VPWR VPWR.n1259 0.047
R12577 VPWR VPWR.n3305 0.047
R12578 VPWR VPWR.n1802 0.047
R12579 VPWR VPWR.n3180 0.047
R12580 VPWR VPWR.n1121 0.047
R12581 VPWR VPWR.n659 0.047
R12582 VPWR VPWR.n1935 0.047
R12583 VPWR VPWR.n1958 0.047
R12584 VPWR VPWR.n1952 0.047
R12585 VPWR.n2385 VPWR 0.047
R12586 VPWR.n2396 VPWR 0.047
R12587 VPWR.n2407 VPWR 0.047
R12588 VPWR VPWR.n2015 0.047
R12589 VPWR.n2730 VPWR 0.047
R12590 VPWR VPWR.n2067 0.047
R12591 VPWR VPWR.n556 0.047
R12592 VPWR VPWR.n1912 0.047
R12593 VPWR VPWR.n1906 0.047
R12594 VPWR.n1447 VPWR 0.0455
R12595 VPWR.n1446 VPWR.n1445 0.0455
R12596 VPWR.n859 VPWR.n858 0.0455
R12597 VPWR.n1677 VPWR.n1676 0.0455
R12598 VPWR.n814 VPWR.n813 0.0455
R12599 VPWR.n2915 VPWR 0.0455
R12600 VPWR.n600 VPWR.n599 0.0455
R12601 VPWR.n400 VPWR 0.0455
R12602 VPWR.n3396 VPWR 0.04475
R12603 VPWR VPWR.n3433 0.04475
R12604 VPWR VPWR.n3173 0.04475
R12605 VPWR VPWR.n164 0.04475
R12606 VPWR VPWR.n646 0.04475
R12607 VPWR VPWR.n3142 0.04475
R12608 VPWR VPWR.n3152 0.04475
R12609 VPWR.n2110 VPWR 0.04475
R12610 VPWR.n2127 VPWR 0.04475
R12611 VPWR VPWR.n2165 0.04475
R12612 VPWR VPWR.n2175 0.04475
R12613 VPWR.n305 VPWR 0.04475
R12614 VPWR VPWR.n329 0.04475
R12615 VPWR VPWR.n2266 0.04475
R12616 VPWR VPWR.n2248 0.04475
R12617 VPWR VPWR.n339 0.04475
R12618 VPWR VPWR.n2306 0.04475
R12619 VPWR VPWR.n2288 0.04475
R12620 VPWR.n2194 VPWR 0.04475
R12621 VPWR VPWR.n2217 0.04475
R12622 VPWR VPWR.n2227 0.04475
R12623 VPWR VPWR.n2824 0.04475
R12624 VPWR VPWR.n2807 0.04475
R12625 VPWR VPWR.n2777 0.04475
R12626 VPWR VPWR.n2758 0.04475
R12627 VPWR VPWR.n2665 0.04475
R12628 VPWR VPWR.n253 0.04475
R12629 VPWR VPWR.n215 0.04475
R12630 VPWR VPWR.n3053 0.04475
R12631 VPWR VPWR.n3099 0.04475
R12632 VPWR VPWR.n3081 0.04475
R12633 VPWR VPWR.n3063 0.04475
R12634 VPWR VPWR.n2431 0.04475
R12635 VPWR VPWR.n2522 0.04475
R12636 VPWR VPWR.n2577 0.04475
R12637 VPWR VPWR.n2543 0.04475
R12638 VPWR VPWR.n22 0.04475
R12639 VPWR VPWR.n3781 0.04475
R12640 VPWR.n82 VPWR 0.04475
R12641 VPWR VPWR.n3719 0.04475
R12642 VPWR.n2323 VPWR 0.04325
R12643 VPWR.n1451 VPWR 0.0425
R12644 VPWR.n1429 VPWR 0.0425
R12645 VPWR.n1647 VPWR.n1646 0.0425
R12646 VPWR.n1681 VPWR.n1680 0.0425
R12647 VPWR.n1787 VPWR.n134 0.0425
R12648 VPWR.n2858 VPWR.n2857 0.0425
R12649 VPWR.n2919 VPWR.n2918 0.0425
R12650 VPWR.n405 VPWR.n404 0.0425
R12651 VPWR.n2942 VPWR.n2941 0.0425
R12652 VPWR.n2393 VPWR 0.04175
R12653 VPWR.n2404 VPWR 0.04175
R12654 VPWR.n2415 VPWR 0.04175
R12655 VPWR.n2382 VPWR 0.04175
R12656 VPWR VPWR.n2457 0.04175
R12657 VPWR.n993 VPWR.n992 0.041
R12658 VPWR.n1264 VPWR 0.041
R12659 VPWR.n1288 VPWR.n1287 0.04025
R12660 VPWR.n3174 VPWR 0.04025
R12661 VPWR.n647 VPWR 0.04025
R12662 VPWR.n3143 VPWR 0.04025
R12663 VPWR VPWR.n2109 0.04025
R12664 VPWR.n2166 VPWR 0.04025
R12665 VPWR VPWR.n304 0.04025
R12666 VPWR.n330 VPWR 0.04025
R12667 VPWR.n2267 VPWR 0.04025
R12668 VPWR.n2249 VPWR 0.04025
R12669 VPWR.n2307 VPWR 0.04025
R12670 VPWR.n2289 VPWR 0.04025
R12671 VPWR VPWR.n2193 0.04025
R12672 VPWR.n2218 VPWR 0.04025
R12673 VPWR.n2825 VPWR 0.04025
R12674 VPWR.n2778 VPWR 0.04025
R12675 VPWR.n1853 VPWR 0.04025
R12676 VPWR.n3054 VPWR 0.04025
R12677 VPWR.n3100 VPWR 0.04025
R12678 VPWR.n3082 VPWR 0.04025
R12679 VPWR VPWR.n1884 0.04025
R12680 VPWR.n983 VPWR.n982 0.0395
R12681 VPWR VPWR.n3249 0.0395
R12682 VPWR.n1195 VPWR 0.0395
R12683 VPWR VPWR.n1187 0.0395
R12684 VPWR VPWR.n1832 0.0395
R12685 VPWR.n1943 VPWR.n1942 0.0395
R12686 VPWR.n2831 VPWR.n189 0.0395
R12687 VPWR.n1872 VPWR.n1871 0.0395
R12688 VPWR.n434 VPWR.n433 0.0395
R12689 VPWR VPWR.n1058 0.03875
R12690 VPWR VPWR.n1068 0.03875
R12691 VPWR VPWR.n1473 0.03875
R12692 VPWR VPWR.n1485 0.03875
R12693 VPWR VPWR.n1827 0.03875
R12694 VPWR.n575 VPWR 0.03875
R12695 VPWR.n901 VPWR.n900 0.038
R12696 VPWR.n1239 VPWR 0.038
R12697 VPWR.n1976 VPWR 0.038
R12698 VPWR VPWR.n2846 0.038
R12699 VPWR.n2018 VPWR 0.038
R12700 VPWR.n2064 VPWR 0.038
R12701 VPWR.n2692 VPWR 0.038
R12702 VPWR VPWR.n459 0.038
R12703 VPWR VPWR.n1860 0.038
R12704 VPWR.n570 VPWR 0.038
R12705 VPWR VPWR.n361 0.038
R12706 VPWR.n368 VPWR 0.038
R12707 VPWR.n455 VPWR 0.038
R12708 VPWR VPWR.n3701 0.038
R12709 VPWR.n2426 VPWR 0.038
R12710 VPWR.n1698 VPWR.n1697 0.0365
R12711 VPWR.n3187 VPWR.n3186 0.0365
R12712 VPWR.n2763 VPWR.n2761 0.0365
R12713 VPWR.n3020 VPWR.n3019 0.0365
R12714 VPWR VPWR.n3123 0.03575
R12715 VPWR VPWR.n356 0.03575
R12716 VPWR VPWR.n2149 0.03575
R12717 VPWR VPWR.n293 0.03575
R12718 VPWR.n276 VPWR 0.03575
R12719 VPWR.n2042 VPWR 0.03575
R12720 VPWR.n2737 VPWR 0.03575
R12721 VPWR.n3008 VPWR 0.03575
R12722 VPWR.n1441 VPWR 0.03425
R12723 VPWR.n1427 VPWR.n1426 0.03425
R12724 VPWR.n864 VPWR.n863 0.03425
R12725 VPWR.n1453 VPWR.n1452 0.0335
R12726 VPWR.n1623 VPWR 0.0335
R12727 VPWR.n1303 VPWR 0.0335
R12728 VPWR.n897 VPWR.n896 0.0335
R12729 VPWR.n892 VPWR.n891 0.0335
R12730 VPWR.n868 VPWR.n867 0.0335
R12731 VPWR.n3334 VPWR.n3333 0.0335
R12732 VPWR VPWR.n789 0.0335
R12733 VPWR.n1208 VPWR 0.0335
R12734 VPWR.n3220 VPWR.n3219 0.0335
R12735 VPWR.n3190 VPWR.n3189 0.0335
R12736 VPWR.n3162 VPWR.n3161 0.0335
R12737 VPWR.n3158 VPWR.n171 0.0335
R12738 VPWR.n509 VPWR 0.0335
R12739 VPWR.n501 VPWR 0.0335
R12740 VPWR.n1854 VPWR 0.0335
R12741 VPWR VPWR.n1850 0.0335
R12742 VPWR.n3070 VPWR.n3069 0.0335
R12743 VPWR.n1894 VPWR.n1893 0.0335
R12744 VPWR VPWR.n423 0.0335
R12745 VPWR.n1284 VPWR 0.03275
R12746 VPWR.n1199 VPWR.n1198 0.032
R12747 VPWR.n1190 VPWR.n1189 0.032
R12748 VPWR.n1184 VPWR.n1183 0.032
R12749 VPWR.n3203 VPWR 0.03125
R12750 VPWR VPWR.n3446 0.0305
R12751 VPWR VPWR.n3461 0.0305
R12752 VPWR VPWR.n3476 0.0305
R12753 VPWR VPWR.n3491 0.0305
R12754 VPWR VPWR.n3506 0.0305
R12755 VPWR VPWR.n3521 0.0305
R12756 VPWR VPWR.n3536 0.0305
R12757 VPWR VPWR.n3551 0.0305
R12758 VPWR VPWR.n3566 0.0305
R12759 VPWR VPWR.n3581 0.0305
R12760 VPWR VPWR.n3596 0.0305
R12761 VPWR VPWR.n3611 0.0305
R12762 VPWR VPWR.n3626 0.0305
R12763 VPWR VPWR.n3641 0.0305
R12764 VPWR VPWR.n3656 0.0305
R12765 VPWR VPWR.n3671 0.0305
R12766 VPWR.n1487 VPWR 0.0305
R12767 VPWR VPWR.n1514 0.0305
R12768 VPWR VPWR.n1603 0.0305
R12769 VPWR VPWR.n1461 0.0305
R12770 VPWR VPWR.n1456 0.0305
R12771 VPWR VPWR.n1455 0.0305
R12772 VPWR.n1442 VPWR 0.0305
R12773 VPWR.n1627 VPWR 0.0305
R12774 VPWR.n1615 VPWR 0.0305
R12775 VPWR.n1016 VPWR 0.0305
R12776 VPWR VPWR.n3381 0.0305
R12777 VPWR.n1335 VPWR 0.0305
R12778 VPWR.n1322 VPWR 0.0305
R12779 VPWR.n1306 VPWR 0.0305
R12780 VPWR.n1298 VPWR 0.0305
R12781 VPWR.n1293 VPWR 0.0305
R12782 VPWR.n1660 VPWR.n1659 0.0305
R12783 VPWR VPWR.n1649 0.0305
R12784 VPWR.n878 VPWR.n877 0.0305
R12785 VPWR.n872 VPWR 0.0305
R12786 VPWR.n3347 VPWR.n3346 0.0305
R12787 VPWR VPWR.n1226 0.0305
R12788 VPWR.n1223 VPWR 0.0305
R12789 VPWR.n1219 VPWR 0.0305
R12790 VPWR.n1258 VPWR 0.0305
R12791 VPWR.n1245 VPWR 0.0305
R12792 VPWR.n1244 VPWR 0.0305
R12793 VPWR.n1694 VPWR 0.0305
R12794 VPWR.n762 VPWR 0.0305
R12795 VPWR.n1170 VPWR 0.0305
R12796 VPWR.n1210 VPWR 0.0305
R12797 VPWR VPWR.n1205 0.0305
R12798 VPWR.n1181 VPWR 0.0305
R12799 VPWR VPWR.n1180 0.0305
R12800 VPWR VPWR.n1712 0.0305
R12801 VPWR VPWR.n1718 0.0305
R12802 VPWR.n1719 VPWR 0.0305
R12803 VPWR.n3178 VPWR 0.0305
R12804 VPWR.n3173 VPWR 0.0305
R12805 VPWR.n1154 VPWR 0.0305
R12806 VPWR VPWR.n1130 0.0305
R12807 VPWR.n1117 VPWR 0.0305
R12808 VPWR VPWR.n688 0.0305
R12809 VPWR.n676 VPWR 0.0305
R12810 VPWR.n675 VPWR 0.0305
R12811 VPWR.n653 VPWR 0.0305
R12812 VPWR.n646 VPWR 0.0305
R12813 VPWR VPWR.n3116 0.0305
R12814 VPWR.n3142 VPWR 0.0305
R12815 VPWR.n1929 VPWR 0.0305
R12816 VPWR VPWR.n1964 0.0305
R12817 VPWR.n1957 VPWR 0.0305
R12818 VPWR.n1956 VPWR 0.0305
R12819 VPWR.n2901 VPWR.n2900 0.0305
R12820 VPWR VPWR.n2110 0.0305
R12821 VPWR VPWR.n2136 0.0305
R12822 VPWR VPWR.n2142 0.0305
R12823 VPWR.n2165 VPWR 0.0305
R12824 VPWR VPWR.n305 0.0305
R12825 VPWR.n329 VPWR 0.0305
R12826 VPWR.n2266 VPWR 0.0305
R12827 VPWR.n2248 VPWR 0.0305
R12828 VPWR.n2306 VPWR 0.0305
R12829 VPWR.n2288 VPWR 0.0305
R12830 VPWR VPWR.n2194 0.0305
R12831 VPWR.n2217 VPWR 0.0305
R12832 VPWR.n2009 VPWR 0.0305
R12833 VPWR.n2031 VPWR 0.0305
R12834 VPWR.n2744 VPWR 0.0305
R12835 VPWR.n2824 VPWR 0.0305
R12836 VPWR.n2783 VPWR 0.0305
R12837 VPWR.n2777 VPWR 0.0305
R12838 VPWR VPWR.n462 0.0305
R12839 VPWR.n463 VPWR 0.0305
R12840 VPWR VPWR.n506 0.0305
R12841 VPWR.n503 VPWR 0.0305
R12842 VPWR.n497 VPWR 0.0305
R12843 VPWR.n561 VPWR 0.0305
R12844 VPWR VPWR.n3038 0.0305
R12845 VPWR.n3053 VPWR 0.0305
R12846 VPWR.n3099 VPWR 0.0305
R12847 VPWR.n3081 VPWR 0.0305
R12848 VPWR.n1902 VPWR 0.0305
R12849 VPWR VPWR.n451 0.0305
R12850 VPWR.n448 VPWR 0.0305
R12851 VPWR.n441 VPWR 0.0305
R12852 VPWR.n438 VPWR 0.0305
R12853 VPWR.n424 VPWR 0.0305
R12854 VPWR.n2941 VPWR 0.0305
R12855 VPWR.n1292 VPWR 0.02975
R12856 VPWR VPWR.n1282 0.02975
R12857 VPWR VPWR.n1748 0.02975
R12858 VPWR.n1749 VPWR 0.02975
R12859 VPWR.n1041 VPWR.n1040 0.029
R12860 VPWR.n1043 VPWR.n1042 0.029
R12861 VPWR.n1470 VPWR.n1033 0.029
R12862 VPWR.n1469 VPWR 0.029
R12863 VPWR.n1626 VPWR 0.029
R12864 VPWR VPWR.n3384 0.029
R12865 VPWR VPWR.n3396 0.029
R12866 VPWR VPWR.n3415 0.029
R12867 VPWR.n1263 VPWR.n1262 0.029
R12868 VPWR.n1707 VPWR.n728 0.029
R12869 VPWR.n1212 VPWR 0.029
R12870 VPWR VPWR.n1714 0.029
R12871 VPWR VPWR.n1727 0.029
R12872 VPWR.n1127 VPWR.n1126 0.029
R12873 VPWR.n1106 VPWR 0.029
R12874 VPWR.n1993 VPWR 0.029
R12875 VPWR.n2275 VPWR.n285 0.029
R12876 VPWR.n2279 VPWR.n2278 0.029
R12877 VPWR.n2363 VPWR.n2362 0.029
R12878 VPWR.n2085 VPWR 0.029
R12879 VPWR.n2079 VPWR.n2078 0.029
R12880 VPWR.n2077 VPWR.n2076 0.029
R12881 VPWR.n2683 VPWR 0.029
R12882 VPWR.n2656 VPWR 0.029
R12883 VPWR.n253 VPWR 0.029
R12884 VPWR.n235 VPWR 0.029
R12885 VPWR.n478 VPWR.n477 0.029
R12886 VPWR.n480 VPWR.n479 0.029
R12887 VPWR.n482 VPWR.n481 0.029
R12888 VPWR.n484 VPWR.n483 0.029
R12889 VPWR.n486 VPWR.n485 0.029
R12890 VPWR.n488 VPWR.n487 0.029
R12891 VPWR.n1878 VPWR 0.029
R12892 VPWR VPWR.n2459 0.029
R12893 VPWR.n2500 VPWR.n265 0.029
R12894 VPWR.n2446 VPWR 0.029
R12895 VPWR.n2503 VPWR.n263 0.029
R12896 VPWR VPWR.n2504 0.029
R12897 VPWR VPWR.n2519 0.029
R12898 VPWR.n2591 VPWR 0.029
R12899 VPWR.n2574 VPWR 0.029
R12900 VPWR.n2558 VPWR 0.029
R12901 VPWR VPWR.n16 0.029
R12902 VPWR.n21 VPWR 0.029
R12903 VPWR.n3798 VPWR 0.029
R12904 VPWR VPWR.n70 0.029
R12905 VPWR VPWR.n82 0.029
R12906 VPWR.n3738 VPWR 0.029
R12907 VPWR.n1667 VPWR.n1666 0.02825
R12908 VPWR.n1707 VPWR.n1706 0.0275
R12909 VPWR.n1676 VPWR.n816 0.0275
R12910 VPWR.n3231 VPWR 0.0275
R12911 VPWR.n1711 VPWR.n1710 0.0275
R12912 VPWR.n1789 VPWR.n1788 0.0275
R12913 VPWR.n685 VPWR.n684 0.0275
R12914 VPWR.n683 VPWR.n682 0.0275
R12915 VPWR.n1881 VPWR.n1880 0.0275
R12916 VPWR VPWR.n1227 0.026
R12917 VPWR.n1222 VPWR 0.026
R12918 VPWR.n1218 VPWR 0.026
R12919 VPWR.n1209 VPWR 0.026
R12920 VPWR VPWR.n1206 0.026
R12921 VPWR VPWR.n1202 0.026
R12922 VPWR.n1201 VPWR 0.026
R12923 VPWR.n1125 VPWR 0.026
R12924 VPWR VPWR.n1965 0.026
R12925 VPWR VPWR.n1961 0.026
R12926 VPWR.n1960 VPWR 0.026
R12927 VPWR.n466 VPWR 0.026
R12928 VPWR VPWR.n467 0.026
R12929 VPWR.n470 VPWR 0.026
R12930 VPWR VPWR.n472 0.026
R12931 VPWR VPWR.n491 0.026
R12932 VPWR VPWR.n507 0.026
R12933 VPWR.n502 VPWR 0.026
R12934 VPWR VPWR.n452 0.026
R12935 VPWR.n447 VPWR 0.026
R12936 VPWR.n2923 VPWR 0.026
R12937 VPWR.n2891 VPWR 0.02525
R12938 VPWR.n2936 VPWR.n2935 0.02525
R12939 VPWR.n1000 VPWR.n999 0.0245
R12940 VPWR.n1342 VPWR 0.0245
R12941 VPWR.n1308 VPWR.n1307 0.0245
R12942 VPWR.n1649 VPWR.n1648 0.0245
R12943 VPWR VPWR.n886 0.0245
R12944 VPWR.n3332 VPWR.n3331 0.0245
R12945 VPWR VPWR.n3344 0.0245
R12946 VPWR.n1254 VPWR.n1253 0.0245
R12947 VPWR.n3225 VPWR.n3224 0.0245
R12948 VPWR VPWR.n3292 0.0245
R12949 VPWR.n1156 VPWR.n1155 0.0245
R12950 VPWR.n1134 VPWR.n1133 0.0245
R12951 VPWR.n1988 VPWR.n1987 0.0245
R12952 VPWR.n1984 VPWR.n1983 0.0245
R12953 VPWR.n1940 VPWR.n189 0.0245
R12954 VPWR.n2027 VPWR.n2026 0.0245
R12955 VPWR.n2723 VPWR.n2722 0.0245
R12956 VPWR.n2072 VPWR.n2071 0.0245
R12957 VPWR.n2705 VPWR.n2704 0.0245
R12958 VPWR.n474 VPWR.n473 0.0245
R12959 VPWR.n496 VPWR.n495 0.0245
R12960 VPWR.n1897 VPWR.n1896 0.0245
R12961 VPWR.n446 VPWR 0.0245
R12962 VPWR.n1669 VPWR 0.02375
R12963 VPWR.n1347 VPWR.n1053 0.023
R12964 VPWR VPWR.n1463 0.023
R12965 VPWR.n876 VPWR 0.023
R12966 VPWR.n3319 VPWR.n119 0.023
R12967 VPWR.n1702 VPWR.n1701 0.023
R12968 VPWR.n1215 VPWR.n1159 0.023
R12969 VPWR.n1834 VPWR.n1833 0.023
R12970 VPWR.n471 VPWR.n470 0.023
R12971 VPWR.n2949 VPWR 0.023
R12972 VPWR.n3285 VPWR 0.02225
R12973 VPWR VPWR.n1434 0.0215
R12974 VPWR VPWR.n990 0.0215
R12975 VPWR.n3367 VPWR.n3366 0.0215
R12976 VPWR.n1682 VPWR 0.0215
R12977 VPWR.n3309 VPWR.n3308 0.0215
R12978 VPWR VPWR.n3220 0.0215
R12979 VPWR.n3184 VPWR.n3183 0.0215
R12980 VPWR.n2909 VPWR.n2908 0.0215
R12981 VPWR.n2184 VPWR.n2183 0.0215
R12982 VPWR.n2239 VPWR.n347 0.0215
R12983 VPWR.n2236 VPWR.n2235 0.0215
R12984 VPWR.n2669 VPWR.n2668 0.0215
R12985 VPWR.n423 VPWR.n422 0.0215
R12986 VPWR.n2926 VPWR.n2925 0.0215
R12987 VPWR.n2599 VPWR.n2598 0.0215
R12988 VPWR VPWR.n2843 0.02075
R12989 VPWR.n1512 VPWR 0.0200652
R12990 VPWR.n1361 VPWR 0.0200652
R12991 VPWR.n883 VPWR 0.0200652
R12992 VPWR.n3198 VPWR 0.0200652
R12993 VPWR.n2909 VPWR 0.0200652
R12994 VPWR.n3457 VPWR.n3444 0.0185
R12995 VPWR.n3472 VPWR.n3459 0.0185
R12996 VPWR.n3487 VPWR.n3474 0.0185
R12997 VPWR.n3502 VPWR.n3489 0.0185
R12998 VPWR.n3517 VPWR.n3504 0.0185
R12999 VPWR.n3532 VPWR.n3519 0.0185
R13000 VPWR.n3547 VPWR.n3534 0.0185
R13001 VPWR.n3562 VPWR.n3549 0.0185
R13002 VPWR.n3577 VPWR.n3564 0.0185
R13003 VPWR.n3592 VPWR.n3579 0.0185
R13004 VPWR.n3607 VPWR.n3594 0.0185
R13005 VPWR.n3622 VPWR.n3609 0.0185
R13006 VPWR.n3637 VPWR.n3624 0.0185
R13007 VPWR.n3652 VPWR.n3639 0.0185
R13008 VPWR.n3667 VPWR.n3654 0.0185
R13009 VPWR.n3682 VPWR.n3669 0.0185
R13010 VPWR.n1605 VPWR.n1018 0.0185
R13011 VPWR.n1543 VPWR.n95 0.0185
R13012 VPWR.n1608 VPWR.n1607 0.0185
R13013 VPWR.n3442 VPWR.n96 0.0185
R13014 VPWR VPWR.n1336 0.0185
R13015 VPWR.n1662 VPWR.n1661 0.0185
R13016 VPWR.n3328 VPWR.n3327 0.0185
R13017 VPWR VPWR.n1228 0.0185
R13018 VPWR.n797 VPWR.n796 0.0185
R13019 VPWR.n793 VPWR.n792 0.0185
R13020 VPWR VPWR.n1171 0.0185
R13021 VPWR VPWR.n1207 0.0185
R13022 VPWR VPWR.n603 0.0185
R13023 VPWR.n696 VPWR.n695 0.0185
R13024 VPWR VPWR.n508 0.0185
R13025 VPWR VPWR.n585 0.0185
R13026 VPWR VPWR.n453 0.0185
R13027 VPWR.n3836 VPWR.n4 0.0185
R13028 VPWR.n3714 VPWR.n3684 0.0185
R13029 VPWR.n3840 VPWR.n3839 0.0185
R13030 VPWR.n3718 VPWR.n3717 0.0185
R13031 VPWR.n1318 VPWR.n1317 0.01775
R13032 VPWR VPWR.n784 0.01775
R13033 VPWR VPWR.n591 0.01775
R13034 VPWR.n1622 VPWR 0.017
R13035 VPWR.n906 VPWR 0.017
R13036 VPWR.n1131 VPWR 0.017
R13037 VPWR VPWR.n1217 0.01625
R13038 VPWR.n1720 VPWR 0.01625
R13039 VPWR VPWR.n1124 0.01625
R13040 VPWR VPWR.n1922 0.01625
R13041 VPWR.n888 VPWR.n887 0.0155
R13042 VPWR VPWR.n686 0.0155
R13043 VPWR.n3279 VPWR 0.01475
R13044 VPWR.n1423 VPWR 0.014
R13045 VPWR.n1639 VPWR.n1638 0.014
R13046 VPWR VPWR.n3302 0.014
R13047 VPWR.n2798 VPWR.n2797 0.014
R13048 VPWR VPWR.n786 0.01325
R13049 VPWR.n786 VPWR.n785 0.01325
R13050 VPWR.n590 VPWR.n589 0.01325
R13051 VPWR VPWR.n1358 0.0125
R13052 VPWR VPWR.n1466 0.0125
R13053 VPWR VPWR.n1442 0.0125
R13054 VPWR.n1413 VPWR 0.0125
R13055 VPWR.n1610 VPWR 0.0125
R13056 VPWR.n1008 VPWR 0.0125
R13057 VPWR.n999 VPWR 0.0125
R13058 VPWR.n995 VPWR 0.0125
R13059 VPWR.n984 VPWR 0.0125
R13060 VPWR VPWR.n3378 0.0125
R13061 VPWR.n1316 VPWR 0.0125
R13062 VPWR VPWR.n1283 0.0125
R13063 VPWR.n904 VPWR 0.0125
R13064 VPWR.n890 VPWR 0.0125
R13065 VPWR.n3321 VPWR 0.0125
R13066 VPWR.n3322 VPWR.n3321 0.0125
R13067 VPWR VPWR.n3329 0.0125
R13068 VPWR.n3351 VPWR 0.0125
R13069 VPWR VPWR.n3350 0.0125
R13070 VPWR.n3365 VPWR 0.0125
R13071 VPWR VPWR.n3364 0.0125
R13072 VPWR.n1234 VPWR 0.0125
R13073 VPWR VPWR.n1230 0.0125
R13074 VPWR VPWR.n1689 0.0125
R13075 VPWR VPWR.n802 0.0125
R13076 VPWR.n787 VPWR 0.0125
R13077 VPWR.n783 VPWR.n782 0.0125
R13078 VPWR.n772 VPWR 0.0125
R13079 VPWR VPWR.n3314 0.0125
R13080 VPWR.n3307 VPWR 0.0125
R13081 VPWR VPWR.n3306 0.0125
R13082 VPWR.n3295 VPWR 0.0125
R13083 VPWR.n3277 VPWR 0.0125
R13084 VPWR.n1197 VPWR 0.0125
R13085 VPWR VPWR.n1185 0.0125
R13086 VPWR.n1800 VPWR 0.0125
R13087 VPWR.n1799 VPWR.n1798 0.0125
R13088 VPWR.n1788 VPWR 0.0125
R13089 VPWR.n3212 VPWR 0.0125
R13090 VPWR.n3204 VPWR 0.0125
R13091 VPWR.n3194 VPWR 0.0125
R13092 VPWR.n3182 VPWR 0.0125
R13093 VPWR VPWR.n3181 0.0125
R13094 VPWR VPWR.n1114 0.0125
R13095 VPWR.n669 VPWR.n668 0.0125
R13096 VPWR.n661 VPWR 0.0125
R13097 VPWR VPWR.n1944 0.0125
R13098 VPWR VPWR.n2858 0.0125
R13099 VPWR.n2856 VPWR.n2855 0.0125
R13100 VPWR.n2852 VPWR.n184 0.0125
R13101 VPWR.n2918 VPWR 0.0125
R13102 VPWR.n2899 VPWR 0.0125
R13103 VPWR.n2892 VPWR 0.0125
R13104 VPWR VPWR.n2799 0.0125
R13105 VPWR VPWR.n1874 0.0125
R13106 VPWR VPWR.n3031 0.0125
R13107 VPWR VPWR.n435 0.0125
R13108 VPWR.n407 VPWR 0.0125
R13109 VPWR.n406 VPWR 0.0125
R13110 VPWR.n3015 VPWR 0.0125
R13111 VPWR.n3445 VPWR 0.01175
R13112 VPWR.n3460 VPWR 0.01175
R13113 VPWR.n3475 VPWR 0.01175
R13114 VPWR.n3490 VPWR 0.01175
R13115 VPWR.n3505 VPWR 0.01175
R13116 VPWR.n3520 VPWR 0.01175
R13117 VPWR.n3535 VPWR 0.01175
R13118 VPWR.n3550 VPWR 0.01175
R13119 VPWR.n3565 VPWR 0.01175
R13120 VPWR.n3580 VPWR 0.01175
R13121 VPWR.n3595 VPWR 0.01175
R13122 VPWR.n3610 VPWR 0.01175
R13123 VPWR.n3625 VPWR 0.01175
R13124 VPWR.n3640 VPWR 0.01175
R13125 VPWR.n3655 VPWR 0.01175
R13126 VPWR.n3670 VPWR 0.01175
R13127 VPWR VPWR.n1428 0.01175
R13128 VPWR VPWR.n980 0.01175
R13129 VPWR.n970 VPWR.n969 0.01175
R13130 VPWR VPWR.n1269 0.01175
R13131 VPWR VPWR.n1296 0.01175
R13132 VPWR VPWR.n1289 0.01175
R13133 VPWR VPWR.n1692 0.01175
R13134 VPWR VPWR.n1082 0.01175
R13135 VPWR VPWR.n1140 0.01175
R13136 VPWR VPWR.n2890 0.01175
R13137 VPWR.n349 VPWR 0.01175
R13138 VPWR.n286 VPWR 0.01175
R13139 VPWR VPWR.n283 0.01175
R13140 VPWR.n2713 VPWR 0.01175
R13141 VPWR.n3032 VPWR 0.01175
R13142 VPWR VPWR.n442 0.01175
R13143 VPWR VPWR.n425 0.01175
R13144 VPWR.n1286 VPWR.n1285 0.01025
R13145 VPWR.n1651 VPWR.n1650 0.0095
R13146 VPWR.n883 VPWR.n882 0.0095
R13147 VPWR.n809 VPWR.n808 0.0095
R13148 VPWR.n671 VPWR.n670 0.0095
R13149 VPWR.n2834 VPWR.n2833 0.0095
R13150 VPWR.n2790 VPWR.n2789 0.0095
R13151 VPWR.n1857 VPWR.n1856 0.0095
R13152 VPWR.n428 VPWR.n427 0.0095
R13153 VPWR.n1010 VPWR 0.008
R13154 VPWR.n2928 VPWR 0.008
R13155 VPWR.n1444 VPWR 0.00725
R13156 VPWR.n1331 VPWR 0.00725
R13157 VPWR.n1652 VPWR 0.00725
R13158 VPWR.n1813 VPWR 0.00725
R13159 VPWR.n1839 VPWR 0.00725
R13160 VPWR.n1437 VPWR 0.0065
R13161 VPWR VPWR.n1011 0.0065
R13162 VPWR VPWR.n988 0.0065
R13163 VPWR.n895 VPWR.n894 0.0065
R13164 VPWR.n3326 VPWR 0.0065
R13165 VPWR.n1684 VPWR 0.0065
R13166 VPWR.n811 VPWR 0.0065
R13167 VPWR VPWR.n3310 0.0065
R13168 VPWR.n1769 VPWR 0.0065
R13169 VPWR.n3221 VPWR.n134 0.0065
R13170 VPWR VPWR.n2897 0.0065
R13171 VPWR.n2102 VPWR.n2101 0.0065
R13172 VPWR.n297 VPWR.n296 0.0065
R13173 VPWR.n2315 VPWR.n2314 0.0065
R13174 VPWR.n1868 VPWR 0.0065
R13175 VPWR.n1924 VPWR.n1923 0.0065
R13176 VPWR.n1473 VPWR.n1472 0.00575
R13177 VPWR.n1344 VPWR 0.00575
R13178 VPWR.n1804 VPWR 0.00575
R13179 VPWR.n682 VPWR 0.00575
R13180 VPWR.n565 VPWR 0.00575
R13181 VPWR.n2934 VPWR.n2933 0.00575
R13182 VPWR.n1221 VPWR.n1220 0.005
R13183 VPWR.n1696 VPWR.n1695 0.005
R13184 VPWR.n1147 VPWR.n1146 0.005
R13185 VPWR.n2920 VPWR.n2919 0.005
R13186 VPWR.n2134 VPWR.n2133 0.005
R13187 VPWR.n2729 VPWR.n2728 0.005
R13188 VPWR.n465 VPWR.n464 0.005
R13189 VPWR.n580 VPWR.n579 0.005
R13190 VPWR.n1071 VPWR 0.0035
R13191 VPWR.n1070 VPWR 0.0035
R13192 VPWR.n1635 VPWR 0.0035
R13193 VPWR.n986 VPWR.n985 0.0035
R13194 VPWR VPWR.n977 0.0035
R13195 VPWR.n1673 VPWR.n818 0.0035
R13196 VPWR.n3241 VPWR 0.0035
R13197 VPWR.n3248 VPWR.n3247 0.0035
R13198 VPWR VPWR.n2377 0.0035
R13199 VPWR.n1848 VPWR.n1847 0.0035
R13200 VPWR VPWR.n2999 0.0035
R13201 VPWR.n2466 VPWR 0.0035
R13202 VPWR VPWR.n3700 0.0035
R13203 VPWR.n972 VPWR.n971 0.00275
R13204 VPWR.n3450 VPWR 0.002
R13205 VPWR.n3465 VPWR 0.002
R13206 VPWR.n3480 VPWR 0.002
R13207 VPWR.n3495 VPWR 0.002
R13208 VPWR.n3510 VPWR 0.002
R13209 VPWR.n3525 VPWR 0.002
R13210 VPWR.n3540 VPWR 0.002
R13211 VPWR.n3555 VPWR 0.002
R13212 VPWR.n3570 VPWR 0.002
R13213 VPWR.n3585 VPWR 0.002
R13214 VPWR.n3600 VPWR 0.002
R13215 VPWR.n3615 VPWR 0.002
R13216 VPWR.n3630 VPWR 0.002
R13217 VPWR.n3645 VPWR 0.002
R13218 VPWR.n3660 VPWR 0.002
R13219 VPWR.n3675 VPWR 0.002
R13220 VPWR VPWR.n1077 0.002
R13221 VPWR VPWR.n1069 0.002
R13222 VPWR.n1474 VPWR 0.002
R13223 VPWR.n1482 VPWR 0.002
R13224 VPWR.n1489 VPWR 0.002
R13225 VPWR.n1506 VPWR 0.002
R13226 VPWR.n1509 VPWR 0.002
R13227 VPWR.n1521 VPWR 0.002
R13228 VPWR VPWR.n1018 0.002
R13229 VPWR VPWR.n1599 0.002
R13230 VPWR VPWR.n1591 0.002
R13231 VPWR.n1590 VPWR.n1589 0.002
R13232 VPWR VPWR.n1582 0.002
R13233 VPWR VPWR.n1573 0.002
R13234 VPWR.n1570 VPWR 0.002
R13235 VPWR VPWR.n1562 0.002
R13236 VPWR VPWR.n1553 0.002
R13237 VPWR VPWR.n1545 0.002
R13238 VPWR.n1350 VPWR 0.002
R13239 VPWR.n1359 VPWR 0.002
R13240 VPWR.n1384 VPWR 0.002
R13241 VPWR VPWR.n1468 0.002
R13242 VPWR VPWR.n1460 0.002
R13243 VPWR VPWR.n1451 0.002
R13244 VPWR VPWR.n1439 0.002
R13245 VPWR VPWR.n1429 0.002
R13246 VPWR VPWR.n1424 0.002
R13247 VPWR.n1418 VPWR 0.002
R13248 VPWR VPWR.n1637 0.002
R13249 VPWR VPWR.n1621 0.002
R13250 VPWR VPWR.n1608 0.002
R13251 VPWR VPWR.n1009 0.002
R13252 VPWR VPWR.n1005 0.002
R13253 VPWR VPWR.n994 0.002
R13254 VPWR.n992 VPWR.n991 0.002
R13255 VPWR VPWR.n981 0.002
R13256 VPWR VPWR.n966 0.002
R13257 VPWR.n3385 VPWR 0.002
R13258 VPWR.n3387 VPWR 0.002
R13259 VPWR.n3397 VPWR 0.002
R13260 VPWR.n3414 VPWR 0.002
R13261 VPWR.n3416 VPWR 0.002
R13262 VPWR.n3434 VPWR 0.002
R13263 VPWR VPWR.n1341 0.002
R13264 VPWR VPWR.n1325 0.002
R13265 VPWR VPWR.n1309 0.002
R13266 VPWR VPWR.n1295 0.002
R13267 VPWR VPWR.n1668 0.002
R13268 VPWR VPWR.n1655 0.002
R13269 VPWR VPWR.n907 0.002
R13270 VPWR VPWR.n895 0.002
R13271 VPWR VPWR.n878 0.002
R13272 VPWR VPWR.n865 0.002
R13273 VPWR.n3320 VPWR.n3319 0.002
R13274 VPWR.n3324 VPWR 0.002
R13275 VPWR.n3353 VPWR 0.002
R13276 VPWR VPWR.n3369 0.002
R13277 VPWR VPWR.n1260 0.002
R13278 VPWR VPWR.n1240 0.002
R13279 VPWR VPWR.n1703 0.002
R13280 VPWR VPWR.n1686 0.002
R13281 VPWR VPWR.n815 0.002
R13282 VPWR VPWR.n798 0.002
R13283 VPWR VPWR.n783 0.002
R13284 VPWR.n3228 VPWR 0.002
R13285 VPWR.n3254 VPWR 0.002
R13286 VPWR VPWR.n3312 0.002
R13287 VPWR VPWR.n3301 0.002
R13288 VPWR VPWR.n3286 0.002
R13289 VPWR VPWR.n1211 0.002
R13290 VPWR VPWR.n1191 0.002
R13291 VPWR.n1715 VPWR 0.002
R13292 VPWR.n1728 VPWR 0.002
R13293 VPWR.n1744 VPWR 0.002
R13294 VPWR.n1777 VPWR 0.002
R13295 VPWR VPWR.n1811 0.002
R13296 VPWR VPWR.n1799 0.002
R13297 VPWR VPWR.n3218 0.002
R13298 VPWR VPWR.n3205 0.002
R13299 VPWR VPWR.n3191 0.002
R13300 VPWR VPWR.n3175 0.002
R13301 VPWR VPWR.n165 0.002
R13302 VPWR VPWR.n1141 0.002
R13303 VPWR.n1126 VPWR 0.002
R13304 VPWR VPWR.n1122 0.002
R13305 VPWR VPWR.n1107 0.002
R13306 VPWR VPWR.n1841 0.002
R13307 VPWR.n1830 VPWR 0.002
R13308 VPWR VPWR.n1829 0.002
R13309 VPWR.n1824 VPWR.n1823 0.002
R13310 VPWR.n1819 VPWR.n1818 0.002
R13311 VPWR VPWR.n694 0.002
R13312 VPWR VPWR.n681 0.002
R13313 VPWR VPWR.n665 0.002
R13314 VPWR VPWR.n648 0.002
R13315 VPWR.n3110 VPWR.n3109 0.002
R13316 VPWR.n3114 VPWR 0.002
R13317 VPWR.n3144 VPWR 0.002
R13318 VPWR VPWR.n3153 0.002
R13319 VPWR VPWR.n2002 0.002
R13320 VPWR VPWR.n1992 0.002
R13321 VPWR.n1974 VPWR 0.002
R13322 VPWR VPWR.n1972 0.002
R13323 VPWR VPWR.n1953 0.002
R13324 VPWR.n2832 VPWR 0.002
R13325 VPWR.n2860 VPWR 0.002
R13326 VPWR.n2917 VPWR 0.002
R13327 VPWR VPWR.n2916 0.002
R13328 VPWR VPWR.n2903 0.002
R13329 VPWR.n2108 VPWR 0.002
R13330 VPWR.n2126 VPWR 0.002
R13331 VPWR.n2140 VPWR 0.002
R13332 VPWR.n2167 VPWR 0.002
R13333 VPWR VPWR.n2176 0.002
R13334 VPWR.n303 VPWR 0.002
R13335 VPWR.n331 VPWR 0.002
R13336 VPWR VPWR.n2268 0.002
R13337 VPWR VPWR.n2250 0.002
R13338 VPWR VPWR.n340 0.002
R13339 VPWR VPWR.n2308 0.002
R13340 VPWR VPWR.n2290 0.002
R13341 VPWR.n2192 VPWR 0.002
R13342 VPWR.n2219 VPWR 0.002
R13343 VPWR VPWR.n2228 0.002
R13344 VPWR.n2319 VPWR 0.002
R13345 VPWR.n2323 VPWR 0.002
R13346 VPWR VPWR.n2368 0.002
R13347 VPWR VPWR.n2358 0.002
R13348 VPWR VPWR.n2349 0.002
R13349 VPWR VPWR.n2339 0.002
R13350 VPWR VPWR.n2051 0.002
R13351 VPWR VPWR.n2033 0.002
R13352 VPWR.n2712 VPWR 0.002
R13353 VPWR.n2746 VPWR 0.002
R13354 VPWR VPWR.n2826 0.002
R13355 VPWR VPWR.n2808 0.002
R13356 VPWR VPWR.n2795 0.002
R13357 VPWR VPWR.n2779 0.002
R13358 VPWR VPWR.n2759 0.002
R13359 VPWR VPWR.n2092 0.002
R13360 VPWR VPWR.n2084 0.002
R13361 VPWR VPWR.n2080 0.002
R13362 VPWR.n2707 VPWR 0.002
R13363 VPWR VPWR.n2700 0.002
R13364 VPWR VPWR.n2685 0.002
R13365 VPWR VPWR.n2682 0.002
R13366 VPWR VPWR.n2664 0.002
R13367 VPWR VPWR.n2655 0.002
R13368 VPWR VPWR.n2653 0.002
R13369 VPWR VPWR.n252 0.002
R13370 VPWR VPWR.n236 0.002
R13371 VPWR VPWR.n234 0.002
R13372 VPWR VPWR.n216 0.002
R13373 VPWR.n475 VPWR 0.002
R13374 VPWR.n510 VPWR 0.002
R13375 VPWR VPWR.n1877 0.002
R13376 VPWR VPWR.n1861 0.002
R13377 VPWR VPWR.n598 0.002
R13378 VPWR VPWR.n588 0.002
R13379 VPWR VPWR.n573 0.002
R13380 VPWR VPWR.n558 0.002
R13381 VPWR.n3026 VPWR 0.002
R13382 VPWR.n3055 VPWR 0.002
R13383 VPWR.n3106 VPWR.n3105 0.002
R13384 VPWR VPWR.n3101 0.002
R13385 VPWR VPWR.n3083 0.002
R13386 VPWR VPWR.n3064 0.002
R13387 VPWR.n369 VPWR 0.002
R13388 VPWR VPWR.n1913 0.002
R13389 VPWR VPWR.n1895 0.002
R13390 VPWR.n1884 VPWR 0.002
R13391 VPWR VPWR.n454 0.002
R13392 VPWR VPWR.n445 0.002
R13393 VPWR VPWR.n429 0.002
R13394 VPWR VPWR.n421 0.002
R13395 VPWR VPWR.n416 0.002
R13396 VPWR VPWR.n405 0.002
R13397 VPWR.n2925 VPWR 0.002
R13398 VPWR.n2929 VPWR 0.002
R13399 VPWR.n2950 VPWR 0.002
R13400 VPWR VPWR.n3018 0.002
R13401 VPWR VPWR.n3013 0.002
R13402 VPWR VPWR.n2997 0.002
R13403 VPWR VPWR.n2987 0.002
R13404 VPWR VPWR.n2978 0.002
R13405 VPWR VPWR.n2968 0.002
R13406 VPWR.n2460 VPWR 0.002
R13407 VPWR.n2479 VPWR 0.002
R13408 VPWR VPWR.n2499 0.002
R13409 VPWR VPWR.n2490 0.002
R13410 VPWR.n2603 VPWR 0.002
R13411 VPWR.n2619 VPWR 0.002
R13412 VPWR VPWR.n2641 0.002
R13413 VPWR VPWR.n2632 0.002
R13414 VPWR VPWR.n4 0.002
R13415 VPWR VPWR.n3827 0.002
R13416 VPWR VPWR.n3818 0.002
R13417 VPWR.n3817 VPWR.n7 0.002
R13418 VPWR.n47 VPWR 0.002
R13419 VPWR.n56 VPWR 0.002
R13420 VPWR VPWR.n3767 0.002
R13421 VPWR VPWR.n3758 0.002
R13422 VPWR.n3693 VPWR 0.002
R13423 VPWR.n3706 VPWR 0.002
R13424 VPWR VPWR.n2451 0.002
R13425 VPWR VPWR.n2445 0.002
R13426 VPWR VPWR.n2437 0.002
R13427 VPWR.n2505 VPWR 0.002
R13428 VPWR.n2515 VPWR 0.002
R13429 VPWR.n2534 VPWR 0.002
R13430 VPWR VPWR.n2597 0.002
R13431 VPWR VPWR.n2590 0.002
R13432 VPWR VPWR.n2584 0.002
R13433 VPWR VPWR.n2573 0.002
R13434 VPWR VPWR.n2561 0.002
R13435 VPWR VPWR.n2557 0.002
R13436 VPWR VPWR.n3840 0.002
R13437 VPWR.n17 VPWR 0.002
R13438 VPWR.n30 VPWR 0.002
R13439 VPWR VPWR.n9 0.002
R13440 VPWR.n3814 VPWR.n3813 0.002
R13441 VPWR VPWR.n3800 0.002
R13442 VPWR VPWR.n3797 0.002
R13443 VPWR VPWR.n3780 0.002
R13444 VPWR.n71 VPWR 0.002
R13445 VPWR.n73 VPWR 0.002
R13446 VPWR.n84 VPWR 0.002
R13447 VPWR VPWR.n3739 0.002
R13448 VPWR VPWR.n3737 0.002
R13449 VPWR VPWR.n3720 0.002
R13450 VGND.n3700 VGND.n38 57115.1
R13451 VGND.n3700 VGND.n21 57115.1
R13452 VGND.n3700 VGND.n37 57115.1
R13453 VGND.n3700 VGND.n36 57115.1
R13454 VGND.n3704 VGND.n3700 57115.1
R13455 VGND.n3700 VGND.n40 57115.1
R13456 VGND.n2953 VGND.n2952 10144.3
R13457 VGND.t4341 VGND.t2012 3324.2
R13458 VGND.t2672 VGND.t699 3324.2
R13459 VGND.t699 VGND.t4405 3324.2
R13460 VGND.t4405 VGND.t5551 3324.2
R13461 VGND.t5858 VGND.t3950 3324.2
R13462 VGND.t3950 VGND.t1274 3324.2
R13463 VGND.t1274 VGND.t4798 3324.2
R13464 VGND.t4798 VGND.t4616 3324.2
R13465 VGND.t4616 VGND.t4020 3324.2
R13466 VGND.t4020 VGND.t1961 3324.2
R13467 VGND.t1961 VGND.t2931 3324.2
R13468 VGND.t2441 VGND.t5763 3324.2
R13469 VGND.t4925 VGND.t2441 3324.2
R13470 VGND.t2424 VGND.t4925 3324.2
R13471 VGND.t1959 VGND.t2424 3324.2
R13472 VGND.t5309 VGND.t1959 3324.2
R13473 VGND.t5042 VGND.t5309 3324.2
R13474 VGND.t1163 VGND.t5042 3324.2
R13475 VGND.t4767 VGND.t1302 3324.2
R13476 VGND.t4012 VGND.t4767 3324.2
R13477 VGND.t3952 VGND.t4012 3324.2
R13478 VGND.t2033 VGND.t3952 3324.2
R13479 VGND.t2548 VGND.t2033 3324.2
R13480 VGND.t2803 VGND.t2548 3324.2
R13481 VGND.t2808 VGND.t2803 3324.2
R13482 VGND.t5942 VGND.t4584 3324.2
R13483 VGND.t4584 VGND.t1258 3324.2
R13484 VGND.t1258 VGND.t5833 3324.2
R13485 VGND.t5833 VGND.t2483 3324.2
R13486 VGND.t2483 VGND.t3732 3324.2
R13487 VGND.t3732 VGND.t5641 3324.2
R13488 VGND.t5641 VGND.t4258 3324.2
R13489 VGND.t4593 VGND.t2776 3324.2
R13490 VGND.t2776 VGND.t3159 3324.2
R13491 VGND.t3159 VGND.t2666 3324.2
R13492 VGND.t2666 VGND.t5546 3324.2
R13493 VGND.t5546 VGND.t627 3324.2
R13494 VGND.t627 VGND.t4239 3324.2
R13495 VGND.t4239 VGND.t1967 3324.2
R13496 VGND.t6753 VGND.t2128 3324.2
R13497 VGND.t6085 VGND.t6753 3324.2
R13498 VGND.t903 VGND.t6085 3324.2
R13499 VGND.t4985 VGND.t903 3324.2
R13500 VGND.t4400 VGND.t4985 3324.2
R13501 VGND.t2530 VGND.t4400 3324.2
R13502 VGND.t3999 VGND.t2530 3324.2
R13503 VGND.t4582 VGND.t2138 3324.2
R13504 VGND.t406 VGND.t4582 3324.2
R13505 VGND.t1551 VGND.t406 3324.2
R13506 VGND.t3366 VGND.t1551 3324.2
R13507 VGND.t4747 VGND.t3366 3324.2
R13508 VGND.t4387 VGND.t4747 3324.2
R13509 VGND.t625 VGND.t4387 3324.2
R13510 VGND.t3179 VGND.t4663 3324.2
R13511 VGND.t4663 VGND.t5258 3324.2
R13512 VGND.t5258 VGND.t836 3324.2
R13513 VGND.t836 VGND.t3207 3324.2
R13514 VGND.t3207 VGND.t615 3324.2
R13515 VGND.t615 VGND.t4630 3324.2
R13516 VGND.t4630 VGND.t2040 3324.2
R13517 VGND.t2206 VGND.t3283 3324.2
R13518 VGND.t3283 VGND.t1718 3324.2
R13519 VGND.t1718 VGND.t5483 3324.2
R13520 VGND.t5483 VGND.t3086 3324.2
R13521 VGND.t3086 VGND.t4708 3324.2
R13522 VGND.t4708 VGND.t3790 3324.2
R13523 VGND.t3790 VGND.t3110 3324.2
R13524 VGND.t1620 VGND.t3765 3324.2
R13525 VGND.t1734 VGND.t1620 3324.2
R13526 VGND.t2553 VGND.t1734 3324.2
R13527 VGND.t4098 VGND.t2553 3324.2
R13528 VGND.t5528 VGND.t4098 3324.2
R13529 VGND.t2975 VGND.t5528 3324.2
R13530 VGND.t3349 VGND.t2975 3324.2
R13531 VGND.t6161 VGND.t1935 3324.2
R13532 VGND.t6813 VGND.t6161 3324.2
R13533 VGND.t5988 VGND.t6813 3324.2
R13534 VGND.t5496 VGND.t5988 3324.2
R13535 VGND.t1583 VGND.t5496 3324.2
R13536 VGND.t6029 VGND.t1583 3324.2
R13537 VGND.t2832 VGND.t6029 3324.2
R13538 VGND.t356 VGND.t935 3324.2
R13539 VGND.t3400 VGND.t356 3324.2
R13540 VGND.t5487 VGND.t3400 3324.2
R13541 VGND.t5290 VGND.t5487 3324.2
R13542 VGND.t5964 VGND.t5290 3324.2
R13543 VGND.t410 VGND.t5964 3324.2
R13544 VGND.t5189 VGND.t410 3324.2
R13545 VGND.t4667 VGND.t4777 3324.2
R13546 VGND.t4144 VGND.t4667 3324.2
R13547 VGND.t6760 VGND.t4144 3324.2
R13548 VGND.t2836 VGND.t6760 3324.2
R13549 VGND.t931 VGND.t2836 3324.2
R13550 VGND.t3465 VGND.t931 3324.2
R13551 VGND.t5519 VGND.t3465 3324.2
R13552 VGND.t4790 VGND.t3692 3324.2
R13553 VGND.t3692 VGND.t1418 3324.2
R13554 VGND.t1418 VGND.t4436 3324.2
R13555 VGND.t4436 VGND.t2853 3324.2
R13556 VGND.t2853 VGND.t5489 3324.2
R13557 VGND.t5489 VGND.t2747 3324.2
R13558 VGND.t2747 VGND.t5966 3324.2
R13559 VGND.t4409 VGND.t5863 3324.2
R13560 VGND.t5863 VGND.t3317 3324.2
R13561 VGND.t3317 VGND.t4627 3324.2
R13562 VGND.t4627 VGND.t4578 3324.2
R13563 VGND.t4578 VGND.t442 3324.2
R13564 VGND.t442 VGND.t2546 3324.2
R13565 VGND.t2546 VGND.t5340 3324.2
R13566 VGND.t5617 VGND.t5944 3324.2
R13567 VGND.t3372 VGND.t5617 3324.2
R13568 VGND.t337 VGND.t3372 3324.2
R13569 VGND.t5934 VGND.t337 3324.2
R13570 VGND.t2114 VGND.t5934 3324.2
R13571 VGND.t1327 VGND.t2114 3324.2
R13572 VGND.t2202 VGND.t1327 3324.2
R13573 VGND.t1300 VGND.t4084 3324.2
R13574 VGND.t2173 VGND.t1300 3324.2
R13575 VGND.t69 VGND.t2173 3324.2
R13576 VGND.t635 VGND.t69 3324.2
R13577 VGND.t4572 VGND.t635 3324.2
R13578 VGND.t3487 VGND.t4572 3324.2
R13579 VGND.t1442 VGND.t3487 3324.2
R13580 VGND.n3700 VGND.n3699 3179.33
R13581 VGND.n380 VGND.t5858 2493.15
R13582 VGND.t5763 VGND.n3019 2493.15
R13583 VGND.t1302 VGND.n3020 2493.15
R13584 VGND.n3021 VGND.t5942 2493.15
R13585 VGND.n372 VGND.t4593 2493.15
R13586 VGND.t2128 VGND.n3124 2493.15
R13587 VGND.t2138 VGND.n3125 2493.15
R13588 VGND.n3126 VGND.t3179 2493.15
R13589 VGND.n365 VGND.t2206 2493.15
R13590 VGND.t3765 VGND.n3230 2493.15
R13591 VGND.t1935 VGND.n3231 2493.15
R13592 VGND.t935 VGND.n3232 2493.15
R13593 VGND.t4777 VGND.n3233 2493.15
R13594 VGND.n3234 VGND.t4790 2493.15
R13595 VGND.n1 VGND.t4409 2493.15
R13596 VGND.t5944 VGND.n3776 2493.15
R13597 VGND.t4084 VGND.n3777 2493.15
R13598 VGND.n3700 VGND.n39 2317.79
R13599 VGND VGND.t4341 2166.67
R13600 VGND VGND.t2672 2166.67
R13601 VGND.t63 VGND.t555 2068.18
R13602 VGND.t2588 VGND.t63 2068.18
R13603 VGND.t1289 VGND.t2588 2068.18
R13604 VGND.t5330 VGND.t1289 2068.18
R13605 VGND.t1316 VGND.t5330 2068.18
R13606 VGND.t650 VGND.t1316 2068.18
R13607 VGND.t2175 VGND.t650 2068.18
R13608 VGND.t2935 VGND.t1365 2068.18
R13609 VGND.t2192 VGND.t2935 2068.18
R13610 VGND.t2943 VGND.t2192 2068.18
R13611 VGND.t2977 VGND.t2943 2068.18
R13612 VGND.t4185 VGND.t2977 2068.18
R13613 VGND.t416 VGND.t4185 2068.18
R13614 VGND.t2681 VGND.t416 2068.18
R13615 VGND.t2883 VGND.t3054 2068.18
R13616 VGND.t3668 VGND.t2883 2068.18
R13617 VGND.t2208 VGND.t3668 2068.18
R13618 VGND.t640 VGND.t2208 2068.18
R13619 VGND.t1314 VGND.t640 2068.18
R13620 VGND.t2187 VGND.t1314 2068.18
R13621 VGND.t3839 VGND.t2187 2068.18
R13622 VGND.t4407 VGND.t4832 2068.18
R13623 VGND.t408 VGND.t4407 2068.18
R13624 VGND.t1398 VGND.t408 2068.18
R13625 VGND.t619 VGND.t1398 2068.18
R13626 VGND.t2281 VGND.t619 2068.18
R13627 VGND.t3343 VGND.t2281 2068.18
R13628 VGND.t766 VGND.t3343 2068.18
R13629 VGND.t3009 VGND.t1574 2068.18
R13630 VGND.t2751 VGND.t3009 2068.18
R13631 VGND.t2683 VGND.t2751 2068.18
R13632 VGND.t4204 VGND.t2683 2068.18
R13633 VGND.t1260 VGND.t4204 2068.18
R13634 VGND.t5798 VGND.t1260 2068.18
R13635 VGND.t4712 VGND.t5798 2068.18
R13636 VGND.t782 VGND.t2126 2068.18
R13637 VGND.t4899 VGND.t782 2068.18
R13638 VGND.t2924 VGND.t4899 2068.18
R13639 VGND.t1839 VGND.t2924 2068.18
R13640 VGND.t1214 VGND.t1839 2068.18
R13641 VGND.t1764 VGND.t1214 2068.18
R13642 VGND.t2006 VGND.t1764 2068.18
R13643 VGND.t1877 VGND.t905 2068.18
R13644 VGND.t2080 VGND.t1877 2068.18
R13645 VGND.t1497 VGND.t2080 2068.18
R13646 VGND.t3511 VGND.t1497 2068.18
R13647 VGND.t1937 VGND.t3511 2068.18
R13648 VGND.t1169 VGND.t1937 2068.18
R13649 VGND.t3970 VGND.t1169 2068.18
R13650 VGND.t4127 VGND.t1030 2068.18
R13651 VGND.t5213 VGND.t4127 2068.18
R13652 VGND.t3076 VGND.t5213 2068.18
R13653 VGND.t557 VGND.t3076 2068.18
R13654 VGND.t1088 VGND.t557 2068.18
R13655 VGND.t2711 VGND.t1088 2068.18
R13656 VGND.t622 VGND.t2711 2068.18
R13657 VGND.t5498 VGND.t2194 2068.18
R13658 VGND.t1722 VGND.t5498 2068.18
R13659 VGND.t354 VGND.t1722 2068.18
R13660 VGND.t489 VGND.t354 2068.18
R13661 VGND.t2849 VGND.t489 2068.18
R13662 VGND.t3507 VGND.t2849 2068.18
R13663 VGND.t61 VGND.t3507 2068.18
R13664 VGND.t3542 VGND.t3444 2068.18
R13665 VGND.t854 VGND.t3542 2068.18
R13666 VGND.t2461 VGND.t854 2068.18
R13667 VGND.t742 VGND.t2461 2068.18
R13668 VGND.t4153 VGND.t742 2068.18
R13669 VGND.t2106 VGND.t4153 2068.18
R13670 VGND.t3193 VGND.t2106 2068.18
R13671 VGND.t997 VGND.t1641 2068.18
R13672 VGND.t646 VGND.t997 2068.18
R13673 VGND.t2586 VGND.t646 2068.18
R13674 VGND.t3845 VGND.t2586 2068.18
R13675 VGND.t3339 VGND.t3845 2068.18
R13676 VGND.t1799 VGND.t3339 2068.18
R13677 VGND.t3890 VGND.t1799 2068.18
R13678 VGND.t5639 VGND.t3031 2068.18
R13679 VGND.t2269 VGND.t5639 2068.18
R13680 VGND.t4074 VGND.t2269 2068.18
R13681 VGND.t607 VGND.t4074 2068.18
R13682 VGND.t652 VGND.t607 2068.18
R13683 VGND.t2439 VGND.t652 2068.18
R13684 VGND.t475 VGND.t2439 2068.18
R13685 VGND.t4080 VGND.t730 2068.18
R13686 VGND.t362 VGND.t4080 2068.18
R13687 VGND.t2086 VGND.t362 2068.18
R13688 VGND.t3755 VGND.t2086 2068.18
R13689 VGND.t0 VGND.t3755 2068.18
R13690 VGND.t3062 VGND.t0 2068.18
R13691 VGND.t352 VGND.t3062 2068.18
R13692 VGND.t1130 VGND.t1375 2068.18
R13693 VGND.t2713 VGND.t1130 2068.18
R13694 VGND.t762 VGND.t2713 2068.18
R13695 VGND.t448 VGND.t762 2068.18
R13696 VGND.t2142 VGND.t448 2068.18
R13697 VGND.t2772 VGND.t2142 2068.18
R13698 VGND.t1406 VGND.t2772 2068.18
R13699 VGND.t4938 VGND.t2540 2068.18
R13700 VGND.t3294 VGND.t4938 2068.18
R13701 VGND.t4200 VGND.t3294 2068.18
R13702 VGND.t371 VGND.t4200 2068.18
R13703 VGND.t3499 VGND.t371 2068.18
R13704 VGND.t501 VGND.t3499 2068.18
R13705 VGND.t320 VGND.t501 2068.18
R13706 VGND.t3501 VGND.t483 2068.18
R13707 VGND.t2767 VGND.t3501 2068.18
R13708 VGND.t458 VGND.t2767 2068.18
R13709 VGND.t1823 VGND.t458 2068.18
R13710 VGND.t1904 VGND.t1823 2068.18
R13711 VGND.t3672 VGND.t1904 2068.18
R13712 VGND.t686 VGND.t3672 2068.18
R13713 VGND.t491 VGND.t2617 2068.18
R13714 VGND.t2341 VGND.t2065 2068.18
R13715 VGND.t907 VGND.t5240 2068.18
R13716 VGND.t1991 VGND.t907 2068.18
R13717 VGND.t1408 VGND.t2023 2068.18
R13718 VGND.t2124 VGND.t1408 2068.18
R13719 VGND.t2491 VGND.t2124 2068.18
R13720 VGND.t2294 VGND.t2491 2068.18
R13721 VGND.t4828 VGND.t2294 2068.18
R13722 VGND.t660 VGND.t4828 2068.18
R13723 VGND.t2217 VGND.t660 2068.18
R13724 VGND.t1329 VGND.t2074 2068.18
R13725 VGND.t551 VGND.t1090 2068.18
R13726 VGND.t360 VGND.t1483 2068.18
R13727 VGND.t2367 VGND.t523 2068.18
R13728 VGND.t523 VGND.t402 2068.18
R13729 VGND.t402 VGND.t1165 2068.18
R13730 VGND.t1165 VGND.t719 2068.18
R13731 VGND.t719 VGND.t2743 2068.18
R13732 VGND.t2743 VGND.t1249 2068.18
R13733 VGND.t1249 VGND.t1879 2068.18
R13734 VGND.t3411 VGND.t1613 2068.18
R13735 VGND.t1613 VGND.t2363 2068.18
R13736 VGND.t2363 VGND.t1561 2068.18
R13737 VGND.t1561 VGND.t2300 2068.18
R13738 VGND.t2300 VGND.t5062 2068.18
R13739 VGND.t5062 VGND.t2343 2068.18
R13740 VGND.t2343 VGND.t3977 2068.18
R13741 VGND.t3300 VGND.t2903 2068.18
R13742 VGND.t49 VGND.t2739 2068.18
R13743 VGND.t2842 VGND.t49 2068.18
R13744 VGND.t1022 VGND.t2842 2068.18
R13745 VGND.t4739 VGND.t1022 2068.18
R13746 VGND.t5150 VGND.t4739 2068.18
R13747 VGND.t3592 VGND.t1883 2068.18
R13748 VGND.t3353 VGND.t3592 2068.18
R13749 VGND.t2582 VGND.t3353 2068.18
R13750 VGND.t5180 VGND.t2582 2068.18
R13751 VGND.t77 VGND.t5180 2068.18
R13752 VGND.t3866 VGND.t77 2068.18
R13753 VGND.t1036 VGND.t3866 2068.18
R13754 VGND.t3078 VGND.t4879 2068.18
R13755 VGND.t4879 VGND.t577 2068.18
R13756 VGND.t577 VGND.t863 2068.18
R13757 VGND.t863 VGND.t5020 2068.18
R13758 VGND.t5020 VGND.t3309 2068.18
R13759 VGND.t3309 VGND.t3288 2068.18
R13760 VGND.t3288 VGND.t2232 2068.18
R13761 VGND.t1321 VGND.t1116 2068.18
R13762 VGND.t1116 VGND.t2594 2068.18
R13763 VGND.t2594 VGND.t5924 2068.18
R13764 VGND.t5924 VGND.t4034 2068.18
R13765 VGND.t4034 VGND.t2947 2068.18
R13766 VGND.t2947 VGND.t2699 2068.18
R13767 VGND.t2699 VGND.t3471 2068.18
R13768 VGND.t4290 VGND.t3385 2068.18
R13769 VGND.t3385 VGND.t2471 2068.18
R13770 VGND.t2471 VGND.t833 2068.18
R13771 VGND.t833 VGND.t966 2068.18
R13772 VGND.t966 VGND.t3096 2068.18
R13773 VGND.t3096 VGND.t4604 2068.18
R13774 VGND.t4604 VGND.t2795 2068.18
R13775 VGND.t5658 VGND.t3523 2068.18
R13776 VGND.t1793 VGND.t5658 2068.18
R13777 VGND.t2640 VGND.t1793 2068.18
R13778 VGND.t464 VGND.t2640 2068.18
R13779 VGND.t670 VGND.t464 2068.18
R13780 VGND.t2960 VGND.t670 2068.18
R13781 VGND.t4548 VGND.t2960 2068.18
R13782 VGND.t1762 VGND.t1643 2068.18
R13783 VGND.t1643 VGND.t553 2068.18
R13784 VGND.t553 VGND.t701 2068.18
R13785 VGND.t701 VGND.t3919 2068.18
R13786 VGND.t3919 VGND.t3718 2068.18
R13787 VGND.t3718 VGND.t964 2068.18
R13788 VGND.t2035 VGND.t3648 2068.18
R13789 VGND.t976 VGND.t5441 2068.18
R13790 VGND.t4883 VGND.t976 2068.18
R13791 VGND.t4983 VGND.t4883 2068.18
R13792 VGND.t2770 VGND.t4983 2068.18
R13793 VGND.t5649 VGND.t2770 2068.18
R13794 VGND.t1939 VGND.t5649 2068.18
R13795 VGND.t1400 VGND.t1939 2068.18
R13796 VGND.t404 VGND.t1132 2068.18
R13797 VGND.t3546 VGND.t404 2068.18
R13798 VGND.t4094 VGND.t3546 2068.18
R13799 VGND.t2877 VGND.t4094 2068.18
R13800 VGND.t1430 VGND.t2877 2068.18
R13801 VGND.t4110 VGND.t1430 2068.18
R13802 VGND.t909 VGND.t4110 2068.18
R13803 VGND.t879 VGND.t968 2068.18
R13804 VGND.t726 VGND.t5023 2068.18
R13805 VGND.t3616 VGND.t726 2068.18
R13806 VGND.t5478 VGND.t3616 2068.18
R13807 VGND.t3066 VGND.t1065 2068.18
R13808 VGND.t2159 VGND.t3066 2068.18
R13809 VGND.t446 VGND.t2159 2068.18
R13810 VGND.t960 VGND.t446 2068.18
R13811 VGND.t1371 VGND.t960 2068.18
R13812 VGND.t375 VGND.t1371 2068.18
R13813 VGND.t3181 VGND.t4302 2068.18
R13814 VGND.t4302 VGND.t2555 2068.18
R13815 VGND.t2555 VGND.t2879 2068.18
R13816 VGND.t2879 VGND.t373 2068.18
R13817 VGND.t373 VGND.t2351 2068.18
R13818 VGND.t1814 VGND.t5038 2068.18
R13819 VGND.t5038 VGND.t1524 2068.18
R13820 VGND.t1524 VGND.t2927 2068.18
R13821 VGND.t2927 VGND.t1339 2068.18
R13822 VGND.t1339 VGND.t2339 2068.18
R13823 VGND.t2339 VGND.t3037 2068.18
R13824 VGND.t3037 VGND.t3217 2068.18
R13825 VGND.t5512 VGND.t2333 2068.18
R13826 VGND.t2333 VGND.t1287 2068.18
R13827 VGND.t1287 VGND.t3703 2068.18
R13828 VGND.t3703 VGND.t2557 2068.18
R13829 VGND.t2557 VGND.t3897 2068.18
R13830 VGND.t3897 VGND.t1154 2068.18
R13831 VGND.t1154 VGND.t339 2068.18
R13832 VGND.t579 VGND.t3571 2068.18
R13833 VGND.t3571 VGND.t2950 2068.18
R13834 VGND.t2950 VGND.t1732 2068.18
R13835 VGND.t1732 VGND.t341 2068.18
R13836 VGND.t341 VGND.t381 2068.18
R13837 VGND.t381 VGND.t3044 2068.18
R13838 VGND.t3044 VGND.t613 2068.18
R13839 VGND.t2729 VGND.t4008 2068.18
R13840 VGND.t2707 VGND.t2729 2068.18
R13841 VGND.t2896 VGND.t2707 2068.18
R13842 VGND.t1049 VGND.t2896 2068.18
R13843 VGND.t1708 VGND.t1049 2068.18
R13844 VGND.t1908 VGND.t1708 2068.18
R13845 VGND.t4372 VGND.t1908 2068.18
R13846 VGND.t369 VGND.t3540 2068.18
R13847 VGND.t3540 VGND.t2025 2068.18
R13848 VGND.t2025 VGND.t1005 2068.18
R13849 VGND.t1005 VGND.t2200 2068.18
R13850 VGND.t2200 VGND.t3165 2068.18
R13851 VGND.t3165 VGND.t1041 2068.18
R13852 VGND.t1041 VGND.t1578 2068.18
R13853 VGND.t1053 VGND.t564 2068.18
R13854 VGND.t980 VGND.t1053 2068.18
R13855 VGND.t1204 VGND.t980 2068.18
R13856 VGND.t956 VGND.t1685 2068.18
R13857 VGND.t1685 VGND.t805 2068.18
R13858 VGND.t805 VGND.t4327 2068.18
R13859 VGND.t4327 VGND.t1024 2068.18
R13860 VGND.t1024 VGND.t751 2068.18
R13861 VGND.t751 VGND.t444 2068.18
R13862 VGND.t444 VGND.t848 2068.18
R13863 VGND.t440 VGND.t3458 2068.18
R13864 VGND.t1867 VGND.t3321 2068.18
R13865 VGND.t1354 VGND.t1867 2068.18
R13866 VGND.t2092 VGND.t1354 2068.18
R13867 VGND.t2969 VGND.t2092 2068.18
R13868 VGND.t638 VGND.t5429 2068.18
R13869 VGND.t5429 VGND.t3517 2068.18
R13870 VGND.t3517 VGND.t923 2068.18
R13871 VGND.t923 VGND.t1176 2068.18
R13872 VGND.t1176 VGND.t809 2068.18
R13873 VGND.t809 VGND.t1971 2068.18
R13874 VGND.t1971 VGND.t4639 2068.18
R13875 VGND.t892 VGND.t4131 2068.18
R13876 VGND.t666 VGND.t892 2068.18
R13877 VGND.t735 VGND.t666 2068.18
R13878 VGND.t1624 VGND.t735 2068.18
R13879 VGND.t367 VGND.t1624 2068.18
R13880 VGND.t2229 VGND.t3177 2068.18
R13881 VGND.t3177 VGND.t2161 2068.18
R13882 VGND.t2161 VGND.t3126 2068.18
R13883 VGND.t3126 VGND.t595 2068.18
R13884 VGND.t595 VGND.t3052 2068.18
R13885 VGND.t3052 VGND.t3947 2068.18
R13886 VGND.t3947 VGND.t1977 2068.18
R13887 VGND.t3163 VGND.t1943 2068.18
R13888 VGND.t1120 VGND.t3163 2068.18
R13889 VGND.t1128 VGND.t1120 2068.18
R13890 VGND.t2493 VGND.t1128 2068.18
R13891 VGND.t1136 VGND.t2493 2068.18
R13892 VGND.t67 VGND.t1136 2068.18
R13893 VGND.t1272 VGND.t3297 2068.18
R13894 VGND.t3297 VGND.t1887 2068.18
R13895 VGND.t1887 VGND.t1206 2068.18
R13896 VGND.t1206 VGND.t377 2068.18
R13897 VGND.t377 VGND.t513 2068.18
R13898 VGND.t513 VGND.t895 2068.18
R13899 VGND.t895 VGND.t549 2068.18
R13900 VGND.t2952 VGND.t4129 2068.18
R13901 VGND.t1171 VGND.t2952 2068.18
R13902 VGND.t1220 VGND.t1171 2068.18
R13903 VGND.t347 VGND.t1220 2068.18
R13904 VGND.t1224 VGND.t347 2068.18
R13905 VGND.t1292 VGND.t1224 2068.18
R13906 VGND.t2922 VGND.t1292 2068.18
R13907 VGND.t3216 VGND.t6307 1869.67
R13908 VGND.t2337 VGND.t1827 1791.19
R13909 VGND.t2459 VGND 1754.26
R13910 VGND.t4532 VGND.t3536 1735.8
R13911 VGND.t2954 VGND.t6670 1735.8
R13912 VGND.n654 VGND.t3124 1717.33
R13913 VGND.t4819 VGND.t2992 1708.1
R13914 VGND.t3640 VGND.t4970 1708.1
R13915 VGND.t2377 VGND.t3943 1708.1
R13916 VGND.t6069 VGND.t6067 1698.86
R13917 VGND.t173 VGND.t171 1698.86
R13918 VGND.t6129 VGND.t6132 1698.86
R13919 VGND.t153 VGND.t151 1698.86
R13920 VGND.n3699 VGND.n41 1655.57
R13921 VGND.n565 VGND.t1807 1569.6
R13922 VGND.t3705 VGND.t1379 1551.14
R13923 VGND.t3882 VGND.t4022 1551.14
R13924 VGND.t1835 VGND.t3004 1551.14
R13925 VGND.t593 VGND.t5395 1551.14
R13926 VGND.t3305 VGND.t5951 1551.14
R13927 VGND.n1124 VGND.t5868 1551.14
R13928 VGND.t4164 VGND.t5125 1551.14
R13929 VGND.t2660 VGND.t3493 1551.14
R13930 VGND.t6092 VGND.t5439 1551.14
R13931 VGND.t1900 VGND.t4339 1551.14
R13932 VGND.t4555 VGND.t333 1551.14
R13933 VGND.t2292 VGND.t5568 1551.14
R13934 VGND.t2405 VGND.t2265 1551.14
R13935 VGND.t710 VGND.t3796 1551.14
R13936 VGND.t697 VGND.t311 1551.14
R13937 VGND.t1440 VGND.t6186 1551.14
R13938 VGND.t1738 VGND.t2309 1551.14
R13939 VGND.t4796 VGND.t5336 1551.14
R13940 VGND.t1997 VGND.t4447 1551.14
R13941 VGND.t5635 VGND.t4743 1551.14
R13942 VGND.t962 VGND.t1980 1551.14
R13943 VGND.t4786 VGND.t2774 1551.14
R13944 VGND.t4491 VGND.t4174 1551.14
R13945 VGND.t2805 VGND.t4380 1551.14
R13946 VGND.t3460 VGND.t1567 1551.14
R13947 VGND.t4552 VGND.t1633 1551.14
R13948 VGND.t3094 VGND.t4090 1551.14
R13949 VGND.t5447 VGND.t807 1551.14
R13950 VGND.t412 VGND.t1308 1551.14
R13951 VGND.t3763 VGND.t1923 1551.14
R13952 VGND.t6078 VGND.t5161 1551.14
R13953 VGND.t4233 VGND.t3359 1551.14
R13954 VGND.t1341 VGND.t2318 1551.14
R13955 VGND.t1247 VGND.t2584 1551.14
R13956 VGND.t3351 VGND.t1570 1551.14
R13957 VGND.t3907 VGND.t2679 1551.14
R13958 VGND.t1635 VGND.t4944 1551.14
R13959 VGND.t3307 VGND.t5137 1551.14
R13960 VGND.t4749 VGND.t5900 1551.14
R13961 VGND.t2069 VGND.t1864 1551.14
R13962 VGND.t5544 VGND.t690 1551.14
R13963 VGND.t4478 VGND.t3534 1551.14
R13964 VGND.t597 VGND.t1528 1551.14
R13965 VGND.t629 VGND.t5841 1551.14
R13966 VGND.t1989 VGND.t875 1551.14
R13967 VGND.t3396 VGND.t1969 1551.14
R13968 VGND.t2409 VGND.t4872 1551.14
R13969 VGND.t1892 VGND.t654 1551.14
R13970 VGND.t3239 VGND.n467 1551.14
R13971 VGND.t562 VGND.t1526 1551.14
R13972 VGND.t728 VGND.t1202 1551.14
R13973 VGND.t5847 VGND.t2500 1551.14
R13974 VGND.t3560 VGND.t5320 1551.14
R13975 VGND.t1436 VGND.t4100 1551.14
R13976 VGND.t3818 VGND.t1359 1551.14
R13977 VGND.t1416 VGND.t764 1551.14
R13978 VGND.t4426 VGND.t5109 1551.14
R13979 VGND.t5127 VGND.t4137 1551.14
R13980 VGND.t2933 VGND.t1724 1551.14
R13981 VGND.t5970 VGND.t3098 1551.14
R13982 VGND.t1278 VGND.t4140 1551.14
R13983 VGND.t2050 VGND.t4217 1551.14
R13984 VGND.t2263 VGND.t5653 1551.14
R13985 VGND.t850 VGND.t5093 1551.14
R13986 VGND.t318 VGND.t2542 1551.14
R13987 VGND.t4696 VGND.t793 1551.14
R13988 VGND.t4507 VGND.t5668 1551.14
R13989 VGND.t3273 VGND.t1414 1551.14
R13990 VGND.t5680 VGND.t5521 1551.14
R13991 VGND.t2565 VGND.t795 1551.14
R13992 VGND.t503 VGND.t4765 1551.14
R13993 VGND.t5313 VGND.t4987 1551.14
R13994 VGND.t1396 VGND.t1019 1551.14
R13995 VGND.t1714 VGND.t3806 1551.14
R13996 VGND.t5357 VGND.t1580 1551.14
R13997 VGND.t1549 VGND.t1559 1551.14
R13998 VGND.t1444 VGND.t6750 1551.14
R13999 VGND.t1489 VGND.t4621 1551.14
R14000 VGND.t4794 VGND.t601 1551.14
R14001 VGND.t2204 VGND.t5433 1551.14
R14002 VGND.t1885 VGND.t4350 1551.14
R14003 VGND.t6076 VGND.t5875 1551.14
R14004 VGND.t4329 VGND.t4188 1551.14
R14005 VGND.t4431 VGND.t2078 1551.14
R14006 VGND.t2151 VGND.t2110 1551.14
R14007 VGND.t1003 VGND.t4876 1551.14
R14008 VGND.t414 VGND.t1493 1551.14
R14009 VGND.t4155 VGND.t5540 1551.14
R14010 VGND.t2311 VGND.t1963 1551.14
R14011 VGND.t3577 VGND.t1438 1551.14
R14012 VGND.t1951 VGND.t4612 1551.14
R14013 VGND.t2574 VGND.t1392 1551.14
R14014 VGND.t2255 VGND.t6796 1551.14
R14015 VGND.t3626 VGND.t852 1551.14
R14016 VGND.t3742 VGND.t5549 1551.14
R14017 VGND.t1647 VGND.t2185 1551.14
R14018 VGND.t1495 VGND.t3573 1551.14
R14019 VGND.t4914 VGND.t2003 1551.14
R14020 VGND.t3720 VGND.t799 1551.14
R14021 VGND.t1871 VGND.t1941 1551.14
R14022 VGND.t1805 VGND.n2495 1551.14
R14023 VGND.n2497 VGND.t497 1551.14
R14024 VGND.n405 VGND.t2887 1551.14
R14025 VGND.t4036 VGND.t5825 1551.14
R14026 VGND.t2029 VGND.t1466 1551.14
R14027 VGND.t978 VGND.t1356 1551.14
R14028 VGND.t1174 VGND.t5647 1551.14
R14029 VGND.t2755 VGND.t3798 1551.14
R14030 VGND.t1043 VGND.t1957 1551.14
R14031 VGND.t2323 VGND.t5326 1551.14
R14032 VGND.t495 VGND.t4271 1551.14
R14033 VGND.t3714 VGND.t1530 1551.14
R14034 VGND.t784 VGND.t5380 1551.14
R14035 VGND.t1833 VGND.t4792 1551.14
R14036 VGND.t2090 VGND.t2365 1551.14
R14037 VGND.t4397 VGND.t4088 1551.14
R14038 VGND.t1337 VGND.t5346 1551.14
R14039 VGND.t3993 VGND.t5888 1551.14
R14040 VGND.t4658 VGND.t3843 1551.14
R14041 VGND.t5186 VGND.t3119 1551.14
R14042 VGND.t4449 VGND.t1343 1551.14
R14043 VGND.t2885 VGND.t3438 1551.14
R14044 VGND.t5838 VGND.t3550 1551.14
R14045 VGND.t3854 VGND.t1818 1551.14
R14046 VGND.t5246 VGND.t3035 1551.14
R14047 VGND.t4891 VGND.t4770 1551.14
R14048 VGND.t5959 VGND.t672 1551.14
R14049 VGND.t51 VGND.t2325 1551.14
R14050 VGND.t3585 VGND.t5717 1551.14
R14051 VGND.t1576 VGND.t533 1551.14
R14052 VGND.t2349 VGND.t4378 1551.14
R14053 VGND.t5407 VGND.t668 1551.14
R14054 VGND.t1657 VGND.t4725 1551.14
R14055 VGND.t1222 VGND.t3205 1551.14
R14056 VGND.t4356 VGND.t5800 1551.14
R14057 VGND.t1210 VGND.t3011 1551.14
R14058 VGND.t1331 VGND.t5103 1551.14
R14059 VGND.t2789 VGND.t3856 1551.14
R14060 VGND.t5468 VGND.t4474 1551.14
R14061 VGND.t3230 VGND.t1797 1551.14
R14062 VGND.t813 VGND.t5738 1551.14
R14063 VGND.t5003 VGND.t958 1551.14
R14064 VGND.t2898 VGND.t1276 1551.14
R14065 VGND.t6767 VGND.t4850 1551.14
R14066 VGND.t379 VGND.t2719 1551.14
R14067 VGND.t4779 VGND.t4249 1551.14
R14068 VGND.t4211 VGND.t1107 1551.14
R14069 VGND.t2122 VGND.t3646 1551.14
R14070 VGND.t2286 VGND.t4927 1551.14
R14071 VGND.t4952 VGND.t2215 1551.14
R14072 VGND.t4215 VGND.t2656 1551.14
R14073 VGND.t5064 VGND.t6802 1551.14
R14074 VGND.t1281 VGND.t3183 1551.14
R14075 VGND.t1987 VGND.t4304 1551.14
R14076 VGND.t4714 VGND.t4482 1551.14
R14077 VGND.t1477 VGND.t2147 1551.14
R14078 VGND.t434 VGND.t2303 1551.14
R14079 VGND.t3927 VGND.t1676 1551.14
R14080 VGND.t4830 VGND.t1597 1551.14
R14081 VGND.t5201 VGND.t1196 1551.14
R14082 VGND.t5574 VGND.t791 1551.14
R14083 VGND.t5861 VGND.t4487 1551.14
R14084 VGND.t1432 VGND.t1915 1551.14
R14085 VGND.t3792 VGND.t3383 1551.14
R14086 VGND.t5269 VGND.t1843 1551.14
R14087 VGND.t5318 VGND.t4502 1551.14
R14088 VGND.t5730 VGND.t5452 1551.14
R14089 VGND.t1599 VGND.t1710 1551.14
R14090 VGND.t65 VGND.t3142 1551.14
R14091 VGND.t6040 VGND.t5977 1551.14
R14092 VGND.t6173 VGND.t499 1551.14
R14093 VGND.t1627 VGND.t1781 1551.14
R14094 VGND.t1156 VGND.t4756 1551.14
R14095 VGND.t4881 VGND.t1367 1551.14
R14096 VGND.t4607 VGND.t1198 1551.14
R14097 VGND.t2650 VGND.t4190 1551.14
R14098 VGND.t4610 VGND.t2622 1551.14
R14099 VGND.t712 VGND.t2824 1551.14
R14100 VGND.t4202 VGND.t3664 1551.14
R14101 VGND.t2307 VGND.t2347 1551.14
R14102 VGND.t5930 VGND.t2369 1551.14
R14103 VGND.t745 VGND.t1534 1551.14
R14104 VGND.t1081 VGND.t3744 1551.14
R14105 VGND.t4822 VGND.t4665 1551.14
R14106 VGND.t5917 VGND.t2402 1551.14
R14107 VGND.t4614 VGND.t4716 1551.14
R14108 VGND.t4142 VGND.t3870 1551.14
R14109 VGND.t1692 VGND.t2104 1551.14
R14110 VGND.t3258 VGND.t732 1551.14
R14111 VGND.t5771 VGND.t5851 1551.14
R14112 VGND.t5602 VGND.t4907 1551.14
R14113 VGND.t3473 VGND.t2576 1551.14
R14114 VGND.t3442 VGND.t1369 1551.14
R14115 VGND.t4444 VGND.t1200 1551.14
R14116 VGND.t4300 VGND.t4194 1551.14
R14117 VGND.t5947 VGND.t3092 1551.14
R14118 VGND.t3656 VGND.t3260 1551.14
R14119 VGND.t3868 VGND.t3115 1551.14
R14120 VGND.t3666 VGND.t418 1551.14
R14121 VGND.t2988 VGND.t2526 1551.14
R14122 VGND.t3525 VGND.t6018 1551.14
R14123 VGND.t5956 VGND.t3394 1551.14
R14124 VGND.t4461 VGND.t4183 1551.14
R14125 VGND.t3997 VGND.t674 1551.14
R14126 VGND.t1760 VGND.t1756 1551.14
R14127 VGND.t5553 VGND.t4463 1551.14
R14128 VGND.t3587 VGND.t5397 1551.14
R14129 VGND.t6034 VGND.t2847 1551.14
R14130 VGND.t3925 VGND.t5481 1551.14
R14131 VGND.t970 VGND.t2223 1551.14
R14132 VGND.t3696 VGND.t2183 1551.14
R14133 VGND.t5949 VGND.t4352 1551.14
R14134 VGND.t566 VGND.t2741 1551.14
R14135 VGND.t1743 VGND.t1298 1551.14
R14136 VGND.t4367 VGND.t3877 1551.14
R14137 VGND.t3090 VGND.t5926 1551.14
R14138 VGND.t3538 VGND.t2061 1551.14
R14139 VGND.t5975 VGND.t2892 1551.14
R14140 VGND.t2871 VGND.t4806 1551.14
R14141 VGND.t3604 VGND.t1789 1551.14
R14142 VGND.t1791 VGND.t4166 1551.14
R14143 VGND.t3694 VGND.t2134 1551.14
R14144 VGND.t5199 VGND.t4267 1551.14
R14145 VGND.t5920 VGND.t4024 1551.14
R14146 VGND.t4901 VGND.t4568 1551.14
R14147 VGND.t995 VGND.t1706 1551.14
R14148 VGND.t4440 VGND.t3406 1551.14
R14149 VGND.t1716 VGND.t2422 1551.14
R14150 VGND.t2749 VGND.t3774 1551.14
R14151 VGND.t2426 VGND.t5525 1551.14
R14152 VGND.t1726 VGND.t972 1551.14
R14153 VGND.t2345 VGND.t4451 1551.14
R14154 VGND.t974 VGND.t3345 1551.14
R14155 VGND.t564 VGND.n2969 1551.14
R14156 VGND.n2971 VGND.t956 1551.14
R14157 VGND.n376 VGND.t2753 1551.14
R14158 VGND.t3321 VGND.n3075 1551.14
R14159 VGND.n3077 VGND.t638 1551.14
R14160 VGND.n368 VGND.t1085 1551.14
R14161 VGND.t4131 VGND.n3181 1551.14
R14162 VGND.n3183 VGND.t2229 1551.14
R14163 VGND.n361 VGND.t3228 1551.14
R14164 VGND.t1943 VGND.n3311 1551.14
R14165 VGND.t4129 VGND.n8 1551.14
R14166 VGND.n1725 VGND.t5632 1532.67
R14167 VGND.t2144 VGND.t3850 1532.67
R14168 VGND VGND.t186 1532.67
R14169 VGND.t6101 VGND.t5694 1514.2
R14170 VGND.t680 VGND.t6473 1514.2
R14171 VGND.t6312 VGND.t856 1514.2
R14172 VGND.t3130 VGND 1504.97
R14173 VGND.t1847 VGND 1504.97
R14174 VGND VGND.t2084 1504.97
R14175 VGND.t3746 VGND 1504.97
R14176 VGND.t5227 VGND 1504.97
R14177 VGND VGND.t1194 1504.97
R14178 VGND.t2277 VGND 1504.97
R14179 VGND.t1243 VGND 1504.97
R14180 VGND VGND.t537 1504.97
R14181 VGND.t605 VGND 1504.97
R14182 VGND.t4495 VGND 1504.97
R14183 VGND VGND.t1631 1504.97
R14184 VGND.t5734 VGND.t428 1495.74
R14185 VGND.t298 VGND.t1455 1495.74
R14186 VGND.t5416 VGND.t990 1495.74
R14187 VGND.t2573 VGND.t2764 1495.74
R14188 VGND.t929 VGND.t5843 1440.34
R14189 VGND.t6349 VGND 1421.88
R14190 VGND.t6569 VGND 1421.88
R14191 VGND.t204 VGND 1421.88
R14192 VGND.t6392 VGND.t6594 1403.41
R14193 VGND.t6719 VGND.t195 1403.41
R14194 VGND.t5365 VGND.t6571 1403.41
R14195 VGND.t6516 VGND.t3245 1403.41
R14196 VGND.t4160 VGND.t718 1403.41
R14197 VGND VGND.t3268 1403.41
R14198 VGND.t1688 VGND.t6468 1398.79
R14199 VGND VGND.t2171 1394.18
R14200 VGND VGND.t4348 1394.18
R14201 VGND.t5592 VGND 1366.48
R14202 VGND.t4016 VGND 1366.48
R14203 VGND VGND.t4227 1348.01
R14204 VGND.t555 VGND 1348.01
R14205 VGND.t4343 VGND 1348.01
R14206 VGND.t1365 VGND 1348.01
R14207 VGND.t3962 VGND 1348.01
R14208 VGND.t3054 VGND 1348.01
R14209 VGND VGND.t4471 1348.01
R14210 VGND.t4832 VGND 1348.01
R14211 VGND.t4752 VGND 1348.01
R14212 VGND.t1574 VGND 1348.01
R14213 VGND.t1694 VGND 1348.01
R14214 VGND.t2126 VGND 1348.01
R14215 VGND.t2487 VGND 1348.01
R14216 VGND.t905 VGND 1348.01
R14217 VGND.t2528 VGND 1348.01
R14218 VGND.t1030 VGND 1348.01
R14219 VGND.t1667 VGND 1348.01
R14220 VGND.t2194 VGND 1348.01
R14221 VGND.t3319 VGND 1348.01
R14222 VGND.t3444 VGND 1348.01
R14223 VGND.t2284 VGND 1348.01
R14224 VGND.t1641 VGND 1348.01
R14225 VGND.t5820 VGND 1348.01
R14226 VGND.t3031 VGND 1348.01
R14227 VGND.t5338 VGND 1348.01
R14228 VGND.t730 VGND 1348.01
R14229 VGND VGND.t5353 1348.01
R14230 VGND.t1375 VGND 1348.01
R14231 VGND.t5117 VGND 1348.01
R14232 VGND.t2540 VGND 1348.01
R14233 VGND.t483 VGND 1348.01
R14234 VGND VGND.t491 1348.01
R14235 VGND.t3567 VGND.t5461 1348.01
R14236 VGND VGND.n891 1348.01
R14237 VGND VGND.t3548 1348.01
R14238 VGND.t2371 VGND 1348.01
R14239 VGND.t1736 VGND 1348.01
R14240 VGND.t2654 VGND 1348.01
R14241 VGND.t350 VGND 1348.01
R14242 VGND.t3303 VGND 1348.01
R14243 VGND VGND.t2341 1348.01
R14244 VGND.t5091 VGND.t6274 1348.01
R14245 VGND.t493 VGND 1348.01
R14246 VGND.t1795 VGND 1348.01
R14247 VGND.t5240 VGND 1348.01
R14248 VGND.t3211 VGND 1348.01
R14249 VGND.t2023 VGND 1348.01
R14250 VGND.t5025 VGND 1348.01
R14251 VGND.t5908 VGND.t5682 1348.01
R14252 VGND.t3237 VGND 1348.01
R14253 VGND.t2074 VGND 1348.01
R14254 VGND.t1090 VGND 1348.01
R14255 VGND.t1306 VGND 1348.01
R14256 VGND.t3558 VGND 1348.01
R14257 VGND VGND.t2367 1348.01
R14258 VGND.n665 VGND.t3575 1348.01
R14259 VGND.t5362 VGND 1348.01
R14260 VGND.t4512 VGND 1348.01
R14261 VGND.t5324 VGND 1348.01
R14262 VGND VGND.t3411 1348.01
R14263 VGND VGND.t1001 1348.01
R14264 VGND.t2638 VGND 1348.01
R14265 VGND.t2890 VGND 1348.01
R14266 VGND VGND.t823 1348.01
R14267 VGND.t1593 VGND 1348.01
R14268 VGND.t2903 VGND 1348.01
R14269 VGND.t2739 VGND 1348.01
R14270 VGND.t3232 VGND 1348.01
R14271 VGND.t1883 VGND 1348.01
R14272 VGND VGND.t3078 1348.01
R14273 VGND VGND.t1321 1348.01
R14274 VGND VGND.t4290 1348.01
R14275 VGND.t3523 VGND 1348.01
R14276 VGND VGND.t1973 1348.01
R14277 VGND VGND.t3967 1348.01
R14278 VGND VGND.t1762 1348.01
R14279 VGND.t3648 VGND 1348.01
R14280 VGND.t2067 VGND 1348.01
R14281 VGND.n529 VGND.t4225 1348.01
R14282 VGND.t5441 VGND 1348.01
R14283 VGND.t617 VGND 1348.01
R14284 VGND.t2289 VGND 1348.01
R14285 VGND.t3024 VGND 1348.01
R14286 VGND.t5624 VGND 1348.01
R14287 VGND.t4480 VGND 1348.01
R14288 VGND VGND.t991 1348.01
R14289 VGND VGND.t4219 1348.01
R14290 VGND VGND.t3621 1348.01
R14291 VGND VGND.t1093 1348.01
R14292 VGND VGND.t3670 1348.01
R14293 VGND.t5359 VGND 1348.01
R14294 VGND.t1132 VGND 1348.01
R14295 VGND.t3921 VGND 1348.01
R14296 VGND.t968 VGND 1348.01
R14297 VGND.t5023 VGND 1348.01
R14298 VGND.t1065 VGND 1348.01
R14299 VGND VGND.t3181 1348.01
R14300 VGND VGND.t3170 1348.01
R14301 VGND VGND.t3712 1348.01
R14302 VGND.t3019 VGND 1348.01
R14303 VGND.t5829 VGND 1348.01
R14304 VGND.t2189 VGND 1348.01
R14305 VGND VGND.t1814 1348.01
R14306 VGND VGND.t5512 1348.01
R14307 VGND.t1565 VGND 1348.01
R14308 VGND.t4698 VGND 1348.01
R14309 VGND VGND.t4133 1348.01
R14310 VGND VGND.t2165 1348.01
R14311 VGND.t487 VGND 1348.01
R14312 VGND VGND.t579 1348.01
R14313 VGND.t4041 VGND 1348.01
R14314 VGND.t4008 VGND 1348.01
R14315 VGND.t2094 VGND 1348.01
R14316 VGND VGND.t369 1348.01
R14317 VGND.t4660 VGND 1348.01
R14318 VGND VGND.t2149 1348.01
R14319 VGND VGND.t440 1348.01
R14320 VGND VGND.t3161 1348.01
R14321 VGND VGND.t1272 1348.01
R14322 VGND VGND.n380 1335.62
R14323 VGND.n3019 VGND 1335.62
R14324 VGND.n3020 VGND 1335.62
R14325 VGND.n3021 VGND 1335.62
R14326 VGND VGND.n372 1335.62
R14327 VGND.n3124 VGND 1335.62
R14328 VGND.n3125 VGND 1335.62
R14329 VGND.n3126 VGND 1335.62
R14330 VGND VGND.n365 1335.62
R14331 VGND.n3230 VGND 1335.62
R14332 VGND.n3231 VGND 1335.62
R14333 VGND.n3232 VGND 1335.62
R14334 VGND.n3233 VGND 1335.62
R14335 VGND.n3234 VGND 1335.62
R14336 VGND VGND.n1 1335.62
R14337 VGND.n3776 VGND 1335.62
R14338 VGND.n3777 VGND 1335.62
R14339 VGND.t4809 VGND.t2971 1329.55
R14340 VGND.t4929 VGND.t6036 1311.08
R14341 VGND VGND.t6693 1311.08
R14342 VGND VGND.t6144 1311.08
R14343 VGND.t456 VGND.t197 1311.08
R14344 VGND.t6191 VGND 1311.08
R14345 VGND.n732 VGND.t1589 1292.61
R14346 VGND.t3046 VGND.t5173 1292.61
R14347 VGND.t6140 VGND.t6134 1290.2
R14348 VGND.t2602 VGND.t117 1255.68
R14349 VGND VGND.t4524 1241.83
R14350 VGND.n899 VGND 1237.22
R14351 VGND.t4296 VGND.t5292 1237.22
R14352 VGND.t3760 VGND 1237.22
R14353 VGND.t1622 VGND 1237.22
R14354 VGND VGND.t4824 1237.22
R14355 VGND VGND.t1151 1237.22
R14356 VGND VGND.n943 1237.22
R14357 VGND.t327 VGND.t585 1237.22
R14358 VGND.t5156 VGND 1237.22
R14359 VGND.t4994 VGND.t5746 1237.22
R14360 VGND.t2765 VGND.t1776 1218.75
R14361 VGND.t5588 VGND.t14 1218.75
R14362 VGND.t144 VGND.t2986 1218.75
R14363 VGND.t6327 VGND.t385 1218.75
R14364 VGND.n783 VGND.t264 1218.75
R14365 VGND.t5562 VGND.t6683 1218.75
R14366 VGND.t92 VGND.t4510 1218.75
R14367 VGND.t5299 VGND.t4654 1218.75
R14368 VGND VGND.t6002 1218.75
R14369 VGND.t6631 VGND.t572 1218.75
R14370 VGND.t6677 VGND.t3375 1200.28
R14371 VGND.t873 VGND.t6008 1200.28
R14372 VGND.t6428 VGND.t3894 1200.28
R14373 VGND VGND.t3767 1200.28
R14374 VGND.t1253 VGND.t831 1200.28
R14375 VGND.t2331 VGND.t3467 1200.28
R14376 VGND.t5506 VGND.t169 1200.28
R14377 VGND.t4863 VGND.n522 1200.28
R14378 VGND VGND.t3784 1195.67
R14379 VGND.t694 VGND.t4117 1191.05
R14380 VGND.t676 VGND.t4277 1191.05
R14381 VGND.t3347 VGND.t1557 1191.05
R14382 VGND.t4694 VGND.t3989 1191.05
R14383 VGND.t3650 VGND.t507 1191.05
R14384 VGND.t5163 VGND.t4955 1191.05
R14385 VGND.t5508 VGND.t2475 1191.05
R14386 VGND.t772 VGND.t4256 1191.05
R14387 VGND.t4489 VGND.t5721 1191.05
R14388 VGND.t6748 VGND.t4974 1191.05
R14389 VGND.t5743 VGND.t5225 1191.05
R14390 VGND.t2038 VGND.t2249 1191.05
R14391 VGND.t6466 VGND.t3728 1181.82
R14392 VGND VGND.t6644 1181.82
R14393 VGND.t2012 VGND 1157.53
R14394 VGND.t5551 VGND 1157.53
R14395 VGND.t2931 VGND 1157.53
R14396 VGND VGND.t1163 1157.53
R14397 VGND VGND.t2808 1157.53
R14398 VGND.t4258 VGND 1157.53
R14399 VGND.t1967 VGND 1157.53
R14400 VGND VGND.t3999 1157.53
R14401 VGND VGND.t625 1157.53
R14402 VGND.t2040 VGND 1157.53
R14403 VGND.t3110 VGND 1157.53
R14404 VGND VGND.t3349 1157.53
R14405 VGND VGND.t2832 1157.53
R14406 VGND VGND.t5189 1157.53
R14407 VGND VGND.t5519 1157.53
R14408 VGND.t5966 VGND 1157.53
R14409 VGND.t5340 VGND 1157.53
R14410 VGND VGND.t2202 1157.53
R14411 VGND VGND.t1442 1157.53
R14412 VGND.t1345 VGND 1126.42
R14413 VGND.t2807 VGND 1126.42
R14414 VGND.t2448 VGND 1126.42
R14415 VGND.t1373 VGND.t452 1126.42
R14416 VGND.t2810 VGND.t2219 1126.42
R14417 VGND.t2136 VGND.t3064 1126.42
R14418 VGND.t1906 VGND.t1264 1126.42
R14419 VGND VGND.t6691 1107.95
R14420 VGND.t1516 VGND.t164 1107.95
R14421 VGND.t6235 VGND.t4978 1104.99
R14422 VGND VGND.t5399 1103.34
R14423 VGND VGND.t3002 1089.49
R14424 VGND.t2797 VGND.t858 1089.49
R14425 VGND VGND.t5600 1084.87
R14426 VGND.t1180 VGND.t6394 1071.02
R14427 VGND.t1849 VGND.t1847 1061.79
R14428 VGND.t2084 VGND.t2082 1061.79
R14429 VGND.t2171 VGND.t2169 1061.79
R14430 VGND.t881 VGND.t883 1061.79
R14431 VGND.t5231 VGND.t5227 1061.79
R14432 VGND.t1194 VGND.t1192 1061.79
R14433 VGND.t4682 VGND.t4684 1061.79
R14434 VGND.t1772 VGND.t1774 1061.79
R14435 VGND.t5982 VGND.t5984 1061.79
R14436 VGND.t541 VGND.t539 1061.79
R14437 VGND.t1239 VGND.t1241 1061.79
R14438 VGND.t1509 VGND.t1507 1061.79
R14439 VGND.t5896 VGND.t5898 1061.79
R14440 VGND.t1653 VGND.t1655 1061.79
R14441 VGND.t537 VGND.t535 1061.79
R14442 VGND.t2251 VGND.t2253 1061.79
R14443 VGND.t4692 VGND.t4690 1061.79
R14444 VGND.t1422 VGND.t1420 1061.79
R14445 VGND.t5302 VGND.t5300 1061.79
R14446 VGND.t5494 VGND.t5492 1061.79
R14447 VGND.t603 VGND.t605 1061.79
R14448 VGND.t944 VGND.t942 1061.79
R14449 VGND.t1428 VGND.t1426 1061.79
R14450 VGND.t1649 VGND.t1651 1061.79
R14451 VGND.t2514 VGND.t4527 1055.25
R14452 VGND.t1563 VGND.t927 1052.56
R14453 VGND.t1976 VGND.t4996 1047.94
R14454 VGND.t3147 VGND.t305 1038.71
R14455 VGND.t1749 VGND.t5906 1034.09
R14456 VGND.t3048 VGND.t1749 1034.09
R14457 VGND.n273 VGND.t299 1034.09
R14458 VGND.t1837 VGND.t6555 1034.09
R14459 VGND.t3332 VGND.t3327 1034.09
R14460 VGND.t4720 VGND.t3642 1034.09
R14461 VGND.t1811 VGND.t5916 1034.09
R14462 VGND.t2047 VGND.t3355 1034.09
R14463 VGND.t2522 VGND.t2524 1034.09
R14464 VGND.t16 VGND.t1013 1034.09
R14465 VGND.t3802 VGND.t644 1034.09
R14466 VGND.t788 VGND 1034.09
R14467 VGND.t4030 VGND.t4026 1034.09
R14468 VGND.t6237 VGND.t3446 1034.09
R14469 VGND.t6244 VGND.t5702 1034.09
R14470 VGND.t5459 VGND.t5178 1034.09
R14471 VGND.t5288 VGND.t2384 1034.09
R14472 VGND.t4686 VGND.t5531 1034.09
R14473 VGND.t1346 VGND.t1348 1034.09
R14474 VGND.t1352 VGND.t1350 1034.09
R14475 VGND.t4834 VGND.t3608 1034.09
R14476 VGND.t6329 VGND.t1862 1034.09
R14477 VGND.t3688 VGND.t6426 1034.09
R14478 VGND.t3674 VGND.t4538 1034.09
R14479 VGND.t3589 VGND.t3676 1034.09
R14480 VGND.t4422 VGND.t5760 1034.09
R14481 VGND.t3117 VGND.t229 1034.09
R14482 VGND.t6355 VGND.t225 1034.09
R14483 VGND.t1931 VGND.t6492 1034.09
R14484 VGND.t3430 VGND.t3424 1034.09
R14485 VGND.t5184 VGND 1034.09
R14486 VGND.t399 VGND.t6539 1034.09
R14487 VGND.t387 VGND.t391 1034.09
R14488 VGND.t6112 VGND.t5415 1034.09
R14489 VGND.t6113 VGND.t6216 1034.09
R14490 VGND.t6700 VGND.t2464 1034.09
R14491 VGND.t2590 VGND.t2592 1034.09
R14492 VGND.t6686 VGND.t725 1034.09
R14493 VGND.t4561 VGND.t6687 1034.09
R14494 VGND.t6460 VGND.t6096 1034.09
R14495 VGND.t6281 VGND.t6279 1034.09
R14496 VGND.t6289 VGND.t6285 1034.09
R14497 VGND.t6285 VGND.t6283 1034.09
R14498 VGND.t18 VGND.t2353 1034.09
R14499 VGND.t2353 VGND.t6276 1034.09
R14500 VGND.t5656 VGND.t569 1034.09
R14501 VGND.t5890 VGND.t5690 1034.09
R14502 VGND.t4688 VGND.t473 1034.09
R14503 VGND.t6385 VGND.t2815 1034.09
R14504 VGND.t5682 VGND.t6786 1034.09
R14505 VGND.t4004 VGND.t1503 1034.09
R14506 VGND.t3155 VGND.t4758 1034.09
R14507 VGND.t186 VGND.t1186 1034.09
R14508 VGND.t1186 VGND.t183 1034.09
R14509 VGND.t183 VGND.t130 1034.09
R14510 VGND.t270 VGND.t272 1034.09
R14511 VGND.t284 VGND.t288 1034.09
R14512 VGND.t3419 VGND.t3418 1034.09
R14513 VGND.t1588 VGND.t5445 1034.09
R14514 VGND.t1813 VGND.t529 1034.09
R14515 VGND.t6049 VGND.t2972 1034.09
R14516 VGND.t6222 VGND.t6115 1034.09
R14517 VGND.t6383 VGND.t2857 1034.09
R14518 VGND.t3247 VGND.t2260 1034.09
R14519 VGND.t3771 VGND.t3247 1034.09
R14520 VGND.t2813 VGND.t3199 1034.09
R14521 VGND.t4325 VGND.t219 1034.09
R14522 VGND.t2685 VGND.t2398 1034.09
R14523 VGND.t2691 VGND.t3594 1034.09
R14524 VGND.t1557 VGND.t5688 1034.09
R14525 VGND.t6309 VGND.t6450 1034.09
R14526 VGND.t23 VGND.t3828 1034.09
R14527 VGND.t4992 VGND.t915 1034.09
R14528 VGND.t260 VGND.t258 1034.09
R14529 VGND.t244 VGND.t246 1034.09
R14530 VGND.t2918 VGND.t4957 1034.09
R14531 VGND.t4256 VGND.t2912 1034.09
R14532 VGND.t303 VGND.t6336 1034.09
R14533 VGND.t3080 VGND.t5243 1034.09
R14534 VGND.t1933 VGND.t6148 1034.09
R14535 VGND.t210 VGND.t6123 1034.09
R14536 VGND.t3017 VGND.t1310 1034.09
R14537 VGND.t1325 VGND.t5872 1034.09
R14538 VGND.t4384 VGND.t5991 1034.09
R14539 VGND.t5723 VGND.t3776 1034.09
R14540 VGND.t5159 VGND.t2840 1034.09
R14541 VGND.t2840 VGND.t755 1034.09
R14542 VGND.t755 VGND.t6181 1034.09
R14543 VGND.t6181 VGND.t5342 1034.09
R14544 VGND.t5342 VGND.t2717 1034.09
R14545 VGND.t2717 VGND.t2909 1034.09
R14546 VGND.t2909 VGND.t4811 1034.09
R14547 VGND.t4811 VGND.t2693 1034.09
R14548 VGND.t2693 VGND.t4370 1034.09
R14549 VGND.t4370 VGND.t5845 1034.09
R14550 VGND.t5845 VGND.t3489 1034.09
R14551 VGND.t3489 VGND.t5248 1034.09
R14552 VGND.t160 VGND.t6367 1034.09
R14553 VGND.t6369 VGND.t6733 1034.09
R14554 VGND.t162 VGND.t4864 1034.09
R14555 VGND.t1522 VGND.t1296 1034.09
R14556 VGND.t1845 VGND.t5558 1034.09
R14557 VGND.t4147 VGND.t1845 1034.09
R14558 VGND.t5107 VGND.t4147 1034.09
R14559 VGND.t2390 VGND.t5107 1034.09
R14560 VGND.t3903 VGND.t2390 1034.09
R14561 VGND.t2211 VGND.t3903 1034.09
R14562 VGND.t4247 VGND.t2211 1034.09
R14563 VGND.t5431 VGND.t4247 1034.09
R14564 VGND.t5485 VGND.t5431 1034.09
R14565 VGND.t5751 VGND.t5485 1034.09
R14566 VGND.t703 VGND.t5751 1034.09
R14567 VGND.t1912 VGND.t703 1034.09
R14568 VGND.t5457 VGND.t1912 1034.09
R14569 VGND.t4393 VGND.t5457 1034.09
R14570 VGND.t2670 VGND.t4393 1034.09
R14571 VGND.t4817 VGND.t1208 1034.09
R14572 VGND.t1208 VGND.t3463 1034.09
R14573 VGND.t3463 VGND.t4705 1034.09
R14574 VGND.t4705 VGND.t4557 1034.09
R14575 VGND.t4557 VGND.t4574 1034.09
R14576 VGND.t4574 VGND.t3875 1034.09
R14577 VGND.t3875 VGND.t2298 1034.09
R14578 VGND.t2298 VGND.t1540 1034.09
R14579 VGND.t1540 VGND.t5348 1034.09
R14580 VGND.t5348 VGND.t5167 1034.09
R14581 VGND.t5167 VGND.t2396 1034.09
R14582 VGND.t2396 VGND.t2612 1034.09
R14583 VGND.t2612 VGND.t59 1034.09
R14584 VGND.t59 VGND.t2335 1034.09
R14585 VGND.t2335 VGND.t521 1034.09
R14586 VGND.t5105 VGND.n2629 1034.09
R14587 VGND.t5449 VGND.n2630 1034.09
R14588 VGND.t6815 VGND.n2631 1034.09
R14589 VGND.t3637 VGND.n2632 1034.09
R14590 VGND.t2453 VGND.t2227 1034.09
R14591 VGND.t6363 VGND.t40 1034.09
R14592 VGND.t5067 VGND.n2095 1034.09
R14593 VGND.n2096 VGND.t2538 1034.09
R14594 VGND.t5014 VGND.t3275 1034.09
R14595 VGND.t5389 VGND.t5001 1034.09
R14596 VGND.t5001 VGND.t5372 1034.09
R14597 VGND.t5372 VGND.t1851 1034.09
R14598 VGND.t1851 VGND.t3256 1034.09
R14599 VGND.t3256 VGND.t1758 1034.09
R14600 VGND.t1758 VGND.t2327 1034.09
R14601 VGND.t185 VGND.t3632 1034.09
R14602 VGND.t1975 VGND.t1007 1034.09
R14603 VGND.t3041 VGND.t202 1034.09
R14604 VGND.t4540 VGND.t4520 1034.09
R14605 VGND.t2072 VGND.t5753 1034.09
R14606 VGND.t6089 VGND.t2072 1034.09
R14607 VGND.t817 VGND.t684 1034.09
R14608 VGND.t5203 VGND.t817 1034.09
R14609 VGND.t365 VGND.t5203 1034.09
R14610 VGND.t821 VGND.t365 1034.09
R14611 VGND.t4800 VGND.t821 1034.09
R14612 VGND.t845 VGND.t4800 1034.09
R14613 VGND.t838 VGND.t4045 1034.09
R14614 VGND.t753 VGND.t2532 1034.09
R14615 VGND.t57 VGND.t753 1034.09
R14616 VGND.t3505 VGND.t57 1034.09
R14617 VGND.t3234 VGND.t3505 1034.09
R14618 VGND.t4465 VGND.t4207 1034.09
R14619 VGND.t4207 VGND.t4285 1034.09
R14620 VGND.t4285 VGND.t1232 1034.09
R14621 VGND.t1232 VGND.t3758 1034.09
R14622 VGND.t3758 VGND.t1167 1034.09
R14623 VGND.t1167 VGND.t4804 1034.09
R14624 VGND.t4804 VGND.t4298 1034.09
R14625 VGND.t4298 VGND.t531 1034.09
R14626 VGND.t4499 VGND.t1690 1034.09
R14627 VGND.t1953 VGND.t4499 1034.09
R14628 VGND.t3598 VGND.t1953 1034.09
R14629 VGND.t4634 VGND.t3598 1034.09
R14630 VGND.t5670 VGND.t4634 1034.09
R14631 VGND.t3006 VGND.t5670 1034.09
R14632 VGND.t2561 VGND.t3006 1034.09
R14633 VGND.t4761 VGND.t2561 1034.09
R14634 VGND.t5405 VGND.t4761 1034.09
R14635 VGND.t3734 VGND.t5405 1034.09
R14636 VGND.t2801 VGND.t3734 1034.09
R14637 VGND.t3864 VGND.t2801 1034.09
R14638 VGND.t2614 VGND.t3864 1034.09
R14639 VGND.t4484 VGND.t2614 1034.09
R14640 VGND.t6055 VGND.t4484 1034.09
R14641 VGND.t3088 VGND.t1134 1034.09
R14642 VGND.t4625 VGND.t5628 1034.09
R14643 VGND.t481 VGND.t4625 1034.09
R14644 VGND.t1752 VGND.t309 1034.09
R14645 VGND.t309 VGND.t2163 1034.09
R14646 VGND.t2163 VGND.t843 1034.09
R14647 VGND.t843 VGND.t4852 1034.09
R14648 VGND.t4852 VGND.t3816 1034.09
R14649 VGND.t3816 VGND.t1896 1034.09
R14650 VGND.t1896 VGND.t6081 1034.09
R14651 VGND.t6081 VGND.t1051 1034.09
R14652 VGND.t1051 VGND.t2668 1034.09
R14653 VGND.t2668 VGND.t2844 1034.09
R14654 VGND.t1983 VGND.t1890 1034.09
R14655 VGND.t633 VGND.t1983 1034.09
R14656 VGND.t2662 VGND.t633 1034.09
R14657 VGND.t383 VGND.t2662 1034.09
R14658 VGND.t815 VGND.t383 1034.09
R14659 VGND.t4619 VGND.t815 1034.09
R14660 VGND.t3872 VGND.t4619 1034.09
R14661 VGND.t1487 VGND.t3872 1034.09
R14662 VGND.t4745 VGND.t1487 1034.09
R14663 VGND.t1720 VGND.t4745 1034.09
R14664 VGND.t714 VGND.t1720 1034.09
R14665 VGND.t4598 VGND.t714 1034.09
R14666 VGND.t2000 VGND.t4598 1034.09
R14667 VGND.t5072 VGND.t2000 1034.09
R14668 VGND.t6176 VGND.t5072 1034.09
R14669 VGND.t1118 VGND.t3337 1034.09
R14670 VGND.t1779 VGND.t4802 1034.09
R14671 VGND.t4802 VGND.t5831 1034.09
R14672 VGND.t5831 VGND.t5962 1034.09
R14673 VGND.t5962 VGND.t5538 1034.09
R14674 VGND.t5538 VGND.t2551 1034.09
R14675 VGND.t2551 VGND.t6053 1034.09
R14676 VGND.t6053 VGND.t3619 1034.09
R14677 VGND.t3619 VGND.t5726 1034.09
R14678 VGND.t5726 VGND.t6061 1034.09
R14679 VGND.t6061 VGND.t1226 1034.09
R14680 VGND.t1226 VGND.t2443 1034.09
R14681 VGND.t2443 VGND.t1712 1034.09
R14682 VGND.t3532 VGND.t5774 1034.09
R14683 VGND.t3810 VGND.t3532 1034.09
R14684 VGND.t1816 VGND.t3810 1034.09
R14685 VGND.t5273 VGND.t1816 1034.09
R14686 VGND.t5266 VGND.t5273 1034.09
R14687 VGND.t1615 VGND.t5266 1034.09
R14688 VGND.t3140 VGND.t1615 1034.09
R14689 VGND.t4947 VGND.t3140 1034.09
R14690 VGND.t3724 VGND.t4947 1034.09
R14691 VGND.t4059 VGND.t3724 1034.09
R14692 VGND.t6772 VGND.t4059 1034.09
R14693 VGND.t6006 VGND.t6772 1034.09
R14694 VGND.t2830 VGND.t6006 1034.09
R14695 VGND.t3082 VGND.t2830 1034.09
R14696 VGND.t3552 VGND.t3082 1034.09
R14697 VGND.t933 VGND.t4591 1034.09
R14698 VGND.t5070 VGND.t933 1034.09
R14699 VGND.t1730 VGND.t5070 1034.09
R14700 VGND.t1474 VGND.t1730 1034.09
R14701 VGND.t4172 VGND.t1474 1034.09
R14702 VGND.t4209 VGND.t4172 1034.09
R14703 VGND.t2851 VGND.t4209 1034.09
R14704 VGND.t3364 VGND.t2851 1034.09
R14705 VGND.t840 VGND.t3364 1034.09
R14706 VGND.t4772 VGND.t840 1034.09
R14707 VGND.t1158 VGND.t4772 1034.09
R14708 VGND.t4181 VGND.t1158 1034.09
R14709 VGND.t4623 VGND.t4181 1034.09
R14710 VGND.t1728 VGND.t4623 1034.09
R14711 VGND.t4354 VGND.t5311 1034.09
R14712 VGND.t5922 VGND.t4354 1034.09
R14713 VGND.t797 VGND.t5922 1034.09
R14714 VGND.t2496 VGND.t797 1034.09
R14715 VGND.t422 VGND.t2496 1034.09
R14716 VGND.t4576 VGND.t422 1034.09
R14717 VGND.t4243 VGND.t4576 1034.09
R14718 VGND.t5637 VGND.t4243 1034.09
R14719 VGND.t2648 VGND.t5637 1034.09
R14720 VGND.t5853 VGND.t2648 1034.09
R14721 VGND.t3544 VGND.t5853 1034.09
R14722 VGND.t631 VGND.t3544 1034.09
R14723 VGND.t4923 VGND.t631 1034.09
R14724 VGND.t3195 VGND.t4923 1034.09
R14725 VGND.t5788 VGND.t6588 1020.24
R14726 VGND.t5796 VGND.t6586 1020.24
R14727 VGND.t3056 VGND.t6236 1018.96
R14728 VGND VGND.t2520 1015.62
R14729 VGND.t4071 VGND.t4294 1015.62
R14730 VGND.t6204 VGND.t6777 1015.62
R14731 VGND.t3748 VGND 1015.62
R14732 VGND.t5827 VGND.t3941 1015.62
R14733 VGND.t3428 VGND.t4055 1015.62
R14734 VGND VGND.t6229 1015.62
R14735 VGND VGND.t954 1015.62
R14736 VGND.t927 VGND.t861 1015.62
R14737 VGND.t2467 VGND 1015.62
R14738 VGND.t32 VGND 1015.62
R14739 VGND.t6706 VGND 1015.62
R14740 VGND.t5910 VGND 1015.62
R14741 VGND.t4361 VGND 1015.62
R14742 VGND.t1034 VGND 1015.62
R14743 VGND.t2512 VGND 1015.62
R14744 VGND.t6520 VGND 1015.62
R14745 VGND.t6543 VGND 1015.62
R14746 VGND.t986 VGND.t21 1015.62
R14747 VGND.t5660 VGND 1015.62
R14748 VGND.t4919 VGND 1015.62
R14749 VGND.t2537 VGND 1015.62
R14750 VGND VGND.t6580 1015.62
R14751 VGND VGND.t2451 1015.62
R14752 VGND VGND.t4312 1015.62
R14753 VGND.t786 VGND.n1483 1011.01
R14754 VGND.t4281 VGND.t331 1006.39
R14755 VGND.t6320 VGND.t6319 998.629
R14756 VGND.t3138 VGND.t776 997.159
R14757 VGND.t525 VGND.t988 997.159
R14758 VGND.t2464 VGND.t1770 997.159
R14759 VGND.t6689 VGND.t4391 997.159
R14760 VGND.t2157 VGND.t6263 997.159
R14761 VGND.t6287 VGND.t2155 997.159
R14762 VGND.t6497 VGND.t6663 997.159
R14763 VGND.t4845 VGND.t6610 997.159
R14764 VGND VGND.t4857 997.159
R14765 VGND.t2757 VGND.t3455 997.159
R14766 VGND VGND.t4981 997.159
R14767 VGND.t2504 VGND 997.159
R14768 VGND.t1532 VGND.t5523 992.543
R14769 VGND.t2359 VGND 987.927
R14770 VGND.t5421 VGND 987.927
R14771 VGND.t2782 VGND 987.927
R14772 VGND.t5027 VGND 987.927
R14773 VGND.t2994 VGND 987.927
R14774 VGND.t6616 VGND.t6620 983.298
R14775 VGND.t664 VGND 978.693
R14776 VGND VGND.t984 978.693
R14777 VGND.t3440 VGND.t1921 978.693
R14778 VGND.t3711 VGND.t2626 978.693
R14779 VGND.t2544 VGND.t16 974.077
R14780 VGND.t292 VGND.t2415 969.461
R14781 VGND.t5255 VGND.t4893 967.966
R14782 VGND.t3958 VGND.t4536 962.963
R14783 VGND.t4537 VGND.t3960 962.963
R14784 VGND.t6600 VGND.t4522 962.963
R14785 VGND.t6606 VGND.t4523 962.963
R14786 VGND.t6602 VGND.t2876 962.963
R14787 VGND.t6604 VGND.t2873 962.963
R14788 VGND.t6626 VGND.t4525 962.963
R14789 VGND.t6624 VGND.t4535 962.963
R14790 VGND.t2894 VGND.t6142 960.227
R14791 VGND.t6200 VGND.t2392 960.227
R14792 VGND.t682 VGND.t6359 960.227
R14793 VGND.t164 VGND.t3945 960.227
R14794 VGND.t6540 VGND.t3940 941.761
R14795 VGND.t835 VGND.t774 941.761
R14796 VGND.t6038 VGND.t6726 941.761
R14797 VGND.t6342 VGND.t6233 941.761
R14798 VGND.t5391 VGND.t2411 941.761
R14799 VGND.t425 VGND.t3837 941.761
R14800 VGND.t6024 VGND.t2058 941.761
R14801 VGND.t4673 VGND.t4073 941.761
R14802 VGND.t937 VGND.t6103 941.761
R14803 VGND.t6306 VGND.t6314 941.761
R14804 VGND.t6108 VGND.t6318 941.761
R14805 VGND.t663 VGND.t4788 924.163
R14806 VGND.t5277 VGND 923.295
R14807 VGND.t6526 VGND.t4643 923.295
R14808 VGND.t3145 VGND.t5299 923.295
R14809 VGND.t5368 VGND.t5085 923.295
R14810 VGND.t266 VGND.t6662 919.782
R14811 VGND.t1026 VGND.t6701 914.063
R14812 VGND VGND.t6721 904.831
R14813 VGND.t5297 VGND.t212 904.831
R14814 VGND.t890 VGND.t6549 904.831
R14815 VGND VGND.t3484 904.831
R14816 VGND VGND.t4121 904.831
R14817 VGND.t200 VGND 904.831
R14818 VGND.t6389 VGND.t6668 904.831
R14819 VGND.t4054 VGND.t6472 904.831
R14820 VGND.t1702 VGND.t5387 904.831
R14821 VGND.t5165 VGND 904.831
R14822 VGND VGND.t2473 904.831
R14823 VGND.t921 VGND.t2510 904.831
R14824 VGND.t2470 VGND.t4317 904.831
R14825 VGND.t1820 VGND.t6025 904.831
R14826 VGND.t5465 VGND.t6125 904.831
R14827 VGND.t1611 VGND.t5264 904.831
R14828 VGND VGND.t4972 904.831
R14829 VGND.t5741 VGND 904.831
R14830 VGND.n3669 VGND.n3480 895.597
R14831 VGND.n3669 VGND.n3481 895.597
R14832 VGND.n3669 VGND.n3482 895.597
R14833 VGND.n3669 VGND.n3668 895.597
R14834 VGND.n3673 VGND.n3669 895.597
R14835 VGND.n3559 VGND.n41 895.597
R14836 VGND.n3591 VGND.n41 895.597
R14837 VGND.n3623 VGND.n41 895.597
R14838 VGND.n3607 VGND.n41 895.597
R14839 VGND.n3575 VGND.n41 895.597
R14840 VGND.n3669 VGND.n42 895.597
R14841 VGND.n3358 VGND.n246 895.597
R14842 VGND.t2240 VGND.t6257 895.597
R14843 VGND.n3358 VGND.n270 895.597
R14844 VGND.n3359 VGND.n3358 895.597
R14845 VGND.n3358 VGND.n271 895.597
R14846 VGND.n3358 VGND.n272 895.597
R14847 VGND.t4855 VGND.t4648 895.597
R14848 VGND.n2207 VGND.n39 895.597
R14849 VGND.n2953 VGND.n388 895.597
R14850 VGND.n2953 VGND.n389 895.597
R14851 VGND.n2953 VGND.n400 895.597
R14852 VGND.n2954 VGND.n2953 895.597
R14853 VGND.n531 VGND.n39 895.597
R14854 VGND.n2332 VGND.n39 895.597
R14855 VGND.n2952 VGND.n401 895.597
R14856 VGND.n2952 VGND.n402 895.597
R14857 VGND.n2952 VGND.n403 895.597
R14858 VGND.n3358 VGND.n3357 895.597
R14859 VGND.t6551 VGND.t4671 890.981
R14860 VGND.t6678 VGND.t4848 886.365
R14861 VGND.t2778 VGND.t1145 886.365
R14862 VGND.t5916 VGND.t2130 886.365
R14863 VGND.t3530 VGND.t3341 886.365
R14864 VGND.t2631 VGND.t6443 886.365
R14865 VGND.t115 VGND.t6724 886.365
R14866 VGND.t3690 VGND.t3674 886.365
R14867 VGND.t6790 VGND.t6486 886.365
R14868 VGND.t106 VGND.t6488 886.365
R14869 VGND.t1603 VGND.t2019 886.365
R14870 VGND.t6614 VGND.t234 886.365
R14871 VGND.t3822 VGND.t4565 886.365
R14872 VGND.t85 VGND.t1126 886.365
R14873 VGND.t6371 VGND.t221 886.365
R14874 VGND.t1450 VGND.t5146 886.365
R14875 VGND.t3039 VGND.t6149 886.365
R14876 VGND.t2763 VGND.t3788 886.365
R14877 VGND.t740 VGND.t3315 886.365
R14878 VGND.t191 VGND.t6424 886.365
R14879 VGND VGND.t4264 886.365
R14880 VGND VGND.t1263 886.365
R14881 VGND.n1483 VGND.t233 881.747
R14882 VGND VGND.t4337 877.131
R14883 VGND.t4277 VGND.t432 877.131
R14884 VGND.t2703 VGND.t2905 877.131
R14885 VGND.t4836 VGND.t284 877.131
R14886 VGND VGND.t2956 877.131
R14887 VGND.t507 VGND.t5121 877.131
R14888 VGND.t917 VGND.t4162 877.131
R14889 VGND VGND.t3911 877.131
R14890 VGND.n1022 VGND.t511 877.131
R14891 VGND.t2120 VGND.t1100 867.899
R14892 VGND.t6254 VGND.t6477 867.899
R14893 VGND.t12 VGND.t6271 867.899
R14894 VGND.t3814 VGND.t5217 867.899
R14895 VGND.t3197 VGND.t5597 867.899
R14896 VGND.t5781 VGND 867.899
R14897 VGND.t3335 VGND.t6210 858.665
R14898 VGND.t6247 VGND.t2979 858.665
R14899 VGND.t5700 VGND.t2983 858.665
R14900 VGND.t5702 VGND.t2981 858.665
R14901 VGND.t4331 VGND.t5425 858.665
R14902 VGND.t4333 VGND.t5423 858.665
R14903 VGND.t2273 VGND.t1768 858.665
R14904 VGND.t2275 VGND.t1766 858.665
R14905 VGND.t3835 VGND.t5607 858.665
R14906 VGND.t3833 VGND.t5609 858.665
R14907 VGND.t3936 VGND.t2432 849.433
R14908 VGND.t3934 VGND.t1180 849.433
R14909 VGND.t5470 VGND.t2600 849.433
R14910 VGND.t6594 VGND.t2920 849.433
R14911 VGND VGND.n246 849.433
R14912 VGND.t3334 VGND.t6657 849.433
R14913 VGND.t6679 VGND.t780 849.433
R14914 VGND.t4119 VGND.t6348 849.433
R14915 VGND.t3168 VGND.t873 849.433
R14916 VGND.t2518 VGND.t2394 849.433
R14917 VGND.t3022 VGND.t5778 849.433
R14918 VGND.t1015 VGND.t19 849.433
R14919 VGND.t1947 VGND 849.433
R14920 VGND.t6250 VGND.t2244 849.433
R14921 VGND.t1776 VGND.t343 849.433
R14922 VGND.t6226 VGND.t4065 849.433
R14923 VGND.t4067 VGND.t6434 849.433
R14924 VGND.t5865 VGND.t144 849.433
R14925 VGND.t5016 VGND.t6327 849.433
R14926 VGND.t2246 VGND.t6259 849.433
R14927 VGND.t468 VGND.t3333 849.433
R14928 VGND.t163 VGND.t3432 849.433
R14929 VGND.t6534 VGND.t3480 849.433
R14930 VGND.n270 VGND 849.433
R14931 VGND.t112 VGND.t18 849.433
R14932 VGND.t3121 VGND.t6510 849.433
R14933 VGND.t2413 VGND.t5393 849.433
R14934 VGND.t6649 VGND.t4411 849.433
R14935 VGND.t6675 VGND.t4413 849.433
R14936 VGND.t6683 VGND.t599 849.433
R14937 VGND.n3359 VGND 849.433
R14938 VGND.t716 VGND.t189 849.433
R14939 VGND.t6511 VGND.t1188 849.433
R14940 VGND.t4964 VGND.t6547 849.433
R14941 VGND VGND.n271 849.433
R14942 VGND.t4847 VGND.t236 849.433
R14943 VGND.t6308 VGND.t937 849.433
R14944 VGND.t5344 VGND.t2271 849.433
R14945 VGND.t5783 VGND 849.433
R14946 VGND.t6323 VGND.t6110 849.433
R14947 VGND.t581 VGND.t92 849.433
R14948 VGND VGND.n272 849.433
R14949 VGND.t248 VGND.t6440 849.433
R14950 VGND.n944 VGND.t6146 849.433
R14951 VGND.t4647 VGND.t135 849.433
R14952 VGND.t232 VGND.t3252 849.433
R14953 VGND.t6518 VGND.t3249 849.433
R14954 VGND.t5364 VGND.t6158 849.433
R14955 VGND.t2569 VGND.t6579 849.433
R14956 VGND.n2207 VGND 849.433
R14957 VGND VGND.n388 849.433
R14958 VGND VGND.n389 849.433
R14959 VGND.n400 VGND 849.433
R14960 VGND.n2954 VGND 849.433
R14961 VGND.t6157 VGND.t6647 849.433
R14962 VGND.t2316 VGND.t6631 849.433
R14963 VGND.n531 VGND 849.433
R14964 VGND.n2332 VGND 849.433
R14965 VGND VGND.n404 849.433
R14966 VGND VGND.n401 849.433
R14967 VGND VGND.n402 849.433
R14968 VGND VGND.n403 849.433
R14969 VGND.t6149 VGND.t3200 849.433
R14970 VGND.t2449 VGND.t6301 849.433
R14971 VGND.n3357 VGND 849.433
R14972 VGND.t3632 VGND.t4505 849.433
R14973 VGND.t6022 VGND.t3770 849.433
R14974 VGND.t3265 VGND.t2382 835.582
R14975 VGND.t6567 VGND.t4905 835.582
R14976 VGND VGND.t1266 830.966
R14977 VGND VGND.t2267 830.966
R14978 VGND.t4544 VGND 830.966
R14979 VGND.t2535 VGND 830.966
R14980 VGND.t1456 VGND 830.966
R14981 VGND.t2646 VGND 830.966
R14982 VGND VGND.t6806 830.966
R14983 VGND VGND.t2008 830.966
R14984 VGND.t3654 VGND 830.966
R14985 VGND.t3414 VGND 830.966
R14986 VGND.t5282 VGND 830.966
R14987 VGND.t6782 VGND 830.966
R14988 VGND.t2088 VGND 830.966
R14989 VGND.t1659 VGND 830.966
R14990 VGND.t6755 VGND 830.966
R14991 VGND.t2225 VGND 830.966
R14992 VGND.t4261 VGND 830.966
R14993 VGND.t4826 VGND 830.966
R14994 VGND.t517 VGND 830.966
R14995 VGND.t2606 VGND 830.966
R14996 VGND.t1230 VGND 830.966
R14997 VGND.t3779 VGND 830.966
R14998 VGND.t1873 VGND 830.966
R14999 VGND.t73 VGND 830.966
R15000 VGND.t3450 VGND 830.966
R15001 VGND.t3581 VGND 830.966
R15002 VGND VGND.t4061 830.966
R15003 VGND VGND.t4178 830.966
R15004 VGND.t3686 VGND 830.966
R15005 VGND.t4213 VGND 830.966
R15006 VGND VGND.n282 830.966
R15007 VGND VGND.t2063 830.966
R15008 VGND VGND.t2735 830.966
R15009 VGND VGND.t5234 830.966
R15010 VGND VGND.n273 830.966
R15011 VGND.n152 VGND 830.966
R15012 VGND VGND.n1348 830.966
R15013 VGND.t4092 VGND 830.966
R15014 VGND.n1355 VGND 830.966
R15015 VGND VGND.n1360 830.966
R15016 VGND.t4032 VGND.t6778 830.966
R15017 VGND.t5698 VGND.t6441 830.966
R15018 VGND.n1371 VGND 830.966
R15019 VGND.t4376 VGND 830.966
R15020 VGND.t4319 VGND 830.966
R15021 VGND.t218 VGND.t4528 830.966
R15022 VGND.t5219 VGND.t143 830.966
R15023 VGND.t919 VGND.t4422 830.966
R15024 VGND.t5007 VGND.t3117 830.966
R15025 VGND.n1490 VGND.t890 830.966
R15026 VGND.t2196 VGND 830.966
R15027 VGND.t3495 VGND 830.966
R15028 VGND.n1499 VGND 830.966
R15029 VGND.t5415 VGND.t5350 830.966
R15030 VGND.t3760 VGND 830.966
R15031 VGND VGND.t2054 830.966
R15032 VGND VGND.n783 830.966
R15033 VGND.t3013 VGND 830.966
R15034 VGND.n1716 VGND 830.966
R15035 VGND.t3633 VGND 830.966
R15036 VGND.t345 VGND 830.966
R15037 VGND.n1721 VGND 830.966
R15038 VGND.t5835 VGND 830.966
R15039 VGND.t5316 VGND 830.966
R15040 VGND.t6682 VGND.t5307 830.966
R15041 VGND.t1333 VGND.t5253 830.966
R15042 VGND VGND.t5113 830.966
R15043 VGND VGND.t3974 830.966
R15044 VGND VGND.t2652 830.966
R15045 VGND.n1122 VGND 830.966
R15046 VGND VGND.n1122 830.966
R15047 VGND.t4252 VGND 830.966
R15048 VGND.t1319 VGND 830.966
R15049 VGND.n1123 VGND 830.966
R15050 VGND.t1151 VGND 830.966
R15051 VGND.t4870 VGND 830.966
R15052 VGND.t6528 VGND.t3151 830.966
R15053 VGND.t6532 VGND.t5385 830.966
R15054 VGND.n737 VGND.t2259 830.966
R15055 VGND.t155 VGND.t2489 830.966
R15056 VGND.t529 VGND.t4550 830.966
R15057 VGND.n1823 VGND 830.966
R15058 VGND.t1898 VGND 830.966
R15059 VGND.t2265 VGND 830.966
R15060 VGND.t3389 VGND 830.966
R15061 VGND.n655 VGND 830.966
R15062 VGND.n659 VGND 830.966
R15063 VGND.t1855 VGND 830.966
R15064 VGND.t2355 VGND 830.966
R15065 VGND.t4174 VGND 830.966
R15066 VGND.t1923 VGND 830.966
R15067 VGND.t4944 VGND 830.966
R15068 VGND.t2257 VGND 830.966
R15069 VGND VGND.t5294 830.966
R15070 VGND.t3707 VGND 830.966
R15071 VGND.t1184 VGND 830.966
R15072 VGND.t5822 VGND 830.966
R15073 VGND.n942 VGND 830.966
R15074 VGND.t6757 VGND 830.966
R15075 VGND.t4690 VGND.t2251 830.966
R15076 VGND.t2674 VGND 830.966
R15077 VGND.t125 VGND.n472 830.966
R15078 VGND.t2759 VGND.t4652 830.966
R15079 VGND.n478 VGND 830.966
R15080 VGND.t75 VGND 830.966
R15081 VGND.t3888 VGND 830.966
R15082 VGND VGND.t5938 830.966
R15083 VGND VGND.t3370 830.966
R15084 VGND VGND.t3491 830.966
R15085 VGND.t3701 VGND 830.966
R15086 VGND VGND.t4784 830.966
R15087 VGND VGND.t2636 830.966
R15088 VGND VGND.t3241 830.966
R15089 VGND.n466 VGND 830.966
R15090 VGND.t1917 VGND 830.966
R15091 VGND.t2580 VGND 830.966
R15092 VGND.t4170 VGND 830.966
R15093 VGND.t4641 VGND 830.966
R15094 VGND.t678 VGND.t6732 830.966
R15095 VGND.t591 VGND 830.966
R15096 VGND.t2042 VGND 830.966
R15097 VGND.t3243 VGND 830.966
R15098 VGND.t6051 VGND 830.966
R15099 VGND.t5677 VGND 830.966
R15100 VGND.t397 VGND 830.966
R15101 VGND.t5077 VGND 830.966
R15102 VGND.t5193 VGND 830.966
R15103 VGND VGND.t1831 830.966
R15104 VGND VGND.t6808 830.966
R15105 VGND VGND.t4580 830.966
R15106 VGND VGND.t1396 830.966
R15107 VGND VGND.t2204 830.966
R15108 VGND VGND.t414 830.966
R15109 VGND.t852 VGND 830.966
R15110 VGND.t4039 VGND 830.966
R15111 VGND.n2492 VGND 830.966
R15112 VGND.n2494 VGND 830.966
R15113 VGND.n2496 VGND 830.966
R15114 VGND VGND.n406 830.966
R15115 VGND VGND.t3172 830.966
R15116 VGND VGND.t2323 830.966
R15117 VGND.t5346 VGND 830.966
R15118 VGND.t1818 VGND 830.966
R15119 VGND.t4378 VGND 830.966
R15120 VGND.t547 VGND 830.966
R15121 VGND VGND.t3398 830.966
R15122 VGND.n2629 VGND 830.966
R15123 VGND.n2630 VGND 830.966
R15124 VGND.t2656 VGND 830.966
R15125 VGND.t3368 VGND 830.966
R15126 VGND.t5556 VGND 830.966
R15127 VGND.t1047 VGND 830.966
R15128 VGND.n2632 VGND 830.966
R15129 VGND.t4999 VGND 830.966
R15130 VGND.t2824 VGND 830.966
R15131 VGND.t5917 VGND 830.966
R15132 VGND VGND.t3473 830.966
R15133 VGND.t418 VGND 830.966
R15134 VGND.t1491 VGND 830.966
R15135 VGND.t1542 VGND 830.966
R15136 VGND.t4363 VGND 830.966
R15137 VGND VGND.n554 830.966
R15138 VGND VGND.t4108 830.966
R15139 VGND VGND.t4700 830.966
R15140 VGND.n2093 VGND 830.966
R15141 VGND.t2741 VGND 830.966
R15142 VGND.t3600 VGND 830.966
R15143 VGND.t2112 VGND 830.966
R15144 VGND.t1434 VGND 830.966
R15145 VGND.n2096 VGND 830.966
R15146 VGND VGND.t993 830.966
R15147 VGND.t5221 VGND 830.966
R15148 VGND.n1021 VGND 830.966
R15149 VGND.t4457 VGND.t315 830.966
R15150 VGND.t511 VGND.t2964 830.966
R15151 VGND VGND.n573 830.966
R15152 VGND VGND.n570 830.966
R15153 VGND.n2970 VGND 830.966
R15154 VGND VGND.n377 830.966
R15155 VGND.n3074 VGND 830.966
R15156 VGND.n3076 VGND 830.966
R15157 VGND VGND.n369 830.966
R15158 VGND.n3180 VGND 830.966
R15159 VGND.n3182 VGND 830.966
R15160 VGND VGND.n362 830.966
R15161 VGND.n3310 VGND 830.966
R15162 VGND.n3312 VGND 830.966
R15163 VGND VGND.n5 830.966
R15164 VGND.n7 VGND 830.966
R15165 VGND.t3751 VGND.t6515 830.966
R15166 VGND.t2329 VGND.t5427 826.35
R15167 VGND.t6253 VGND.t2243 820.303
R15168 VGND.t2245 VGND.t6256 820.303
R15169 VGND.t3935 VGND.t2428 812.5
R15170 VGND.t2437 VGND.t4731 812.5
R15171 VGND.t2503 VGND.t4231 812.5
R15172 VGND.t2505 VGND.t6584 812.5
R15173 VGND.t6653 VGND.n144 812.5
R15174 VGND.t4065 VGND.t6463 812.5
R15175 VGND.t5323 VGND.t3606 812.5
R15176 VGND.t3879 VGND.t5886 812.5
R15177 VGND.t3477 VGND.n776 812.5
R15178 VGND.t167 VGND.t6138 812.5
R15179 VGND.t911 VGND.t6135 812.5
R15180 VGND.t5376 VGND.t847 812.5
R15181 VGND.t238 VGND.t6608 812.5
R15182 VGND.t240 VGND.t6612 812.5
R15183 VGND.t1126 VGND.t82 812.5
R15184 VGND.t5087 VGND 812.5
R15185 VGND.t6639 VGND.t4965 807.885
R15186 VGND.t6232 VGND.t87 802.47
R15187 VGND.t252 VGND.t6723 802.47
R15188 VGND.t256 VGND.t9 802.47
R15189 VGND.t254 VGND.t8 802.47
R15190 VGND.t250 VGND.t6716 802.47
R15191 VGND.t5792 VGND.t5808 798.652
R15192 VGND.t1114 VGND.t4002 798.652
R15193 VGND.t769 VGND.t6703 798.652
R15194 VGND VGND.t2237 794.034
R15195 VGND.t1595 VGND.t3070 794.034
R15196 VGND.t2153 VGND.t6287 794.034
R15197 VGND.t26 VGND.t3956 794.034
R15198 VGND.t4933 VGND.t6387 794.034
R15199 VGND.t169 VGND.t1102 794.034
R15200 VGND.t6596 VGND.t2875 794.034
R15201 VGND.t6622 VGND.t4844 794.034
R15202 VGND.t4416 VGND.t126 794.034
R15203 VGND.t3455 VGND.t5244 794.034
R15204 VGND.t4940 VGND.t6127 794.034
R15205 VGND.t3583 VGND.t1514 794.034
R15206 VGND.t4977 VGND 784.636
R15207 VGND.t4159 VGND.t460 780.186
R15208 VGND.t6141 VGND.t6398 775.568
R15209 VGND.n278 VGND.t3521 775.568
R15210 VGND.t89 VGND.t3381 775.568
R15211 VGND.t90 VGND.t835 775.568
R15212 VGND.t4722 VGND.t6560 775.568
R15213 VGND.t4703 VGND.t6685 775.568
R15214 VGND.t1783 VGND.t3023 775.568
R15215 VGND.t5292 VGND.t4071 775.568
R15216 VGND.t789 VGND.t1412 775.568
R15217 VGND.t1949 VGND.t6739 775.568
R15218 VGND.t141 VGND.t5323 775.568
R15219 VGND.t801 VGND 775.568
R15220 VGND.t6324 VGND.t3879 775.568
R15221 VGND.t6298 VGND.t6352 775.568
R15222 VGND.t6295 VGND.t6342 775.568
R15223 VGND.t6338 VGND.t6293 775.568
R15224 VGND.t3509 VGND.n200 775.568
R15225 VGND.t6071 VGND.t925 775.568
R15226 VGND.n250 VGND.t1268 775.568
R15227 VGND VGND.t395 775.568
R15228 VGND.t6705 VGND.t4198 775.568
R15229 VGND.t1009 VGND.t6696 775.568
R15230 VGND.t3134 VGND.t5578 775.568
R15231 VGND.t30 VGND.t5817 775.568
R15232 VGND.t6027 VGND.t911 775.568
R15233 VGND.t5630 VGND 775.568
R15234 VGND.t3852 VGND 775.568
R15235 VGND.t5736 VGND.t4669 775.568
R15236 VGND.t847 VGND.t6680 775.568
R15237 VGND.t869 VGND.t4646 775.568
R15238 VGND.t1700 VGND.t1698 775.568
R15239 VGND.t1921 VGND.t6131 775.568
R15240 VGND.t452 VGND.t1587 775.568
R15241 VGND.t2644 VGND.t6119 775.568
R15242 VGND.t2219 VGND.t6050 775.568
R15243 VGND.t1395 VGND.t1955 775.568
R15244 VGND.t94 VGND.t5286 775.568
R15245 VGND.t3102 VGND.t6311 775.568
R15246 VGND.t2799 VGND.t3829 775.568
R15247 VGND.t1404 VGND.t4076 775.568
R15248 VGND.t4997 VGND.t6418 775.568
R15249 VGND.t2761 VGND.t125 775.568
R15250 VGND.t6713 VGND.t1064 775.568
R15251 VGND.t84 VGND.t5502 775.568
R15252 VGND.t1263 VGND.t2031 775.568
R15253 VGND.t5713 VGND.t3046 775.568
R15254 VGND.t6732 VGND.t4018 775.568
R15255 VGND.t4103 VGND.t1704 775.568
R15256 VGND.t1754 VGND.t1745 775.568
R15257 VGND.t6628 VGND.t6042 775.568
R15258 VGND.t44 VGND.t1671 775.568
R15259 VGND.t4310 VGND.t5749 775.568
R15260 VGND.t5355 VGND.t1976 775.568
R15261 VGND.t3679 VGND.t3681 775.568
R15262 VGND.t3214 VGND.t3469 770.952
R15263 VGND.t3768 VGND.t568 770.952
R15264 VGND.t3954 VGND.t4537 766.804
R15265 VGND.t6257 VGND.t6740 766.336
R15266 VGND.t6637 VGND 766.336
R15267 VGND.t6728 VGND.t6038 757.102
R15268 VGND.t2863 VGND.t4066 757.102
R15269 VGND.t611 VGND.t2191 757.102
R15270 VGND.t5444 VGND.t5472 757.102
R15271 VGND.t184 VGND.t2604 757.102
R15272 VGND.t6158 VGND.t6074 757.102
R15273 VGND.t206 VGND.t3860 757.102
R15274 VGND.t2411 VGND.t4526 752.486
R15275 VGND.t4497 VGND.t662 748.971
R15276 VGND.t1011 VGND.t2374 747.87
R15277 VGND VGND.t4837 747.87
R15278 VGND.t1965 VGND.t5849 743.254
R15279 VGND.n3480 VGND 738.636
R15280 VGND VGND.n3481 738.636
R15281 VGND VGND.n3482 738.636
R15282 VGND.n3668 VGND 738.636
R15283 VGND VGND.n3673 738.636
R15284 VGND VGND.n3559 738.636
R15285 VGND VGND.n3591 738.636
R15286 VGND VGND.n3623 738.636
R15287 VGND VGND.n3607 738.636
R15288 VGND VGND.n3575 738.636
R15289 VGND VGND.n38 738.636
R15290 VGND VGND.n21 738.636
R15291 VGND VGND.n37 738.636
R15292 VGND.n36 VGND 738.636
R15293 VGND VGND.n3704 738.636
R15294 VGND.t2457 VGND.t6591 738.636
R15295 VGND.t6558 VGND.t6535 738.636
R15296 VGND.t3736 VGND.t3738 738.636
R15297 VGND.n206 VGND.t5958 738.636
R15298 VGND.t5169 VGND.t6269 738.636
R15299 VGND.t3135 VGND.t6265 738.636
R15300 VGND.t6098 VGND.t6261 738.636
R15301 VGND.t2296 VGND.t2817 738.636
R15302 VGND.t3151 VGND 738.636
R15303 VGND VGND.t242 738.636
R15304 VGND.t1000 VGND.t4595 738.636
R15305 VGND.t2971 VGND.t4842 738.636
R15306 VGND VGND.t587 738.636
R15307 VGND VGND.n40 738.636
R15308 VGND.t4559 VGND.t2573 738.636
R15309 VGND VGND.t6639 724.788
R15310 VGND.t1902 VGND 720.17
R15311 VGND.t2267 VGND 720.17
R15312 VGND VGND.t2175 720.17
R15313 VGND VGND.t3136 720.17
R15314 VGND VGND.t2535 720.17
R15315 VGND VGND.t2681 720.17
R15316 VGND VGND.t1747 720.17
R15317 VGND VGND.t2646 720.17
R15318 VGND VGND.t3839 720.17
R15319 VGND.t420 VGND 720.17
R15320 VGND.t2008 VGND 720.17
R15321 VGND VGND.t766 720.17
R15322 VGND VGND.t5332 720.17
R15323 VGND VGND.t3414 720.17
R15324 VGND VGND.t4712 720.17
R15325 VGND VGND.t5119 720.17
R15326 VGND VGND.t6782 720.17
R15327 VGND VGND.t2006 720.17
R15328 VGND VGND.t2715 720.17
R15329 VGND VGND.t1659 720.17
R15330 VGND VGND.t3970 720.17
R15331 VGND VGND.t1083 720.17
R15332 VGND VGND.t2225 720.17
R15333 VGND VGND.t622 720.17
R15334 VGND VGND.t3503 720.17
R15335 VGND VGND.t4826 720.17
R15336 VGND VGND.t61 720.17
R15337 VGND VGND.t5195 720.17
R15338 VGND VGND.t2606 720.17
R15339 VGND VGND.t3193 720.17
R15340 VGND VGND.t4636 720.17
R15341 VGND VGND.t3779 720.17
R15342 VGND VGND.t3890 720.17
R15343 VGND VGND.t3964 720.17
R15344 VGND VGND.t73 720.17
R15345 VGND VGND.t475 720.17
R15346 VGND VGND.t5139 720.17
R15347 VGND VGND.t3581 720.17
R15348 VGND VGND.t352 720.17
R15349 VGND.t3579 VGND 720.17
R15350 VGND.t4178 VGND 720.17
R15351 VGND VGND.t1406 720.17
R15352 VGND VGND.t2059 720.17
R15353 VGND VGND.t4213 720.17
R15354 VGND VGND.t320 720.17
R15355 VGND VGND.t5096 720.17
R15356 VGND VGND.t3048 720.17
R15357 VGND VGND.t686 720.17
R15358 VGND.n283 VGND 720.17
R15359 VGND.t2617 VGND 720.17
R15360 VGND.t2076 VGND 720.17
R15361 VGND.t4903 VGND 720.17
R15362 VGND.t4112 VGND 720.17
R15363 VGND.t5696 VGND 720.17
R15364 VGND.n887 VGND 720.17
R15365 VGND VGND.t5036 720.17
R15366 VGND VGND.n1354 720.17
R15367 VGND VGND.t5435 720.17
R15368 VGND.n1371 VGND 720.17
R15369 VGND VGND.n1245 720.17
R15370 VGND.t4376 VGND 720.17
R15371 VGND.t5178 VGND 720.17
R15372 VGND VGND.t982 720.17
R15373 VGND VGND.t3929 720.17
R15374 VGND VGND.t4319 720.17
R15375 VGND VGND.t4834 720.17
R15376 VGND VGND.t5588 720.17
R15377 VGND VGND.t3271 720.17
R15378 VGND VGND.n1484 720.17
R15379 VGND.t5566 VGND 720.17
R15380 VGND.t861 VGND 720.17
R15381 VGND VGND.t4229 720.17
R15382 VGND VGND.t3475 720.17
R15383 VGND VGND.t2654 720.17
R15384 VGND VGND.t350 720.17
R15385 VGND.t4601 VGND 720.17
R15386 VGND.t2065 VGND 720.17
R15387 VGND VGND.t3709 720.17
R15388 VGND VGND.t694 720.17
R15389 VGND.t901 VGND 720.17
R15390 VGND.t4420 VGND 720.17
R15391 VGND.t5504 VGND 720.17
R15392 VGND.t2786 VGND 720.17
R15393 VGND.t3820 VGND 720.17
R15394 VGND VGND.t3013 720.17
R15395 VGND VGND.t493 720.17
R15396 VGND VGND.t1795 720.17
R15397 VGND VGND.t1991 720.17
R15398 VGND.t168 VGND.t6028 720.17
R15399 VGND.n1731 VGND.t6682 720.17
R15400 VGND.t3033 VGND 720.17
R15401 VGND.t5997 VGND 720.17
R15402 VGND VGND.t2652 720.17
R15403 VGND VGND.t2217 720.17
R15404 VGND VGND.t3237 720.17
R15405 VGND VGND.t1329 720.17
R15406 VGND VGND.t551 720.17
R15407 VGND.t10 VGND.t294 720.17
R15408 VGND VGND.n605 720.17
R15409 VGND.t3773 VGND 720.17
R15410 VGND.t2259 VGND.t1696 720.17
R15411 VGND.t5191 VGND.t1588 720.17
R15412 VGND.t5031 VGND 720.17
R15413 VGND.n726 VGND 720.17
R15414 VGND.t707 VGND 720.17
R15415 VGND.t692 VGND.t6049 720.17
R15416 VGND VGND.t360 720.17
R15417 VGND VGND.t2954 720.17
R15418 VGND VGND.t53 720.17
R15419 VGND VGND.t658 720.17
R15420 VGND.t3389 VGND 720.17
R15421 VGND.t1879 VGND 720.17
R15422 VGND VGND.t2937 720.17
R15423 VGND VGND.t3635 720.17
R15424 VGND VGND.t1122 720.17
R15425 VGND VGND.t5205 720.17
R15426 VGND VGND.t4424 720.17
R15427 VGND VGND.t5098 720.17
R15428 VGND.t2257 VGND 720.17
R15429 VGND.t3977 VGND 720.17
R15430 VGND VGND.t5262 720.17
R15431 VGND VGND.n1076 720.17
R15432 VGND VGND.t55 720.17
R15433 VGND VGND.t3650 720.17
R15434 VGND VGND.t2638 720.17
R15435 VGND.n1077 VGND 720.17
R15436 VGND.t4955 VGND 720.17
R15437 VGND.t823 VGND 720.17
R15438 VGND.t2479 VGND.t5413 720.17
R15439 VGND.t4158 VGND.t429 720.17
R15440 VGND.t3404 VGND 720.17
R15441 VGND VGND.t4245 720.17
R15442 VGND VGND.t1017 720.17
R15443 VGND VGND.t5822 720.17
R15444 VGND VGND.t3300 720.17
R15445 VGND VGND.t5150 720.17
R15446 VGND VGND.t1546 720.17
R15447 VGND VGND.t5818 720.17
R15448 VGND.t4273 VGND 720.17
R15449 VGND VGND.t4586 720.17
R15450 VGND VGND.t2388 720.17
R15451 VGND.n2175 VGND 720.17
R15452 VGND.t865 VGND 720.17
R15453 VGND VGND.t3888 720.17
R15454 VGND VGND.t1036 720.17
R15455 VGND.t5938 VGND 720.17
R15456 VGND.t2232 VGND 720.17
R15457 VGND.t3370 VGND 720.17
R15458 VGND.t3471 VGND 720.17
R15459 VGND.t3491 VGND 720.17
R15460 VGND.t2795 VGND 720.17
R15461 VGND VGND.t3701 720.17
R15462 VGND VGND.t4548 720.17
R15463 VGND.t1591 VGND 720.17
R15464 VGND.t3917 VGND 720.17
R15465 VGND.t3241 VGND 720.17
R15466 VGND.t3967 VGND 720.17
R15467 VGND.t964 VGND 720.17
R15468 VGND VGND.t3915 720.17
R15469 VGND VGND.t358 720.17
R15470 VGND VGND.t3628 720.17
R15471 VGND VGND.t3900 720.17
R15472 VGND VGND.t4265 720.17
R15473 VGND VGND.t3239 720.17
R15474 VGND VGND.t2035 720.17
R15475 VGND.t1070 VGND.t2015 720.17
R15476 VGND VGND.t5238 720.17
R15477 VGND VGND.t1917 720.17
R15478 VGND VGND.t4196 720.17
R15479 VGND.t4170 VGND 720.17
R15480 VGND.t3776 VGND 720.17
R15481 VGND.t5248 VGND 720.17
R15482 VGND VGND.n521 720.17
R15483 VGND.t5732 VGND.t6513 720.17
R15484 VGND VGND.t1485 720.17
R15485 VGND VGND.t2234 720.17
R15486 VGND VGND.t560 720.17
R15487 VGND VGND.t3243 720.17
R15488 VGND VGND.t1400 720.17
R15489 VGND VGND.t6184 720.17
R15490 VGND VGND.t1825 720.17
R15491 VGND VGND.t397 720.17
R15492 VGND VGND.t3662 720.17
R15493 VGND VGND.t5193 720.17
R15494 VGND VGND.t3024 720.17
R15495 VGND VGND.t6748 720.17
R15496 VGND.t4546 VGND 720.17
R15497 VGND.t6808 VGND 720.17
R15498 VGND.t4428 VGND 720.17
R15499 VGND.t3987 VGND 720.17
R15500 VGND.t1283 VGND 720.17
R15501 VGND.t2498 VGND 720.17
R15502 VGND VGND.t3913 720.17
R15503 VGND VGND.t4039 720.17
R15504 VGND VGND.t909 720.17
R15505 VGND VGND.t3921 720.17
R15506 VGND VGND.t879 720.17
R15507 VGND VGND.t5478 720.17
R15508 VGND VGND.t2670 720.17
R15509 VGND VGND.t3862 720.17
R15510 VGND VGND.t1805 720.17
R15511 VGND VGND.t375 720.17
R15512 VGND VGND.t3782 720.17
R15513 VGND.t497 VGND 720.17
R15514 VGND.t2351 VGND 720.17
R15515 VGND.t521 VGND 720.17
R15516 VGND.t2887 VGND 720.17
R15517 VGND.t5626 VGND 720.17
R15518 VGND.t5802 VGND 720.17
R15519 VGND VGND.t3391 720.17
R15520 VGND VGND.t3569 720.17
R15521 VGND VGND.t2701 720.17
R15522 VGND.t547 VGND 720.17
R15523 VGND.t3217 VGND 720.17
R15524 VGND VGND.t5594 720.17
R15525 VGND VGND.t1995 720.17
R15526 VGND VGND.t3368 720.17
R15527 VGND VGND.t5556 720.17
R15528 VGND.t339 VGND 720.17
R15529 VGND VGND.t3028 720.17
R15530 VGND VGND.t3880 720.17
R15531 VGND.t3074 VGND 720.17
R15532 VGND.t1386 VGND 720.17
R15533 VGND VGND.t4237 720.17
R15534 VGND.t1491 VGND 720.17
R15535 VGND.t613 VGND 720.17
R15536 VGND VGND.t5810 720.17
R15537 VGND VGND.t4363 720.17
R15538 VGND VGND.t4372 720.17
R15539 VGND.t1741 VGND 720.17
R15540 VGND VGND.n2092 720.17
R15541 VGND VGND.t5417 720.17
R15542 VGND VGND.t4735 720.17
R15543 VGND VGND.t2966 720.17
R15544 VGND VGND.t3600 720.17
R15545 VGND VGND.t2112 720.17
R15546 VGND.t1578 VGND 720.17
R15547 VGND VGND.t5221 720.17
R15548 VGND VGND.t5175 720.17
R15549 VGND.t3279 VGND.t2723 720.17
R15550 VGND.t5986 VGND 720.17
R15551 VGND.t2327 VGND 720.17
R15552 VGND VGND.t6089 720.17
R15553 VGND VGND.t2998 720.17
R15554 VGND VGND.t845 720.17
R15555 VGND VGND.t1204 720.17
R15556 VGND VGND.t838 720.17
R15557 VGND VGND.t3234 720.17
R15558 VGND.t848 VGND 720.17
R15559 VGND.t531 VGND 720.17
R15560 VGND.t2753 VGND 720.17
R15561 VGND.t3458 VGND 720.17
R15562 VGND VGND.t6055 720.17
R15563 VGND VGND.t2969 720.17
R15564 VGND VGND.t3088 720.17
R15565 VGND VGND.t481 720.17
R15566 VGND.t4639 VGND 720.17
R15567 VGND.t2844 VGND 720.17
R15568 VGND.t1085 VGND 720.17
R15569 VGND.t3161 VGND 720.17
R15570 VGND VGND.t6176 720.17
R15571 VGND VGND.t367 720.17
R15572 VGND VGND.t1118 720.17
R15573 VGND VGND.t4389 720.17
R15574 VGND.t1977 VGND 720.17
R15575 VGND.t1712 VGND 720.17
R15576 VGND.t3228 VGND 720.17
R15577 VGND VGND.t3552 720.17
R15578 VGND VGND.t67 720.17
R15579 VGND VGND.t5454 720.17
R15580 VGND.t549 VGND 720.17
R15581 VGND VGND.t1728 720.17
R15582 VGND VGND.t656 720.17
R15583 VGND VGND.t3195 720.17
R15584 VGND VGND.t2922 720.17
R15585 VGND.t6291 VGND.t6792 715.554
R15586 VGND VGND.t6231 713.307
R15587 VGND.t3478 VGND.t4534 713.307
R15588 VGND.t6031 VGND.t29 713.307
R15589 VGND.t175 VGND.t28 713.307
R15590 VGND.t6693 VGND.t3740 710.938
R15591 VGND.t3937 VGND.n283 701.706
R15592 VGND.t5046 VGND.n887 701.706
R15593 VGND.t6553 VGND.n1370 701.706
R15594 VGND.t2361 VGND.t5776 701.706
R15595 VGND.t2305 VGND.t899 701.706
R15596 VGND.t5787 VGND.t4168 701.706
R15597 VGND.t5533 VGND.n840 701.706
R15598 VGND.t6057 VGND.t1346 701.706
R15599 VGND.t3929 VGND.t1352 701.706
R15600 VGND.t37 VGND.t2196 701.706
R15601 VGND.t2241 VGND.t471 701.706
R15602 VGND.t6788 VGND.t3495 701.706
R15603 VGND.t1785 VGND.t3426 701.706
R15604 VGND.t5229 VGND.t1161 701.706
R15605 VGND.t2465 VGND.t4874 701.706
R15606 VGND.t2592 VGND.t705 701.706
R15607 VGND.t6096 VGND.t5504 701.706
R15608 VGND.t6155 VGND.t4936 701.706
R15609 VGND.t479 VGND.t3416 701.706
R15610 VGND.t569 VGND.t3995 701.706
R15611 VGND VGND.t3726 701.706
R15612 VGND.t6197 VGND.t5995 701.706
R15613 VGND.t6202 VGND.t5059 701.706
R15614 VGND.t2279 VGND.t5034 701.706
R15615 VGND.t286 VGND 701.706
R15616 VGND.t3884 VGND.t6379 701.706
R15617 VGND.t2642 VGND 701.706
R15618 VGND.t2260 VGND.n655 701.706
R15619 VGND.t3100 VGND.t2797 701.706
R15620 VGND.n625 VGND.t181 701.706
R15621 VGND.t2567 VGND.n2206 701.706
R15622 VGND.t1446 VGND.t3623 701.706
R15623 VGND.t3453 VGND.t4968 701.706
R15624 VGND.t4493 VGND.t5081 701.706
R15625 VGND.t6577 VGND.t6300 701.706
R15626 VGND VGND.t1673 701.706
R15627 VGND.t3652 VGND.t6045 701.706
R15628 VGND.t5029 VGND.t2213 701.706
R15629 VGND.t5141 VGND.t2731 701.706
R15630 VGND.t2386 VGND.t1629 701.706
R15631 VGND.t6413 VGND.n565 701.706
R15632 VGND.t2380 VGND.t2812 700.943
R15633 VGND.t4192 VGND.n1349 697.088
R15634 VGND.t718 VGND.t4163 697.088
R15635 VGND VGND.n151 695.473
R15636 VGND.t2941 VGND.t6347 692.472
R15637 VGND.t6319 VGND.t2379 686.558
R15638 VGND.t3379 VGND.t6655 683.24
R15639 VGND VGND.t771 683.24
R15640 VGND VGND.t6436 683.24
R15641 VGND.t3606 VGND.t5759 683.24
R15642 VGND.t5886 VGND.t5298 683.24
R15643 VGND VGND.t97 683.24
R15644 VGND.t4283 VGND 683.24
R15645 VGND.n776 VGND.t6032 683.24
R15646 VGND.t3536 VGND.t948 683.24
R15647 VGND.t5691 VGND.t3325 683.24
R15648 VGND.t6650 VGND.t345 683.24
R15649 VGND VGND.t6708 683.24
R15650 VGND.t4669 VGND.t5376 683.24
R15651 VGND.t280 VGND.t1187 683.24
R15652 VGND.t276 VGND.t6430 683.24
R15653 VGND.t272 VGND.t6502 683.24
R15654 VGND.t6117 VGND 683.24
R15655 VGND.t2937 VGND.t1395 683.24
R15656 VGND.t24 VGND.t986 683.24
R15657 VGND.t1485 VGND.t1754 683.24
R15658 VGND VGND.t42 683.24
R15659 VGND VGND.t6506 683.24
R15660 VGND.t6507 VGND 678.622
R15661 VGND.t1538 VGND.t233 678.622
R15662 VGND.t6433 VGND 678.622
R15663 VGND VGND.t6575 678.622
R15664 VGND.t1216 VGND.t301 678.622
R15665 VGND.t6537 VGND.t6556 677.641
R15666 VGND.t4223 VGND.n899 674.006
R15667 VGND.t2608 VGND 674.006
R15668 VGND.t5395 VGND.t2608 674.006
R15669 VGND.t3434 VGND 674.006
R15670 VGND.t4824 VGND.t3434 674.006
R15671 VGND.t1774 VGND.t4252 674.006
R15672 VGND.t5984 VGND.t1319 674.006
R15673 VGND.t1507 VGND.t4870 674.006
R15674 VGND.t5662 VGND.t6757 674.006
R15675 VGND.t1546 VGND.t1422 674.006
R15676 VGND.t5666 VGND 674.006
R15677 VGND.t3628 VGND.t5666 674.006
R15678 VGND.t942 VGND.t3640 674.006
R15679 VGND.t1426 VGND.t4660 674.006
R15680 VGND.t315 VGND 674.006
R15681 VGND VGND.t4457 674.006
R15682 VGND.t2964 VGND 674.006
R15683 VGND.t5175 VGND.t1649 674.006
R15684 VGND.t5257 VGND.t2814 674.006
R15685 VGND.t3410 VGND.t6737 665.745
R15686 VGND.t1838 VGND 664.774
R15687 VGND.t6012 VGND.t5048 664.774
R15688 VGND.t6010 VGND.t5044 664.774
R15689 VGND.t771 VGND.t5284 664.774
R15690 VGND.t5759 VGND 664.774
R15691 VGND.t5298 VGND 664.774
R15692 VGND VGND.t36 664.774
R15693 VGND.t4962 VGND.t6106 664.774
R15694 VGND.t6530 VGND.t871 664.774
R15695 VGND VGND.t1812 664.774
R15696 VGND.t6665 VGND 664.774
R15697 VGND.t3064 VGND.t5783 664.774
R15698 VGND.t2469 VGND 664.774
R15699 VGND.t6515 VGND.t326 664.774
R15700 VGND.t2677 VGND.t6160 664.774
R15701 VGND.t6780 VGND.t6413 664.774
R15702 VGND.t2600 VGND 660.157
R15703 VGND VGND.t4414 660.157
R15704 VGND.t5849 VGND 660.157
R15705 VGND.t6153 VGND.t938 655.54
R15706 VGND.t6666 VGND.t3058 650.923
R15707 VGND.t6641 VGND.t4895 650.893
R15708 VGND.t1100 VGND 646.308
R15709 VGND.t6593 VGND.t6582 646.308
R15710 VGND.t6443 VGND 646.308
R15711 VGND.t1424 VGND 646.308
R15712 VGND.t6240 VGND.t6541 646.308
R15713 VGND VGND.t5787 646.308
R15714 VGND.t3026 VGND.t2241 646.308
R15715 VGND.t6251 VGND.t3328 646.308
R15716 VGND.t6477 VGND 646.308
R15717 VGND.t6486 VGND 646.308
R15718 VGND.t3070 VGND.t4086 646.308
R15719 VGND.t2374 VGND 646.308
R15720 VGND.t4053 VGND.t4049 646.308
R15721 VGND.t3104 VGND.t4263 646.308
R15722 VGND.t6387 VGND.t4589 646.308
R15723 VGND.t6522 VGND 646.308
R15724 VGND.t6316 VGND.t1394 646.308
R15725 VGND.t1512 VGND.t3583 646.308
R15726 VGND.t214 VGND.t1755 646.308
R15727 VGND.t4856 VGND.n567 646.308
R15728 VGND.n289 VGND.t6536 641.976
R15729 VGND.t6584 VGND.t1787 627.841
R15730 VGND.t264 VGND.t6648 627.841
R15731 VGND.t5393 VGND 627.841
R15732 VGND.t3324 VGND.t5692 627.841
R15733 VGND.t6135 VGND.t2827 627.841
R15734 VGND VGND.t4933 627.841
R15735 VGND.t4846 VGND.t6598 627.841
R15736 VGND VGND.t4846 627.841
R15737 VGND.t1678 VGND.t6520 627.841
R15738 VGND.t4146 VGND.t6578 627.841
R15739 VGND VGND.t84 627.841
R15740 VGND.t6647 VGND.t1377 627.841
R15741 VGND VGND.t2763 627.841
R15742 VGND.t6137 VGND 624.144
R15743 VGND.t4057 VGND.t4412 623.225
R15744 VGND.t4524 VGND.t1410 623.225
R15745 VGND.t4837 VGND.t274 618.609
R15746 VGND.t4076 VGND 613.991
R15747 VGND.t2818 VGND.t919 609.375
R15748 VGND.t5645 VGND.t5277 609.375
R15749 VGND.t4861 VGND.n1490 609.375
R15750 VGND.t2191 VGND 609.375
R15751 VGND.t5692 VGND.t6466 609.375
R15752 VGND.t3730 VGND.t3324 609.375
R15753 VGND.t5817 VGND 609.375
R15754 VGND.t2817 VGND 609.375
R15755 VGND.t5253 VGND.t5736 609.375
R15756 VGND VGND.t5444 609.375
R15757 VGND.t4550 VGND.t3753 609.375
R15758 VGND VGND.t1000 609.375
R15759 VGND.t5893 VGND.t6456 609.375
R15760 VGND.t6311 VGND.t5813 609.375
R15761 VGND.t4859 VGND.t1402 609.375
R15762 VGND.t637 VGND 609.375
R15763 VGND.t4991 VGND 609.375
R15764 VGND.t2243 VGND.t3410 606.311
R15765 VGND.t4905 VGND.t6349 604.76
R15766 VGND.t230 VGND.t5643 604.76
R15767 VGND VGND.t208 595.527
R15768 VGND.t6422 VGND 595.527
R15769 VGND.t4530 VGND.t304 595.527
R15770 VGND.t6695 VGND.t3658 590.909
R15771 VGND.t3336 VGND.t2238 590.909
R15772 VGND.n1494 VGND.t2246 590.909
R15773 VGND.t6315 VGND 590.909
R15774 VGND.t6148 VGND.t865 590.909
R15775 VGND VGND.t4644 586.293
R15776 VGND.t2664 VGND.t6433 581.677
R15777 VGND.t5794 VGND 572.443
R15778 VGND VGND.t3519 572.443
R15779 VGND VGND.t4897 572.443
R15780 VGND.t6775 VGND.t4028 572.443
R15781 VGND.t2869 VGND.t6227 572.443
R15782 VGND.t2867 VGND.t6226 572.443
R15783 VGND.t5279 VGND 572.443
R15784 VGND.t5305 VGND.t801 572.443
R15785 VGND VGND.t6260 572.443
R15786 VGND VGND.t393 572.443
R15787 VGND.t395 VGND.t3262 572.443
R15788 VGND.t1218 VGND.n583 572.443
R15789 VGND VGND.t2178 572.443
R15790 VGND.t6333 VGND.t3144 572.443
R15791 VGND.t179 VGND.t3148 572.443
R15792 VGND.t326 VGND.t3250 572.443
R15793 VGND.t1704 VGND 572.443
R15794 VGND.t2419 VGND.t6151 567.827
R15795 VGND.t1860 VGND 563.211
R15796 VGND VGND.t5912 563.211
R15797 VGND VGND.t1607 563.211
R15798 VGND VGND.t2100 563.211
R15799 VGND VGND.t3420 563.211
R15800 VGND.t2725 VGND 563.211
R15801 VGND VGND.t2544 558.595
R15802 VGND.t3224 VGND.t786 558.595
R15803 VGND.t2596 VGND.t2504 553.977
R15804 VGND.t4365 VGND.t6678 553.977
R15805 VGND.t774 VGND.t3139 553.977
R15806 VGND.t227 VGND.t5182 553.977
R15807 VGND.t450 VGND.t6101 553.977
R15808 VGND.t6099 VGND.n794 553.977
R15809 VGND.t6473 VGND.t4781 553.977
R15810 VGND.t831 VGND.t6522 553.977
R15811 VGND.t121 VGND.t296 553.977
R15812 VGND.t6717 VGND.t290 553.977
R15813 VGND.t515 VGND.t6312 553.977
R15814 VGND.t1112 VGND.t6422 553.977
R15815 VGND.t5242 VGND 553.977
R15816 VGND.t6002 VGND.t5087 553.977
R15817 VGND.t526 VGND.t3156 549.361
R15818 VGND.t1251 VGND.t177 549.361
R15819 VGND.t6341 VGND.t6661 549.361
R15820 VGND.t165 VGND.t6671 549.361
R15821 VGND.t3128 VGND.t1460 544.745
R15822 VGND.t2118 VGND.t2990 544.745
R15823 VGND.t5419 VGND.t827 544.745
R15824 VGND.t1057 VGND.t4335 544.745
R15825 VGND.t2784 VGND.t1072 544.745
R15826 VGND.t5403 VGND.t3909 544.745
R15827 VGND.t1681 VGND.t4346 544.745
R15828 VGND.t2996 VGND.t721 544.745
R15829 VGND.t2375 VGND.t3191 544.745
R15830 VGND.t2945 VGND 540.129
R15831 VGND VGND.t6343 540.129
R15832 VGND.t2697 VGND 540.129
R15833 VGND VGND.t1251 540.129
R15834 VGND VGND.t1255 540.129
R15835 VGND VGND.t5747 540.129
R15836 VGND.t6671 VGND 540.129
R15837 VGND.t301 VGND 540.129
R15838 VGND.t3252 VGND 540.129
R15839 VGND VGND.t2430 535.511
R15840 VGND VGND.t2434 535.511
R15841 VGND VGND.t4729 535.511
R15842 VGND VGND.t2436 535.511
R15843 VGND.t3939 VGND 535.511
R15844 VGND.t6212 VGND 535.511
R15845 VGND VGND.t4980 535.511
R15846 VGND VGND.t3334 535.511
R15847 VGND VGND.t3565 535.511
R15848 VGND.t1665 VGND 535.511
R15849 VGND VGND.t4221 535.511
R15850 VGND.t5463 VGND 535.511
R15851 VGND.t4718 VGND 535.511
R15852 VGND.t3644 VGND 535.511
R15853 VGND VGND.t2132 535.511
R15854 VGND VGND.t323 535.511
R15855 VGND VGND.t3357 535.511
R15856 VGND.t2516 VGND 535.511
R15857 VGND.t2524 VGND 535.511
R15858 VGND VGND.t5050 535.511
R15859 VGND.t6014 VGND 535.511
R15860 VGND VGND.t4885 535.511
R15861 VGND.t3341 VGND 535.511
R15862 VGND VGND.t2631 535.511
R15863 VGND.t2629 VGND 535.511
R15864 VGND.t885 VGND 535.511
R15865 VGND.t3800 VGND 535.511
R15866 VGND.t2321 VGND 535.511
R15867 VGND.t4294 VGND.n1355 535.511
R15868 VGND.t4930 VGND.t6504 535.511
R15869 VGND VGND.t6498 535.511
R15870 VGND.t1455 VGND.t1609 535.511
R15871 VGND VGND.t6220 535.511
R15872 VGND.t3446 VGND 535.511
R15873 VGND VGND.t6553 535.511
R15874 VGND VGND.t1849 535.511
R15875 VGND.t2082 VGND 535.511
R15876 VGND.t2169 VGND 535.511
R15877 VGND.t899 VGND 535.511
R15878 VGND.t768 VGND 535.511
R15879 VGND.t5054 VGND 535.511
R15880 VGND.t3886 VGND 535.511
R15881 VGND.t14 VGND 535.511
R15882 VGND.t3156 VGND 535.511
R15883 VGND.t1862 VGND 535.511
R15884 VGND VGND.t115 535.511
R15885 VGND.t642 VGND 535.511
R15886 VGND VGND.t187 535.511
R15887 VGND.t4063 VGND 535.511
R15888 VGND VGND.t6373 535.511
R15889 VGND VGND.t6355 535.511
R15890 VGND VGND.t6353 535.511
R15891 VGND.t6258 VGND 535.511
R15892 VGND.t104 VGND 535.511
R15893 VGND.t952 VGND 535.511
R15894 VGND.t3432 VGND 535.511
R15895 VGND VGND.t3482 535.511
R15896 VGND.t3485 VGND 535.511
R15897 VGND.t3268 VGND.t6396 535.511
R15898 VGND VGND.t6206 535.511
R15899 VGND.t3060 VGND 535.511
R15900 VGND.t6216 VGND 535.511
R15901 VGND.t5425 VGND 535.511
R15902 VGND VGND.t4333 535.511
R15903 VGND VGND.t5231 535.511
R15904 VGND.t1192 VGND 535.511
R15905 VGND.t1028 VGND 535.511
R15906 VGND VGND.t2465 535.511
R15907 VGND.t4275 VGND 535.511
R15908 VGND VGND.t329 535.511
R15909 VGND VGND.t1009 535.511
R15910 VGND.t110 VGND 535.511
R15911 VGND.t6662 VGND 535.511
R15912 VGND.t757 VGND 535.511
R15913 VGND VGND.t27 535.511
R15914 VGND VGND.t6155 535.511
R15915 VGND.t3416 VGND 535.511
R15916 VGND VGND.t2056 535.511
R15917 VGND.t6545 VGND 535.511
R15918 VGND VGND.t466 535.511
R15919 VGND VGND.t470 535.511
R15920 VGND VGND.t5954 535.511
R15921 VGND VGND.t6197 535.511
R15922 VGND VGND.t6649 535.511
R15923 VGND VGND.t6475 535.511
R15924 VGND.t6673 VGND 535.511
R15925 VGND VGND.t6202 535.511
R15926 VGND.t3850 VGND.t5316 535.511
R15927 VGND.t6193 VGND 535.511
R15928 VGND.t5684 VGND 535.511
R15929 VGND.t1768 VGND 535.511
R15930 VGND VGND.t2275 535.511
R15931 VGND VGND.t1605 535.511
R15932 VGND VGND.t1501 535.511
R15933 VGND VGND.t2907 535.511
R15934 VGND VGND.t5902 535.511
R15935 VGND.t913 VGND 535.511
R15936 VGND VGND.t3814 535.511
R15937 VGND.t189 VGND 535.511
R15938 VGND.t130 VGND 535.511
R15939 VGND VGND.t3157 535.511
R15940 VGND.t3149 VGND.n593 535.511
R15941 VGND.t950 VGND 535.511
R15942 VGND VGND.t4057 535.511
R15943 VGND VGND.t3771 535.511
R15944 VGND VGND.t2813 535.511
R15945 VGND VGND.t5089 535.511
R15946 VGND.t6321 VGND 535.511
R15947 VGND VGND.t5344 535.511
R15948 VGND.t6104 VGND 535.511
R15949 VGND VGND.t6365 535.511
R15950 VGND VGND.t2400 535.511
R15951 VGND.t2689 VGND 535.511
R15952 VGND.t5686 VGND 535.511
R15953 VGND.t1555 VGND 535.511
R15954 VGND.t2958 VGND 535.511
R15955 VGND.t3991 VGND 535.511
R15956 VGND.t5898 VGND 535.511
R15957 VGND.t505 VGND 535.511
R15958 VGND VGND.t1653 535.511
R15959 VGND.t535 VGND 535.511
R15960 VGND VGND.t5411 535.511
R15961 VGND.t2477 VGND 535.511
R15962 VGND VGND.t887 535.511
R15963 VGND.t4315 VGND 535.511
R15964 VGND.t6416 VGND 535.511
R15965 VGND VGND.t248 535.511
R15966 VGND.t2874 VGND 535.511
R15967 VGND VGND.t4959 535.511
R15968 VGND.t4254 VGND 535.511
R15969 VGND.t6452 VGND 535.511
R15970 VGND VGND.t6448 535.511
R15971 VGND.t117 VGND.t4418 535.511
R15972 VGND VGND.t4656 535.511
R15973 VGND VGND.t131 535.511
R15974 VGND.t6375 VGND 535.511
R15975 VGND VGND.t6357 535.511
R15976 VGND VGND.t6120 535.511
R15977 VGND.t6122 VGND 535.511
R15978 VGND.t6514 VGND.t5769 535.511
R15979 VGND.t6415 VGND.t3752 535.511
R15980 VGND.t6500 VGND.t6188 535.511
R15981 VGND.n2175 VGND.t583 535.511
R15982 VGND.t5366 VGND 535.511
R15983 VGND VGND.t5370 535.511
R15984 VGND VGND.t2567 535.511
R15985 VGND.t6579 VGND 535.511
R15986 VGND.t2571 VGND 535.511
R15987 VGND VGND.t6371 535.511
R15988 VGND VGND.t1312 535.511
R15989 VGND.t1323 VGND 535.511
R15990 VGND.t5993 VGND 535.511
R15991 VGND.t4382 VGND 535.511
R15992 VGND.t5664 VGND 535.511
R15993 VGND VGND.t603 535.511
R15994 VGND.t1068 VGND 535.511
R15995 VGND VGND.t2017 535.511
R15996 VGND.t5719 VGND 535.511
R15997 VGND.t6127 VGND 535.511
R15998 VGND VGND.t3711 535.511
R15999 VGND.t2502 VGND 535.511
R16000 VGND.t216 VGND.t4863 535.511
R16001 VGND VGND.t4889 535.511
R16002 VGND.t4403 VGND 535.511
R16003 VGND VGND.t6377 535.511
R16004 VGND VGND.t2102 535.511
R16005 VGND.t2096 VGND 535.511
R16006 VGND VGND.t5757 535.511
R16007 VGND.t1294 VGND 535.511
R16008 VGND.t1520 VGND 535.511
R16009 VGND.t4972 VGND 535.511
R16010 VGND VGND.t1446 535.511
R16011 VGND.t4968 VGND 535.511
R16012 VGND.t2247 VGND 535.511
R16013 VGND.t6045 VGND 535.511
R16014 VGND.t313 VGND 535.511
R16015 VGND VGND.t509 535.511
R16016 VGND.t2731 VGND 535.511
R16017 VGND VGND.t3835 535.511
R16018 VGND.t5609 VGND 535.511
R16019 VGND.t2727 VGND 535.511
R16020 VGND VGND.t2721 535.511
R16021 VGND.t3281 VGND 535.511
R16022 VGND VGND.t3277 535.511
R16023 VGND.t3785 VGND 535.511
R16024 VGND.t6331 VGND 535.511
R16025 VGND VGND.t128 535.511
R16026 VGND.t3979 VGND 535.511
R16027 VGND.t6361 VGND 535.511
R16028 VGND VGND.t4540 535.511
R16029 VGND.t3610 VGND.t6746 521.663
R16030 VGND.t4841 VGND.t6573 521.663
R16031 VGND.t4680 VGND.t1679 521.663
R16032 VGND.t4308 VGND.t3812 521.663
R16033 VGND.t5980 VGND.t6022 521.663
R16034 VGND VGND.t6218 517.148
R16035 VGND VGND.t1105 517.148
R16036 VGND VGND.t6214 517.148
R16037 VGND.t4227 VGND.t1902 517.045
R16038 VGND.t3136 VGND.t4343 517.045
R16039 VGND.t1747 VGND.t3962 517.045
R16040 VGND.t4471 VGND.t420 517.045
R16041 VGND.t5332 VGND.t4752 517.045
R16042 VGND.t5119 VGND.t1694 517.045
R16043 VGND.t2715 VGND.t2487 517.045
R16044 VGND.t1083 VGND.t2528 517.045
R16045 VGND.t3503 VGND.t1667 517.045
R16046 VGND.t5195 VGND.t3319 517.045
R16047 VGND.t4636 VGND.t2284 517.045
R16048 VGND.t3964 VGND.t5820 517.045
R16049 VGND.t5139 VGND.t5338 517.045
R16050 VGND.t5353 VGND.t3579 517.045
R16051 VGND.t2059 VGND.t5117 517.045
R16052 VGND.n43 VGND.t1237 517.045
R16053 VGND.n282 VGND.t5928 517.045
R16054 VGND.t2063 VGND.t1618 517.045
R16055 VGND.t2735 VGND.t2076 517.045
R16056 VGND.t5234 VGND.t2737 517.045
R16057 VGND.t299 VGND.t3705 517.045
R16058 VGND.t1379 VGND.t3882 517.045
R16059 VGND.t4022 VGND.t4269 517.045
R16060 VGND.t1462 VGND.t3128 517.045
R16061 VGND.t1460 VGND.t3130 517.045
R16062 VGND.n895 VGND.n894 517.045
R16063 VGND.t3614 VGND.t6569 517.045
R16064 VGND.t3528 VGND.t5673 517.045
R16065 VGND.t2520 VGND.t3528 517.045
R16066 VGND VGND.t1454 517.045
R16067 VGND.t2838 VGND 517.045
R16068 VGND.t2990 VGND.t2116 517.045
R16069 VGND.t2992 VGND.t2118 517.045
R16070 VGND.t3290 VGND.t2371 517.045
R16071 VGND.t3004 VGND.t1736 517.045
R16072 VGND.t1777 VGND.t1835 517.045
R16073 VGND.t6350 VGND.t5288 517.045
R16074 VGND.t982 VGND.t593 517.045
R16075 VGND.t143 VGND 517.045
R16076 VGND VGND.t527 517.045
R16077 VGND.t99 VGND 517.045
R16078 VGND VGND.t99 517.045
R16079 VGND.t3267 VGND 517.045
R16080 VGND.t827 VGND.t5421 517.045
R16081 VGND.t825 VGND.t5419 517.045
R16082 VGND.t4335 VGND.t1055 517.045
R16083 VGND.t4337 VGND.t1057 517.045
R16084 VGND.t2054 VGND.t4420 517.045
R16085 VGND.t119 VGND.t6446 517.045
R16086 VGND.t6446 VGND.t3153 517.045
R16087 VGND.t3153 VGND.t173 517.045
R16088 VGND.t1553 VGND.t3633 517.045
R16089 VGND.t6710 VGND 517.045
R16090 VGND.t4670 VGND 517.045
R16091 VGND VGND.t1333 517.045
R16092 VGND.t5113 VGND.t3033 517.045
R16093 VGND.t3974 VGND.t3305 517.045
R16094 VGND.t5951 VGND.t5997 517.045
R16095 VGND.n1124 VGND.t5223 517.045
R16096 VGND VGND.t155 517.045
R16097 VGND.t436 VGND.t1898 517.045
R16098 VGND.t5125 VGND.t1306 517.045
R16099 VGND.t3493 VGND.t4164 517.045
R16100 VGND.t5439 VGND.t2660 517.045
R16101 VGND.t4339 VGND.t6092 517.045
R16102 VGND.t333 VGND.t1900 517.045
R16103 VGND.t5568 VGND.t4555 517.045
R16104 VGND.t53 VGND.t2292 517.045
R16105 VGND.t2485 VGND.t2405 517.045
R16106 VGND.t3796 VGND.t3558 517.045
R16107 VGND.t311 VGND.t710 517.045
R16108 VGND.t6186 VGND.t697 517.045
R16109 VGND.t2309 VGND.t1440 517.045
R16110 VGND.t5336 VGND.t1738 517.045
R16111 VGND.t4447 VGND.t4796 517.045
R16112 VGND.t658 VGND.t1997 517.045
R16113 VGND.t3203 VGND.t6543 517.045
R16114 VGND.t6302 VGND.t3203 517.045
R16115 VGND.t4323 VGND.t6302 517.045
R16116 VGND.t96 VGND 517.045
R16117 VGND.t3635 VGND.t1855 517.045
R16118 VGND.t4743 VGND.t2355 517.045
R16119 VGND.t1980 VGND.t5635 517.045
R16120 VGND.t2774 VGND.t962 517.045
R16121 VGND.t1122 VGND.t4786 517.045
R16122 VGND.t4287 VGND.t4491 517.045
R16123 VGND.t4380 VGND.t5362 517.045
R16124 VGND.t1567 VGND.t2805 517.045
R16125 VGND.t1633 VGND.t3460 517.045
R16126 VGND.t4090 VGND.t4552 517.045
R16127 VGND.t807 VGND.t3094 517.045
R16128 VGND.t1308 VGND.t5447 517.045
R16129 VGND.t5205 VGND.t412 517.045
R16130 VGND.t4676 VGND.t3763 517.045
R16131 VGND.t5161 VGND.t4512 517.045
R16132 VGND.t3359 VGND.t6078 517.045
R16133 VGND.t2318 VGND.t4233 517.045
R16134 VGND.t2584 VGND.t1341 517.045
R16135 VGND.t1570 VGND.t1247 517.045
R16136 VGND.t2679 VGND.t3351 517.045
R16137 VGND.t4424 VGND.t3907 517.045
R16138 VGND.t3841 VGND.t1635 517.045
R16139 VGND.t5137 VGND.t5324 517.045
R16140 VGND.t5900 VGND.t3307 517.045
R16141 VGND.t1864 VGND.t4749 517.045
R16142 VGND.t690 VGND.t2069 517.045
R16143 VGND.t3534 VGND.t5544 517.045
R16144 VGND.t1528 VGND.t4478 517.045
R16145 VGND.t5098 VGND.t597 517.045
R16146 VGND.n1077 VGND.t4989 517.045
R16147 VGND.t4245 VGND.t3707 517.045
R16148 VGND.t4674 VGND.t1184 517.045
R16149 VGND.t5841 VGND.t1593 517.045
R16150 VGND.t875 VGND.t629 517.045
R16151 VGND.t1017 VGND.t1989 517.045
R16152 VGND.t1639 VGND.n942 517.045
R16153 VGND.n943 VGND.t5619 517.045
R16154 VGND.t1969 VGND.t2674 517.045
R16155 VGND.t4542 VGND.t3396 517.045
R16156 VGND.t4784 VGND.t1591 517.045
R16157 VGND.t2636 VGND.t1637 517.045
R16158 VGND.t1973 VGND.t2409 517.045
R16159 VGND.t4872 VGND.t1892 517.045
R16160 VGND.t654 VGND.t3917 517.045
R16161 VGND.t3915 VGND.n466 517.045
R16162 VGND.n467 VGND.t6043 517.045
R16163 VGND.t3387 VGND.t2580 517.045
R16164 VGND.t1526 VGND.t2067 517.045
R16165 VGND.t1202 VGND.t562 517.045
R16166 VGND.t2500 VGND.t728 517.045
R16167 VGND.t5320 VGND.t5847 517.045
R16168 VGND.t4100 VGND.t3560 517.045
R16169 VGND.t1359 VGND.t1436 517.045
R16170 VGND.t4196 VGND.t3818 517.045
R16171 VGND.n521 VGND.t1234 517.045
R16172 VGND.t575 VGND.t4641 517.045
R16173 VGND VGND.t5733 517.045
R16174 VGND.t47 VGND 517.045
R16175 VGND.t2626 VGND.t5732 517.045
R16176 VGND.t6630 VGND 517.045
R16177 VGND.t2234 VGND.t591 517.045
R16178 VGND.t764 VGND.t2042 517.045
R16179 VGND.t5109 VGND.t1416 517.045
R16180 VGND.t4137 VGND.t4426 517.045
R16181 VGND.t560 VGND.t5127 517.045
R16182 VGND.t6184 VGND.t6051 517.045
R16183 VGND.t6166 VGND.t5677 517.045
R16184 VGND.t1724 VGND.t617 517.045
R16185 VGND.t3098 VGND.t2933 517.045
R16186 VGND.t1825 VGND.t5970 517.045
R16187 VGND.t4140 VGND.t5077 517.045
R16188 VGND.t4469 VGND.t1278 517.045
R16189 VGND.t4217 VGND.t2289 517.045
R16190 VGND.t5653 VGND.t2050 517.045
R16191 VGND.t5093 VGND.t2263 517.045
R16192 VGND.t2542 VGND.t850 517.045
R16193 VGND.t793 VGND.t318 517.045
R16194 VGND.t3662 VGND.t4696 517.045
R16195 VGND.t1074 VGND.t2784 517.045
R16196 VGND.t1072 VGND.t2782 517.045
R16197 VGND.t1831 VGND.t2634 517.045
R16198 VGND.t991 VGND.t4546 517.045
R16199 VGND.t4580 VGND.t6765 517.045
R16200 VGND.t4219 VGND.t4507 517.045
R16201 VGND.t5668 VGND.t3273 517.045
R16202 VGND.t1414 VGND.t5680 517.045
R16203 VGND.t5521 VGND.t2565 517.045
R16204 VGND.t795 VGND.t503 517.045
R16205 VGND.t4765 VGND.t5313 517.045
R16206 VGND.t4987 VGND.t4428 517.045
R16207 VGND.t1019 VGND.t940 517.045
R16208 VGND.t3621 VGND.t1714 517.045
R16209 VGND.t3806 VGND.t5357 517.045
R16210 VGND.t1580 VGND.t1549 517.045
R16211 VGND.t1559 VGND.t1444 517.045
R16212 VGND.t6750 VGND.t1489 517.045
R16213 VGND.t4621 VGND.t4794 517.045
R16214 VGND.t601 VGND.t3987 517.045
R16215 VGND.t5433 VGND.t1124 517.045
R16216 VGND.t1093 VGND.t1885 517.045
R16217 VGND.t4350 VGND.t6076 517.045
R16218 VGND.t5875 VGND.t4329 517.045
R16219 VGND.t4188 VGND.t4431 517.045
R16220 VGND.t2078 VGND.t2151 517.045
R16221 VGND.t2110 VGND.t1003 517.045
R16222 VGND.t4876 VGND.t1283 517.045
R16223 VGND.t1493 VGND.t2791 517.045
R16224 VGND.t3670 VGND.t4155 517.045
R16225 VGND.t5540 VGND.t2311 517.045
R16226 VGND.t1963 VGND.t3577 517.045
R16227 VGND.t1438 VGND.t1951 517.045
R16228 VGND.t4612 VGND.t2574 517.045
R16229 VGND.t1392 VGND.t2255 517.045
R16230 VGND.t6796 VGND.t2498 517.045
R16231 VGND.t4114 VGND.t3626 517.045
R16232 VGND.t5549 VGND.t5359 517.045
R16233 VGND.t2185 VGND.t3742 517.045
R16234 VGND.t3573 VGND.t1647 517.045
R16235 VGND.t2003 VGND.t1495 517.045
R16236 VGND.t799 VGND.t4914 517.045
R16237 VGND.t1941 VGND.t3720 517.045
R16238 VGND.t3913 VGND.t1871 517.045
R16239 VGND.t5558 VGND.n2492 517.045
R16240 VGND.n2493 VGND.t2108 517.045
R16241 VGND.t3909 VGND.t5401 517.045
R16242 VGND.t3911 VGND.t5403 517.045
R16243 VGND.n2495 VGND.t2038 517.045
R16244 VGND.t3782 VGND.n2496 517.045
R16245 VGND.n2497 VGND.t2855 517.045
R16246 VGND.n406 VGND.t4817 517.045
R16247 VGND.t3068 VGND.n405 517.045
R16248 VGND.t3170 VGND.t4036 517.045
R16249 VGND.t5825 VGND.t2029 517.045
R16250 VGND.t1466 VGND.t978 517.045
R16251 VGND.t1356 VGND.t1174 517.045
R16252 VGND.t5647 VGND.t2755 517.045
R16253 VGND.t3798 VGND.t1043 517.045
R16254 VGND.t1957 VGND.t5626 517.045
R16255 VGND.t5326 VGND.t4710 517.045
R16256 VGND.t3712 VGND.t495 517.045
R16257 VGND.t4271 VGND.t3714 517.045
R16258 VGND.t1530 VGND.t784 517.045
R16259 VGND.t5380 VGND.t1833 517.045
R16260 VGND.t4792 VGND.t2090 517.045
R16261 VGND.t2365 VGND.t4397 517.045
R16262 VGND.t4088 VGND.t5802 517.045
R16263 VGND.t5010 VGND.t1337 517.045
R16264 VGND.t5888 VGND.t3019 517.045
R16265 VGND.t3843 VGND.t3993 517.045
R16266 VGND.t3119 VGND.t4658 517.045
R16267 VGND.t1343 VGND.t5186 517.045
R16268 VGND.t3438 VGND.t4449 517.045
R16269 VGND.t3550 VGND.t2885 517.045
R16270 VGND.t3391 VGND.t5838 517.045
R16271 VGND.t5074 VGND.t3854 517.045
R16272 VGND.t3035 VGND.t5829 517.045
R16273 VGND.t4770 VGND.t5246 517.045
R16274 VGND.t672 VGND.t4891 517.045
R16275 VGND.t2325 VGND.t5959 517.045
R16276 VGND.t5717 VGND.t51 517.045
R16277 VGND.t533 VGND.t3585 517.045
R16278 VGND.t3569 VGND.t1576 517.045
R16279 VGND.t4763 VGND.t2349 517.045
R16280 VGND.t668 VGND.t2189 517.045
R16281 VGND.t4725 VGND.t5407 517.045
R16282 VGND.t3205 VGND.t1657 517.045
R16283 VGND.t5800 VGND.t1222 517.045
R16284 VGND.t3011 VGND.t4356 517.045
R16285 VGND.t5103 VGND.t1210 517.045
R16286 VGND.t2701 VGND.t1331 517.045
R16287 VGND.t3856 VGND.t5105 517.045
R16288 VGND.t4474 VGND.t2789 517.045
R16289 VGND.t1797 VGND.t5468 517.045
R16290 VGND.t5738 VGND.t3230 517.045
R16291 VGND.t958 VGND.t813 517.045
R16292 VGND.t1276 VGND.t5003 517.045
R16293 VGND.t1388 VGND.t2898 517.045
R16294 VGND.t462 VGND.t5449 517.045
R16295 VGND.t4850 VGND.t6815 517.045
R16296 VGND.t2719 VGND.t6767 517.045
R16297 VGND.t4249 VGND.t379 517.045
R16298 VGND.t1107 VGND.t4779 517.045
R16299 VGND.t3646 VGND.t4211 517.045
R16300 VGND.t4927 VGND.t2122 517.045
R16301 VGND.t2215 VGND.t2286 517.045
R16302 VGND.t5594 VGND.t4952 517.045
R16303 VGND.t6802 VGND.t4215 517.045
R16304 VGND.t3183 VGND.t5064 517.045
R16305 VGND.t4304 VGND.t1281 517.045
R16306 VGND.t4482 VGND.t1987 517.045
R16307 VGND.t2147 VGND.t4714 517.045
R16308 VGND.t2303 VGND.t1477 517.045
R16309 VGND.t1995 VGND.t434 517.045
R16310 VGND.t1676 VGND.t1047 517.045
R16311 VGND.t1597 VGND.t3927 517.045
R16312 VGND.t1196 VGND.t4830 517.045
R16313 VGND.t791 VGND.t5201 517.045
R16314 VGND.t4487 VGND.t5574 517.045
R16315 VGND.t1915 VGND.t5861 517.045
R16316 VGND.t3383 VGND.t1432 517.045
R16317 VGND.t3187 VGND.t3792 517.045
R16318 VGND.t1843 VGND.t3637 517.045
R16319 VGND.t4502 VGND.t5269 517.045
R16320 VGND.t5452 VGND.t5318 517.045
R16321 VGND.t1710 VGND.t5730 517.045
R16322 VGND.t3142 VGND.t1599 517.045
R16323 VGND.t5977 VGND.t65 517.045
R16324 VGND.t499 VGND.t6040 517.045
R16325 VGND.t5144 VGND.t6173 517.045
R16326 VGND.n2634 VGND.n2633 517.045
R16327 VGND.t1781 VGND.t1565 517.045
R16328 VGND.t4756 VGND.t1627 517.045
R16329 VGND.t1367 VGND.t1156 517.045
R16330 VGND.t1198 VGND.t4881 517.045
R16331 VGND.t4190 VGND.t4607 517.045
R16332 VGND.t2622 VGND.t2650 517.045
R16333 VGND.t3028 VGND.t4610 517.045
R16334 VGND.t4292 VGND.t712 517.045
R16335 VGND.t3664 VGND.t4698 517.045
R16336 VGND.t2347 VGND.t4202 517.045
R16337 VGND.t2369 VGND.t2307 517.045
R16338 VGND.t1534 VGND.t5930 517.045
R16339 VGND.t3744 VGND.t745 517.045
R16340 VGND.t4665 VGND.t1081 517.045
R16341 VGND.t3880 VGND.t4822 517.045
R16342 VGND.t2402 VGND.t589 517.045
R16343 VGND.t4133 VGND.t4614 517.045
R16344 VGND.t4716 VGND.t4142 517.045
R16345 VGND.t3870 VGND.t1692 517.045
R16346 VGND.t2104 VGND.t3258 517.045
R16347 VGND.t732 VGND.t5771 517.045
R16348 VGND.t5851 VGND.t5602 517.045
R16349 VGND.t4907 VGND.t3074 517.045
R16350 VGND.t2576 VGND.t5437 517.045
R16351 VGND.t2165 VGND.t3442 517.045
R16352 VGND.t1369 VGND.t4444 517.045
R16353 VGND.t1200 VGND.t4300 517.045
R16354 VGND.t4194 VGND.t5947 517.045
R16355 VGND.t3092 VGND.t3656 517.045
R16356 VGND.t3260 VGND.t3868 517.045
R16357 VGND.t3115 VGND.t1386 517.045
R16358 VGND.t1480 VGND.t3666 517.045
R16359 VGND.t2526 VGND.t487 517.045
R16360 VGND.t6018 VGND.t2988 517.045
R16361 VGND.t3394 VGND.t3525 517.045
R16362 VGND.t4183 VGND.t5956 517.045
R16363 VGND.t674 VGND.t4461 517.045
R16364 VGND.t1756 VGND.t3997 517.045
R16365 VGND.t4237 VGND.t1760 517.045
R16366 VGND.t5810 VGND.t4041 517.045
R16367 VGND.t4108 VGND.t1741 517.045
R16368 VGND.t4700 VGND.t485 517.045
R16369 VGND.t6580 VGND.t6304 517.045
R16370 VGND.t4463 VGND.t5067 517.045
R16371 VGND.t5397 VGND.t5553 517.045
R16372 VGND.t2847 VGND.t3587 517.045
R16373 VGND.t5481 VGND.t6034 517.045
R16374 VGND.t2223 VGND.t3925 517.045
R16375 VGND.t2183 VGND.t970 517.045
R16376 VGND.t4352 VGND.t3696 517.045
R16377 VGND.t4735 VGND.t5949 517.045
R16378 VGND.t1298 VGND.t566 517.045
R16379 VGND.t3877 VGND.t1743 517.045
R16380 VGND.t5926 VGND.t4367 517.045
R16381 VGND.t2061 VGND.t3090 517.045
R16382 VGND.t2892 VGND.t3538 517.045
R16383 VGND.t4806 VGND.t5975 517.045
R16384 VGND.t2966 VGND.t2871 517.045
R16385 VGND.t1789 VGND.t1434 517.045
R16386 VGND.t4166 VGND.t3604 517.045
R16387 VGND.t2134 VGND.t1791 517.045
R16388 VGND.t4267 VGND.t3694 517.045
R16389 VGND.t4024 VGND.t5199 517.045
R16390 VGND.t4568 VGND.t5920 517.045
R16391 VGND.t1706 VGND.t4901 517.045
R16392 VGND.t3050 VGND.t995 517.045
R16393 VGND.t2538 VGND.t4440 517.045
R16394 VGND.t3406 VGND.t1716 517.045
R16395 VGND.t2422 VGND.t2749 517.045
R16396 VGND.t3774 VGND.t2426 517.045
R16397 VGND.t5525 VGND.t1726 517.045
R16398 VGND.t972 VGND.t2345 517.045
R16399 VGND.t4451 VGND.t974 517.045
R16400 VGND.t3345 VGND.t1390 517.045
R16401 VGND.n358 VGND.n357 517.045
R16402 VGND.t4346 VGND.t1683 517.045
R16403 VGND.t4348 VGND.t1681 517.045
R16404 VGND.t721 VGND.t2994 517.045
R16405 VGND.t723 VGND.t2996 517.045
R16406 VGND.t3189 VGND.t2375 517.045
R16407 VGND.t3191 VGND.t2377 517.045
R16408 VGND.t3943 VGND.t1869 517.045
R16409 VGND.t4650 VGND 517.045
R16410 VGND.n2969 VGND.t1109 517.045
R16411 VGND.t4045 VGND.n2970 517.045
R16412 VGND.n2971 VGND.t4632 517.045
R16413 VGND.n377 VGND.t4465 517.045
R16414 VGND.t2793 VGND.n376 517.045
R16415 VGND.t1690 VGND.n3074 517.045
R16416 VGND.n3075 VGND.t1645 517.045
R16417 VGND.t1134 VGND.n3076 517.045
R16418 VGND.n3077 VGND.t2578 517.045
R16419 VGND.n369 VGND.t1752 517.045
R16420 VGND.t3402 VGND.n368 517.045
R16421 VGND.t1890 VGND.n3180 517.045
R16422 VGND.n3181 VGND.t747 517.045
R16423 VGND.t3337 VGND.n3182 517.045
R16424 VGND.n3183 VGND.t1993 517.045
R16425 VGND.n362 VGND.t1779 517.045
R16426 VGND.t3292 VGND.n361 517.045
R16427 VGND.t5774 VGND.n3310 517.045
R16428 VGND.n3311 VGND.t519 517.045
R16429 VGND.t5454 VGND.n3312 517.045
R16430 VGND.n3313 VGND.t829 517.045
R16431 VGND.t4591 VGND.n5 517.045
R16432 VGND.n6 VGND.t1045 517.045
R16433 VGND.t656 VGND.n7 517.045
R16434 VGND.n8 VGND.t5761 517.045
R16435 VGND.t401 VGND.t6381 512.429
R16436 VGND.t6442 VGND.t3610 512.429
R16437 VGND.t5510 VGND.t4680 512.429
R16438 VGND.t1910 VGND.t4308 512.429
R16439 VGND.t2430 VGND 498.58
R16440 VGND.t4909 VGND.t3934 498.58
R16441 VGND VGND.t3302 498.58
R16442 VGND.t6659 VGND 498.58
R16443 VGND.t3377 VGND.t3332 498.58
R16444 VGND VGND.t3644 498.58
R16445 VGND VGND.t1858 498.58
R16446 VGND.t2045 VGND 498.58
R16447 VGND VGND.t2518 498.58
R16448 VGND VGND.t6016 498.58
R16449 VGND VGND.t6438 498.58
R16450 VGND VGND.t885 498.58
R16451 VGND.t6504 VGND.t788 498.58
R16452 VGND.t6498 VGND.t4930 498.58
R16453 VGND VGND.t5827 498.58
R16454 VGND.t888 VGND 498.58
R16455 VGND.n1484 VGND.t803 498.58
R16456 VGND.t471 VGND.t1985 498.58
R16457 VGND VGND.t3428 498.58
R16458 VGND.t1099 VGND.t6538 498.58
R16459 VGND.t3484 VGND.t4374 498.58
R16460 VGND.t4279 VGND 498.58
R16461 VGND.t331 VGND 498.58
R16462 VGND VGND.t759 498.58
R16463 VGND.t3837 VGND.t5890 498.58
R16464 VGND.t6208 VGND 498.58
R16465 VGND.t5914 VGND 498.58
R16466 VGND VGND.t6784 498.58
R16467 VGND.t1605 VGND 498.58
R16468 VGND.t4006 VGND 498.58
R16469 VGND.t1245 VGND 498.58
R16470 VGND.t5387 VGND.n593 498.58
R16471 VGND VGND.t1212 498.58
R16472 VGND.t1919 VGND.n732 498.58
R16473 VGND.t6642 VGND 498.58
R16474 VGND.t5089 VGND 498.58
R16475 VGND VGND.t5605 498.58
R16476 VGND.t2687 VGND 498.58
R16477 VGND VGND.t3596 498.58
R16478 VGND VGND.t5686 498.58
R16479 VGND VGND.t3639 498.58
R16480 VGND.t887 VGND 498.58
R16481 VGND.t3630 VGND 498.58
R16482 VGND.t262 VGND 498.58
R16483 VGND.t6618 VGND.n654 498.58
R16484 VGND.t2916 VGND 498.58
R16485 VGND VGND.t2914 498.58
R16486 VGND.t4656 VGND.t3080 498.58
R16487 VGND.t6711 VGND 498.58
R16488 VGND.t5769 VGND.t6122 498.58
R16489 VGND.t3752 VGND.t6514 498.58
R16490 VGND.t6188 VGND.t6415 498.58
R16491 VGND.t3015 VGND 498.58
R16492 VGND VGND.t5870 498.58
R16493 VGND VGND.t5993 498.58
R16494 VGND.t5173 VGND.t4016 498.58
R16495 VGND.t2102 VGND 498.58
R16496 VGND VGND.t1294 498.58
R16497 VGND.t3422 VGND 498.58
R16498 VGND.n404 VGND.t5135 498.58
R16499 VGND VGND.t2727 498.58
R16500 VGND.t5012 VGND 498.58
R16501 VGND VGND.t5215 498.58
R16502 VGND VGND.t191 498.58
R16503 VGND VGND.t6420 498.58
R16504 VGND.t6343 VGND 493.964
R16505 VGND.t3677 VGND 493.964
R16506 VGND VGND.t6577 493.964
R16507 VGND.t4359 VGND.t5910 489.348
R16508 VGND.t1032 VGND.t4361 489.348
R16509 VGND.t4917 VGND.t5660 489.348
R16510 VGND.t2859 VGND.t4919 489.348
R16511 VGND.t2253 VGND.t5572 489.348
R16512 VGND.t114 VGND.t5622 484.731
R16513 VGND.t3590 VGND.t3419 484.731
R16514 VGND.t3139 VGND.t778 480.115
R16515 VGND VGND.t6565 480.115
R16516 VGND.t1572 VGND.t4929 480.115
R16517 VGND VGND.t3972 480.115
R16518 VGND.t2986 VGND.t141 480.115
R16519 VGND.t385 VGND.t6324 480.115
R16520 VGND.t6142 VGND.t5184 480.115
R16521 VGND VGND.t2417 480.115
R16522 VGND.t6680 VGND.t5562 480.115
R16523 VGND.t296 VGND.t1253 480.115
R16524 VGND.t290 VGND.t121 480.115
R16525 VGND.t294 VGND.t6717 480.115
R16526 VGND.t3698 VGND 480.115
R16527 VGND.t4510 VGND.t94 480.115
R16528 VGND.t133 VGND.t4158 480.115
R16529 VGND.t6418 VGND.t1112 480.115
R16530 VGND VGND.t5242 480.115
R16531 VGND.t2388 VGND.t6713 480.115
R16532 VGND.t572 VGND.t6628 480.115
R16533 VGND.t4151 VGND 475.498
R16534 VGND VGND.t1663 470.882
R16535 VGND VGND.t4720 470.882
R16536 VGND VGND.t2941 470.882
R16537 VGND.t1503 VGND 470.882
R16538 VGND.t2905 VGND 470.882
R16539 VGND.t2398 VGND 470.882
R16540 VGND VGND.t2691 470.882
R16541 VGND VGND.t4854 470.882
R16542 VGND.t4957 VGND 470.882
R16543 VGND.t1310 VGND 470.882
R16544 VGND VGND.t1325 470.882
R16545 VGND VGND.t4384 470.882
R16546 VGND.t5755 VGND 470.882
R16547 VGND VGND.t2098 470.882
R16548 VGND VGND.t1522 470.882
R16549 VGND.t1076 VGND 466.264
R16550 VGND.t2820 VGND.t3589 466.264
R16551 VGND.t2432 VGND 461.649
R16552 VGND VGND.t5792 461.649
R16553 VGND.t3521 VGND 461.649
R16554 VGND VGND.t946 461.649
R16555 VGND.t4026 VGND.t6775 461.649
R16556 VGND.t6227 VGND.t2867 461.649
R16557 VGND VGND.t5279 461.649
R16558 VGND.t925 VGND.n200 461.649
R16559 VGND.t389 VGND 461.649
R16560 VGND.t1270 VGND 461.649
R16561 VGND.t454 VGND 461.649
R16562 VGND VGND.t3923 461.649
R16563 VGND VGND.t5615 461.649
R16564 VGND VGND.t1702 461.649
R16565 VGND.t6318 VGND 461.649
R16566 VGND.t3144 VGND.t133 461.649
R16567 VGND.t3148 VGND.t6333 461.649
R16568 VGND.t4651 VGND 461.649
R16569 VGND.t6164 VGND.t5364 461.649
R16570 VGND.t4018 VGND.t5713 461.649
R16571 VGND.t6000 VGND.t4103 461.649
R16572 VGND.t3892 VGND 461.649
R16573 VGND.t5383 VGND 447.798
R16574 VGND.t4961 VGND 447.798
R16575 VGND.t4996 VGND.t4314 447.798
R16576 VGND.t1985 VGND.t3336 443.183
R16577 VGND.t2237 VGND.n1494 443.183
R16578 VGND.t126 VGND.t2602 443.183
R16579 VGND.t6074 VGND.t1933 443.183
R16580 VGND.t2929 VGND.t3979 443.183
R16581 VGND VGND.t6562 438.565
R16582 VGND.t6646 VGND.t2380 436.901
R16583 VGND.t6381 VGND.t5470 429.332
R16584 VGND.t5399 VGND.t230 429.332
R16585 VGND.t5643 VGND.t3768 429.332
R16586 VGND.t5843 VGND.t2221 424.716
R16587 VGND.t21 VGND.t5893 424.716
R16588 VGND.t5813 VGND.t3794 424.716
R16589 VGND.t4654 VGND 424.716
R16590 VGND VGND.t5621 424.716
R16591 VGND.t1402 VGND.t4997 424.716
R16592 VGND.t5085 VGND.t877 424.716
R16593 VGND VGND.t4991 424.716
R16594 VGND VGND.t4077 420.099
R16595 VGND.t1147 VGND 410.866
R16596 VGND.t2939 VGND.t1464 406.25
R16597 VGND.t1412 VGND 406.25
R16598 VGND.t6431 VGND 406.25
R16599 VGND.t6326 VGND 406.25
R16600 VGND.t6578 VGND.t1678 406.25
R16601 VGND.t3199 VGND.t4146 406.25
R16602 VGND.t427 VGND 406.25
R16603 VGND.t1383 VGND 406.25
R16604 VGND.t6715 VGND 406.25
R16605 VGND VGND.t2559 406.25
R16606 VGND.t1262 VGND 406.25
R16607 VGND.t3858 VGND 406.25
R16608 VGND VGND.t4306 406.25
R16609 VGND.t5746 VGND.t2929 406.25
R16610 VGND VGND.t190 406.25
R16611 VGND.t6703 VGND.t6705 401.635
R16612 VGND.t4314 VGND.t3981 401.635
R16613 VGND VGND.t1182 387.784
R16614 VGND.t1178 VGND 387.784
R16615 VGND.t5790 VGND.t2598 387.784
R16616 VGND.t2598 VGND.t6593 387.784
R16617 VGND.t6582 VGND.t2503 387.784
R16618 VGND.t317 VGND 387.784
R16619 VGND.t3684 VGND 387.784
R16620 VGND.t323 VGND 387.784
R16621 VGND VGND.t6744 387.784
R16622 VGND VGND.t4068 387.784
R16623 VGND VGND.t5131 387.784
R16624 VGND.t6541 VGND.t6244 387.784
R16625 VGND.t2384 VGND 387.784
R16626 VGND.t3413 VGND 387.784
R16627 VGND VGND.t2610 387.784
R16628 VGND.t3328 VGND.t104 387.784
R16629 VGND VGND.t1925 387.784
R16630 VGND VGND.t1927 387.784
R16631 VGND VGND.t1929 387.784
R16632 VGND.t4086 VGND.t3485 387.784
R16633 VGND.t100 VGND 387.784
R16634 VGND.t1505 VGND 387.784
R16635 VGND VGND.t6686 387.784
R16636 VGND.t4263 VGND.t6673 387.784
R16637 VGND.t4589 VGND.t3104 387.784
R16638 VGND VGND.t3436 387.784
R16639 VGND VGND.t6524 387.784
R16640 VGND VGND.t3202 387.784
R16641 VGND.t1394 VGND.t6104 387.784
R16642 VGND.t3575 VGND.t6316 387.784
R16643 VGND VGND.t4315 387.784
R16644 VGND.t2861 VGND 387.784
R16645 VGND VGND.t5570 387.784
R16646 VGND.t6146 VGND 387.784
R16647 VGND VGND.t6189 387.784
R16648 VGND VGND.t223 387.784
R16649 VGND VGND.t5664 387.784
R16650 VGND.t4889 VGND.t1512 387.784
R16651 VGND.t1755 VGND.t4403 387.784
R16652 VGND.t4225 VGND.t214 387.784
R16653 VGND VGND.t313 387.784
R16654 VGND.t4459 VGND 387.784
R16655 VGND VGND.t2962 387.784
R16656 VGND VGND.t5056 383.168
R16657 VGND.t208 VGND.t2820 383.168
R16658 VGND.t6635 VGND.t2329 373.935
R16659 VGND.t3981 VGND.t193 373.935
R16660 VGND VGND.t1838 369.318
R16661 VGND.t3565 VGND.t1665 369.318
R16662 VGND.t4221 VGND.t5463 369.318
R16663 VGND.t6347 VGND.t2939 369.318
R16664 VGND.t6345 VGND 369.318
R16665 VGND.t5050 VGND.t6012 369.318
R16666 VGND.t5048 VGND.t6010 369.318
R16667 VGND.t5044 VGND.t6014 369.318
R16668 VGND.t6426 VGND.t218 369.318
R16669 VGND.t187 VGND.t4063 369.318
R16670 VGND VGND.t3118 369.318
R16671 VGND VGND.t5590 369.318
R16672 VGND.t5392 VGND 369.318
R16673 VGND.t2056 VGND.t4962 369.318
R16674 VGND.t6106 VGND.t6545 369.318
R16675 VGND.t4413 VGND.n1721 369.318
R16676 VGND VGND.t6027 369.318
R16677 VGND.t871 VGND.t6532 369.318
R16678 VGND.t3795 VGND 369.318
R16679 VGND.t258 VGND.t6416 369.318
R16680 VGND VGND.t1829 369.318
R16681 VGND VGND.t2469 369.318
R16682 VGND.t6357 VGND.t6375 369.318
R16683 VGND.t6733 VGND.t160 369.318
R16684 VGND.t5757 VGND.t2096 369.318
R16685 VGND.t128 VGND.t6780 369.318
R16686 VGND.t1809 VGND 369.318
R16687 VGND.t6685 VGND.t3265 364.702
R16688 VGND.t6228 VGND.t4092 364.702
R16689 VGND.t5622 VGND.t2697 364.702
R16690 VGND.t202 VGND.t5355 364.702
R16691 VGND.t3940 VGND 360.086
R16692 VGND VGND.t1143 360.086
R16693 VGND.t2780 VGND 360.086
R16694 VGND.t3355 VGND 360.086
R16695 VGND.t5776 VGND.t2359 360.086
R16696 VGND.t897 VGND.t2305 360.086
R16697 VGND VGND.t897 360.086
R16698 VGND.t5034 VGND.t2277 360.086
R16699 VGND.t1601 VGND 360.086
R16700 VGND VGND.t2021 360.086
R16701 VGND VGND.t4563 360.086
R16702 VGND.t3824 VGND 360.086
R16703 VGND.t3623 VGND.t1448 360.086
R16704 VGND.t1448 VGND 360.086
R16705 VGND VGND.t5148 360.086
R16706 VGND.t1452 VGND 360.086
R16707 VGND.t4970 VGND.t3453 360.086
R16708 VGND.t5081 VGND.t4495 360.086
R16709 VGND.t6047 VGND.t3652 360.086
R16710 VGND VGND.t6047 360.086
R16711 VGND.t738 VGND 360.086
R16712 VGND VGND.t3313 360.086
R16713 VGND.t2213 VGND.t5027 360.086
R16714 VGND.t2733 VGND.t5141 360.086
R16715 VGND VGND.t2733 360.086
R16716 VGND.t1631 VGND.t2386 360.086
R16717 VGND.t3275 VGND 360.086
R16718 VGND.t4520 VGND.t5257 360.086
R16719 VGND VGND.t6568 355.469
R16720 VGND VGND.t6228 355.469
R16721 VGND.t6655 VGND.t3377 350.853
R16722 VGND.t6657 VGND.t3379 350.853
R16723 VGND.t3482 VGND.t1099 350.853
R16724 VGND.t2221 VGND.t5416 350.853
R16725 VGND VGND.t4283 350.853
R16726 VGND VGND.t6689 350.853
R16727 VGND.t470 VGND.t5691 350.853
R16728 VGND.t1038 VGND 350.853
R16729 VGND.t4051 VGND.t6675 350.853
R16730 VGND VGND.t1190 350.853
R16731 VGND.t1187 VGND.t278 350.853
R16732 VGND.t6430 VGND.t280 350.853
R16733 VGND.t6502 VGND.t276 350.853
R16734 VGND.t3794 VGND.t24 350.853
R16735 VGND.t858 VGND.t2799 350.853
R16736 VGND.t4857 VGND.t3404 350.853
R16737 VGND.t877 VGND.t162 350.853
R16738 VGND.t4981 VGND.t3039 350.853
R16739 VGND.t6509 VGND 350.853
R16740 VGND.t6506 VGND 350.853
R16741 VGND.t4895 VGND.t6320 347.738
R16742 VGND.t587 VGND.t232 346.236
R16743 VGND.t5411 VGND.t2479 341.62
R16744 VGND.t5413 VGND.t2477 341.62
R16745 VGND.t2015 VGND.t1068 341.62
R16746 VGND.t2017 VGND.t1070 341.62
R16747 VGND.t2721 VGND.t3279 341.62
R16748 VGND.t2723 VGND.t3281 341.62
R16749 VGND.t4788 VGND.t2245 338.82
R16750 VGND.t5600 VGND.t6442 337.003
R16751 VGND.t4163 VGND.t1910 337.003
R16752 VGND.t6648 VGND.t252 335.373
R16753 VGND.n1370 VGND.t6428 332.387
R16754 VGND.t1945 VGND 332.387
R16755 VGND.t5209 VGND.t3748 332.387
R16756 VGND.t4168 VGND.t3413 332.387
R16757 VGND.t5531 VGND.n840 332.387
R16758 VGND.t2610 VGND.t3311 332.387
R16759 VGND.t1348 VGND.t3113 332.387
R16760 VGND.t1350 VGND.t6057 332.387
R16761 VGND.n1448 VGND.t3688 332.387
R16762 VGND VGND.t2865 332.387
R16763 VGND.t803 VGND 332.387
R16764 VGND.t6229 VGND.t1785 332.387
R16765 VGND.t954 VGND.t3185 332.387
R16766 VGND.t391 VGND.t3060 332.387
R16767 VGND.t4121 VGND.n1202 332.387
R16768 VGND.t4874 VGND.t2467 332.387
R16769 VGND.t477 VGND.t2590 332.387
R16770 VGND.t705 VGND.t1505 332.387
R16771 VGND.n798 VGND.t4279 332.387
R16772 VGND.t3107 VGND.t6460 332.387
R16773 VGND VGND.t6267 332.387
R16774 VGND.t4936 VGND.t4532 332.387
R16775 VGND.t6798 VGND.t5656 332.387
R16776 VGND.t3995 VGND.t204 332.387
R16777 VGND.t3728 VGND 332.387
R16778 VGND.t5995 VGND.t32 332.387
R16779 VGND.t5059 VGND.t6706 332.387
R16780 VGND.t749 VGND.t1034 332.387
R16781 VGND.t3436 VGND.t1470 332.387
R16782 VGND.t3269 VGND.t1772 332.387
R16783 VGND.t2619 VGND.t5982 332.387
R16784 VGND.t5585 VGND.t1509 332.387
R16785 VGND VGND.t268 332.387
R16786 VGND VGND.t1919 332.387
R16787 VGND.t151 VGND.t3884 332.387
R16788 VGND VGND.t2642 332.387
R16789 VGND.t4737 VGND.t6222 332.387
R16790 VGND.t6670 VGND.t1516 332.387
R16791 VGND.t3202 VGND.t1585 332.387
R16792 VGND.t2473 VGND.n577 332.387
R16793 VGND.t3828 VGND.t3100 332.387
R16794 VGND.n625 VGND.t4992 332.387
R16795 VGND VGND.t6618 332.387
R16796 VGND.t1420 VGND.t2140 332.387
R16797 VGND.n2206 VGND.t6571 332.387
R16798 VGND.t5500 VGND 332.387
R16799 VGND.n2223 VGND.t3422 332.387
R16800 VGND.t1518 VGND.t944 332.387
R16801 VGND.n555 VGND.t6516 332.387
R16802 VGND.t3200 VGND.t5904 332.387
R16803 VGND.t2451 VGND.t5582 332.387
R16804 VGND.t4395 VGND.t6363 332.387
R16805 VGND.t4433 VGND.t1428 332.387
R16806 VGND.t1651 VGND.t543 332.387
R16807 VGND.n572 VGND.t5012 332.387
R16808 VGND.t4312 VGND.t2901 332.387
R16809 VGND VGND.t3983 332.387
R16810 VGND.t6420 VGND.n560 332.387
R16811 VGND.t6307 VGND.t4841 327.771
R16812 VGND.t3740 VGND.t3736 323.154
R16813 VGND.t1536 VGND 323.154
R16814 VGND.t4162 VGND.t179 323.154
R16815 VGND.t6218 VGND.t6537 320.988
R16816 VGND.t4644 VGND.t757 318.538
R16817 VGND.t5906 VGND 313.921
R16818 VGND.t1237 VGND 313.921
R16819 VGND VGND.n895 313.921
R16820 VGND VGND.t4112 313.921
R16821 VGND VGND.t5696 313.921
R16822 VGND.n1360 VGND.t2838 313.921
R16823 VGND.n1245 VGND 313.921
R16824 VGND VGND.t5459 313.921
R16825 VGND VGND.t2765 313.921
R16826 VGND.t3608 VGND 313.921
R16827 VGND.t5260 VGND 313.921
R16828 VGND VGND.t5260 313.921
R16829 VGND.t3271 VGND 313.921
R16830 VGND VGND.t5566 313.921
R16831 VGND VGND.t1563 313.921
R16832 VGND.t4229 VGND.t6071 313.921
R16833 VGND VGND.t4601 313.921
R16834 VGND VGND.t901 313.921
R16835 VGND VGND.t676 313.921
R16836 VGND.t4391 VGND 313.921
R16837 VGND VGND.n771 313.921
R16838 VGND.n771 VGND 313.921
R16839 VGND VGND.t3820 313.921
R16840 VGND.t2827 VGND.t168 313.921
R16841 VGND.t1241 VGND.t541 313.921
R16842 VGND.t1188 VGND.t123 313.921
R16843 VGND.t282 VGND.t10 313.921
R16844 VGND.t6131 VGND.t5191 313.921
R16845 VGND.t5445 VGND.t1373 313.921
R16846 VGND.t6119 VGND.t692 313.921
R16847 VGND.t2972 VGND.t2810 313.921
R16848 VGND.t5262 VGND 313.921
R16849 VGND VGND.t4694 313.921
R16850 VGND.t4989 VGND 313.921
R16851 VGND VGND.t5508 313.921
R16852 VGND.t5619 VGND 313.921
R16853 VGND.t5818 VGND 313.921
R16854 VGND.t5492 VGND.t5302 313.921
R16855 VGND.t358 VGND 313.921
R16856 VGND.t3900 VGND 313.921
R16857 VGND.t4265 VGND 313.921
R16858 VGND.t6043 VGND 313.921
R16859 VGND VGND.t5723 313.921
R16860 VGND VGND.t5159 313.921
R16861 VGND VGND.t1234 313.921
R16862 VGND.t1377 VGND.t5368 313.921
R16863 VGND.t5083 VGND.t6157 313.921
R16864 VGND.t2108 VGND 313.921
R16865 VGND.t2855 VGND 313.921
R16866 VGND VGND.t3068 313.921
R16867 VGND.n2631 VGND 313.921
R16868 VGND.n2633 VGND 313.921
R16869 VGND.n2092 VGND 313.921
R16870 VGND.t5417 VGND 313.921
R16871 VGND.t1671 VGND.t2449 313.921
R16872 VGND.n2095 VGND 313.921
R16873 VGND VGND.n358 313.921
R16874 VGND VGND.n1021 313.921
R16875 VGND.n1023 VGND 313.921
R16876 VGND.n1023 VGND 313.921
R16877 VGND VGND.t5986 313.921
R16878 VGND VGND.t5389 313.921
R16879 VGND VGND.t1669 313.921
R16880 VGND.t1669 VGND 313.921
R16881 VGND.t5753 VGND 313.921
R16882 VGND.t2998 VGND 313.921
R16883 VGND.t684 VGND 313.921
R16884 VGND.t1109 VGND 313.921
R16885 VGND.t2532 VGND 313.921
R16886 VGND.t4632 VGND 313.921
R16887 VGND VGND.t2793 313.921
R16888 VGND.t1645 VGND 313.921
R16889 VGND.t5628 VGND 313.921
R16890 VGND.t2578 VGND 313.921
R16891 VGND VGND.t3402 313.921
R16892 VGND.t747 VGND 313.921
R16893 VGND.t4389 VGND 313.921
R16894 VGND.t1993 VGND 313.921
R16895 VGND VGND.t3292 313.921
R16896 VGND.t519 VGND 313.921
R16897 VGND.t829 VGND 313.921
R16898 VGND.t1045 VGND 313.921
R16899 VGND.t5311 VGND 313.921
R16900 VGND.t5761 VGND 313.921
R16901 VGND.t2379 VGND.t6646 312.072
R16902 VGND VGND.t3201 309.305
R16903 VGND VGND.t1536 304.688
R16904 VGND.t177 VGND.t526 300.072
R16905 VGND.t4414 VGND.t6341 300.072
R16906 VGND.t6591 VGND.t6392 295.455
R16907 VGND.t778 VGND.t4365 295.455
R16908 VGND.t6726 VGND.t1572 295.455
R16909 VGND.t1544 VGND 295.455
R16910 VGND.t2865 VGND 295.455
R16911 VGND.t6259 VGND.t6251 295.455
R16912 VGND.t1925 VGND.t3330 295.455
R16913 VGND.t6279 VGND.t5169 295.455
R16914 VGND.t6269 VGND.t3135 295.455
R16915 VGND.t6265 VGND.t6098 295.455
R16916 VGND VGND.t3149 295.455
R16917 VGND.t242 VGND 295.455
R16918 VGND.t268 VGND 295.455
R16919 VGND.t1064 VGND.n478 295.455
R16920 VGND.t583 VGND 295.455
R16921 VGND VGND.t5500 295.455
R16922 VGND.t6367 VGND.t6730 295.455
R16923 VGND.t158 VGND.t6369 295.455
R16924 VGND.n522 VGND.t2502 295.455
R16925 VGND.t3983 VGND 295.455
R16926 VGND.t3676 VGND.t3224 290.839
R16927 VGND.t3467 VGND.t3590 290.839
R16928 VGND.t6696 VGND.t1011 286.223
R16929 VGND.t4839 VGND 286.223
R16930 VGND.t4979 VGND 285.322
R16931 VGND.t6231 VGND 285.322
R16932 VGND.t6236 VGND 285.322
R16933 VGND.t4527 VGND.t3478 285.322
R16934 VGND.t4534 VGND.t6031 285.322
R16935 VGND.t29 VGND.t175 285.322
R16936 VGND.t4526 VGND.t2419 281.606
R16937 VGND.t6151 VGND.t5394 281.606
R16938 VGND.t3201 VGND.t6308 281.606
R16939 VGND.t5530 VGND 276.99
R16940 VGND.t4066 VGND.t2869 276.99
R16941 VGND.t6538 VGND.t2894 276.99
R16942 VGND.t609 VGND.t6200 276.99
R16943 VGND VGND.t6099 276.99
R16944 VGND.t1190 VGND 276.99
R16945 VGND.t6359 VGND.t5474 276.99
R16946 VGND.t5785 VGND.t6323 276.99
R16947 VGND.t2604 VGND.t303 276.99
R16948 VGND.t2031 VGND.t210 276.99
R16949 VGND.t3860 VGND.t2453 276.99
R16950 VGND.t1483 VGND.t6383 272.373
R16951 VGND.t1410 VGND.t4961 272.373
R16952 VGND.t5747 VGND.t2664 267.757
R16953 VGND.t3681 VGND 267.757
R16954 VGND.t568 VGND.t5510 263.139
R16955 VGND.t3519 VGND.n278 258.524
R16956 VGND.t4897 VGND.n152 258.524
R16957 VGND.t4978 VGND.t90 258.524
R16958 VGND VGND.t6345 258.524
R16959 VGND VGND.t1949 258.524
R16960 VGND.t3738 VGND.t5530 258.524
R16961 VGND.t3226 VGND 258.524
R16962 VGND VGND.t3226 258.524
R16963 VGND.t5590 VGND 258.524
R16964 VGND.t2238 VGND.t6258 258.524
R16965 VGND VGND.t609 258.524
R16966 VGND.n250 VGND.t1270 258.524
R16967 VGND.t5394 VGND 258.524
R16968 VGND VGND.t5392 258.524
R16969 VGND.t3923 VGND.n1725 258.524
R16970 VGND VGND.t5630 258.524
R16971 VGND.t5615 VGND.t2144 258.524
R16972 VGND.t1589 VGND.t3440 258.524
R16973 VGND.t5474 VGND 258.524
R16974 VGND.t3002 VGND.t707 258.524
R16975 VGND VGND.t2644 258.524
R16976 VGND VGND.t5785 258.524
R16977 VGND.t4586 VGND.t2337 258.524
R16978 VGND.t1829 VGND 258.524
R16979 VGND VGND.t6000 258.524
R16980 VGND VGND.t1809 258.524
R16981 VGND.t6573 VGND.t4839 253.906
R16982 VGND.t4306 VGND.t4530 253.906
R16983 VGND.t304 VGND.t4159 253.906
R16984 VGND.t2812 VGND.t6637 249.291
R16985 VGND.t1609 VGND.t1544 240.058
R16986 VGND.t3330 VGND 240.058
R16987 VGND.t6396 VGND.t1595 240.058
R16988 VGND.t6263 VGND.t2153 240.058
R16989 VGND.t3956 VGND.t5391 240.058
R16990 VGND.t466 VGND.t3730 240.058
R16991 VGND.t4844 VGND.t6596 240.058
R16992 VGND.t6448 VGND.t4416 240.058
R16993 VGND.t4418 VGND.t2537 240.058
R16994 VGND.t5244 VGND.t4647 240.058
R16995 VGND.t585 VGND.t6500 240.058
R16996 VGND.t6730 VGND 240.058
R16997 VGND VGND.t158 240.058
R16998 VGND.t1514 VGND.t216 240.058
R16999 VGND.t5808 VGND.t5788 235.44
R17000 VGND.t4002 VGND.t769 235.44
R17001 VGND.t6256 VGND.t4497 231.825
R17002 VGND.t4536 VGND.t3954 231.825
R17003 VGND.t6661 VGND.t6291 226.208
R17004 VGND.t4412 VGND.t165 226.208
R17005 VGND.t4729 VGND.t3935 221.591
R17006 VGND.t2428 VGND.t3936 221.591
R17007 VGND.t4231 VGND.t2505 221.591
R17008 VGND.t1787 VGND.t2596 221.591
R17009 VGND.t5182 VGND.t2807 221.591
R17010 VGND.t990 VGND.t450 221.591
R17011 VGND.n794 VGND.t5091 221.591
R17012 VGND.t6138 VGND.t454 221.591
R17013 VGND.t4781 VGND.t2448 221.591
R17014 VGND.t123 VGND 221.591
R17015 VGND VGND.t282 221.591
R17016 VGND VGND.t6635 221.591
R17017 VGND.t6612 VGND.t238 221.591
R17018 VGND.t6598 VGND.t240 221.591
R17019 VGND.t3639 VGND.t515 221.591
R17020 VGND VGND.t1383 221.591
R17021 VGND.t2559 VGND 221.591
R17022 VGND.t82 VGND.t2571 221.591
R17023 VGND VGND.t5083 221.591
R17024 VGND.t6691 VGND.t4119 216.975
R17025 VGND VGND.t4979 213.993
R17026 VGND.t5427 VGND.t2331 207.742
R17027 VGND.t1266 VGND 203.125
R17028 VGND VGND.t4544 203.125
R17029 VGND VGND.t1456 203.125
R17030 VGND.t6806 VGND 203.125
R17031 VGND VGND.t3654 203.125
R17032 VGND VGND.t5282 203.125
R17033 VGND VGND.t2088 203.125
R17034 VGND VGND.t6755 203.125
R17035 VGND VGND.t4261 203.125
R17036 VGND VGND.t517 203.125
R17037 VGND VGND.t1230 203.125
R17038 VGND VGND.t1873 203.125
R17039 VGND VGND.t3450 203.125
R17040 VGND.t4061 VGND 203.125
R17041 VGND VGND.t3686 203.125
R17042 VGND VGND.n43 203.125
R17043 VGND.t5928 VGND 203.125
R17044 VGND.t1618 VGND 203.125
R17045 VGND.t2737 VGND 203.125
R17046 VGND.t4269 VGND 203.125
R17047 VGND.n894 VGND 203.125
R17048 VGND.t4028 VGND.t298 203.125
R17049 VGND.t6778 VGND.t4030 203.125
R17050 VGND.t6220 VGND.t4032 203.125
R17051 VGND.t6441 VGND.t6240 203.125
R17052 VGND.t3894 VGND.t5698 203.125
R17053 VGND VGND.t5209 203.125
R17054 VGND VGND.t4819 203.125
R17055 VGND VGND.t3290 203.125
R17056 VGND VGND.t1777 203.125
R17057 VGND.t3311 VGND 203.125
R17058 VGND.t3113 VGND 203.125
R17059 VGND.t4528 VGND.t525 203.125
R17060 VGND.n1448 VGND 203.125
R17061 VGND.t5760 VGND.t5219 203.125
R17062 VGND.t229 VGND.t5305 203.125
R17063 VGND.t527 VGND.t5007 203.125
R17064 VGND.t36 VGND.t3026 203.125
R17065 VGND.t3185 VGND 203.125
R17066 VGND.t3262 VGND.t6112 203.125
R17067 VGND.t5350 VGND.t929 203.125
R17068 VGND.t5423 VGND.t4331 203.125
R17069 VGND.n1202 VGND 203.125
R17070 VGND VGND.t477 203.125
R17071 VGND VGND.n798 203.125
R17072 VGND VGND.t3107 203.125
R17073 VGND VGND.t6798 203.125
R17074 VGND.t5690 VGND.n1716 203.125
R17075 VGND VGND.t1553 203.125
R17076 VGND.t4049 VGND.t167 203.125
R17077 VGND.t5632 VGND.t6385 203.125
R17078 VGND VGND.t5835 203.125
R17079 VGND.t5307 VGND.t4670 203.125
R17080 VGND VGND.t749 203.125
R17081 VGND.t1470 VGND 203.125
R17082 VGND VGND.t3269 203.125
R17083 VGND.t1766 VGND.t2273 203.125
R17084 VGND VGND.t2619 203.125
R17085 VGND VGND.t5585 203.125
R17086 VGND.t5223 VGND 203.125
R17087 VGND.t5385 VGND.t6528 203.125
R17088 VGND.t2489 VGND.t1813 203.125
R17089 VGND VGND.t4737 203.125
R17090 VGND VGND.t436 203.125
R17091 VGND VGND.t2485 203.125
R17092 VGND.t1585 VGND 203.125
R17093 VGND VGND.t4287 203.125
R17094 VGND VGND.t4676 203.125
R17095 VGND VGND.t3841 203.125
R17096 VGND VGND.t3347 203.125
R17097 VGND.t5294 VGND 203.125
R17098 VGND VGND.n577 203.125
R17099 VGND.n583 VGND.t23 203.125
R17100 VGND VGND.t4674 203.125
R17101 VGND VGND.t1639 203.125
R17102 VGND.t2140 VGND 203.125
R17103 VGND VGND.t772 203.125
R17104 VGND VGND.t4542 203.125
R17105 VGND.t5243 VGND.n472 203.125
R17106 VGND.t4652 VGND.t2757 203.125
R17107 VGND.t131 VGND.t2759 203.125
R17108 VGND.t3250 VGND.t6191 203.125
R17109 VGND VGND.t6164 203.125
R17110 VGND VGND.t75 203.125
R17111 VGND.t1637 VGND 203.125
R17112 VGND VGND.t4489 203.125
R17113 VGND VGND.t3387 203.125
R17114 VGND VGND.t575 203.125
R17115 VGND.t5733 VGND.t678 203.125
R17116 VGND VGND.t6166 203.125
R17117 VGND VGND.t4469 203.125
R17118 VGND.n2223 VGND 203.125
R17119 VGND.t5225 VGND 203.125
R17120 VGND.t2634 VGND 203.125
R17121 VGND.t6765 VGND 203.125
R17122 VGND.t940 VGND 203.125
R17123 VGND.t1124 VGND 203.125
R17124 VGND.t2791 VGND 203.125
R17125 VGND VGND.t4114 203.125
R17126 VGND VGND.n2493 203.125
R17127 VGND VGND.n2494 203.125
R17128 VGND VGND.t1518 203.125
R17129 VGND.t3172 VGND 203.125
R17130 VGND.t4710 VGND 203.125
R17131 VGND VGND.t5010 203.125
R17132 VGND VGND.t5074 203.125
R17133 VGND VGND.t4763 203.125
R17134 VGND.t3398 VGND 203.125
R17135 VGND VGND.t1388 203.125
R17136 VGND VGND.t462 203.125
R17137 VGND VGND.t3187 203.125
R17138 VGND VGND.t5144 203.125
R17139 VGND.n2634 VGND 203.125
R17140 VGND VGND.t4999 203.125
R17141 VGND VGND.t4292 203.125
R17142 VGND.t589 VGND 203.125
R17143 VGND.t5437 VGND 203.125
R17144 VGND VGND.t1480 203.125
R17145 VGND VGND.t1542 203.125
R17146 VGND VGND.n555 203.125
R17147 VGND.n554 VGND 203.125
R17148 VGND.t485 VGND 203.125
R17149 VGND.t5904 VGND 203.125
R17150 VGND.t5582 VGND 203.125
R17151 VGND VGND.t4395 203.125
R17152 VGND VGND.t3050 203.125
R17153 VGND.t1390 VGND 203.125
R17154 VGND.n357 VGND 203.125
R17155 VGND.t993 VGND 203.125
R17156 VGND VGND.t4433 203.125
R17157 VGND.t543 VGND 203.125
R17158 VGND.t5607 VGND.t3833 203.125
R17159 VGND.t1869 VGND 203.125
R17160 VGND VGND.n572 203.125
R17161 VGND.t2901 VGND 203.125
R17162 VGND.n567 VGND.t4650 203.125
R17163 VGND.n560 VGND 203.125
R17164 VGND.n3313 VGND 203.125
R17165 VGND VGND.n6 203.125
R17166 VGND.t2382 VGND.t6567 198.51
R17167 VGND.t725 VGND.t1114 198.51
R17168 VGND.t87 VGND.t6235 196.16
R17169 VGND.t6214 VGND.t6232 196.16
R17170 VGND.t6723 VGND.t256 196.16
R17171 VGND.t9 VGND.t254 196.16
R17172 VGND.t8 VGND.t250 196.16
R17173 VGND.t6716 VGND.t266 196.16
R17174 VGND.t288 VGND.t1700 193.893
R17175 VGND.t6300 VGND.t6153 193.893
R17176 VGND.t6562 VGND 189.276
R17177 VGND.t6547 VGND.t4673 189.276
R17178 VGND.t2920 VGND.t6212 184.66
R17179 VGND.t2132 VGND.t3168 184.66
R17180 VGND.t3548 VGND.t2516 184.66
R17181 VGND.t2394 VGND.t2522 184.66
R17182 VGND.n1348 VGND.t4885 184.66
R17183 VGND.t5036 VGND.t2629 184.66
R17184 VGND.n1354 VGND.t1424 184.66
R17185 VGND.t6036 VGND.t789 184.66
R17186 VGND VGND.t1945 184.66
R17187 VGND VGND.t1947 184.66
R17188 VGND.t343 VGND.t768 184.66
R17189 VGND.t5284 VGND.t3886 184.66
R17190 VGND.t3658 VGND.t4686 184.66
R17191 VGND.t6373 VGND.t5865 184.66
R17192 VGND.t6353 VGND.t5016 184.66
R17193 VGND VGND.t6298 184.66
R17194 VGND.t3424 VGND.t163 184.66
R17195 VGND.t3475 VGND.t399 184.66
R17196 VGND.t5694 VGND.t6113 184.66
R17197 VGND.t6687 VGND.t2459 184.66
R17198 VGND.t432 VGND.t4275 184.66
R17199 VGND.t6283 VGND.t112 184.66
R17200 VGND.t6267 VGND 184.66
R17201 VGND.t473 VGND.t1038 184.66
R17202 VGND VGND.t4051 184.66
R17203 VGND.t6475 VGND.t680 184.66
R17204 VGND.t599 VGND.t6193 184.66
R17205 VGND.t2907 VGND.t2703 184.66
R17206 VGND.t5868 VGND.t913 184.66
R17207 VGND.t278 VGND 184.66
R17208 VGND.t6115 VGND.n1823 184.66
R17209 VGND.t2271 VGND.t4325 184.66
R17210 VGND.t6365 VGND.t581 184.66
R17211 VGND.n1076 VGND.t2958 184.66
R17212 VGND.t55 VGND.t3991 184.66
R17213 VGND.t5121 VGND.t505 184.66
R17214 VGND.t856 VGND.t6309 184.66
R17215 VGND.t6440 VGND.t244 184.66
R17216 VGND.n944 VGND.t6452 184.66
R17217 VGND.t5370 VGND.t2677 184.66
R17218 VGND.t5238 VGND.t5719 184.66
R17219 VGND.t6377 VGND.t2316 184.66
R17220 VGND.t3862 VGND.t2247 184.66
R17221 VGND.t40 VGND.n2093 184.66
R17222 VGND.t509 VGND.n1022 184.66
R17223 VGND.n570 VGND.t3785 184.66
R17224 VGND.t2149 VGND.t185 184.66
R17225 VGND.t4505 VGND.t6331 184.66
R17226 VGND VGND.t4856 184.66
R17227 VGND.t6568 VGND.t1811 180.043
R17228 VGND.t1013 VGND.t3022 180.043
R17229 VGND.t4538 VGND.t4067 180.043
R17230 VGND VGND.t5383 180.043
R17231 VGND.n289 VGND.t6137 178.327
R17232 VGND.t6740 VGND.t3335 175.427
R17233 VGND.t1143 VGND.t2778 175.427
R17234 VGND.t1145 VGND.t2780 175.427
R17235 VGND.t2979 VGND.t6237 175.427
R17236 VGND.t2983 VGND.t6247 175.427
R17237 VGND.t2981 VGND.t5700 175.427
R17238 VGND.t2019 VGND.t1601 175.427
R17239 VGND.t2021 VGND.t1603 175.427
R17240 VGND.t4563 VGND.t3822 175.427
R17241 VGND.t4565 VGND.t3824 175.427
R17242 VGND.t429 VGND.t4855 175.427
R17243 VGND.t5148 VGND.t1450 175.427
R17244 VGND.t5146 VGND.t1452 175.427
R17245 VGND.t3315 VGND.t738 175.427
R17246 VGND.t3313 VGND.t740 175.427
R17247 VGND.t1255 VGND.t1538 170.81
R17248 VGND.t3784 VGND.t1216 170.81
R17249 VGND.t6394 VGND.t2120 166.194
R17250 VGND.t946 VGND 166.194
R17251 VGND.t3118 VGND.t5645 166.194
R17252 VGND VGND.t227 166.194
R17253 VGND.t225 VGND.t5592 166.194
R17254 VGND.t6492 VGND.t6254 166.194
R17255 VGND.t6293 VGND.t952 166.194
R17256 VGND VGND.t389 166.194
R17257 VGND.t6276 VGND.t12 166.194
R17258 VGND.t6271 VGND.t110 166.194
R17259 VGND.t5217 VGND.t3155 166.194
R17260 VGND.t1587 VGND.t5031 166.194
R17261 VGND.t1812 VGND.n726 166.194
R17262 VGND.t6050 VGND.t4809 166.194
R17263 VGND.t5597 VGND.t6321 166.194
R17264 VGND.t6456 VGND.t3795 166.194
R17265 VGND.t4077 VGND.t4859 166.194
R17266 VGND VGND.t4651 166.194
R17267 VGND VGND.t5781 166.194
R17268 VGND.t6644 VGND.t5156 166.194
R17269 VGND.t193 VGND 166.194
R17270 VGND VGND.t6509 166.194
R17271 VGND VGND.t1076 161.577
R17272 VGND.t460 VGND.t3147 161.577
R17273 VGND.t5542 VGND.t4570 160.672
R17274 VGND.t4570 VGND.t5973 160.672
R17275 VGND.t5973 VGND.t1148 160.672
R17276 VGND.t1148 VGND.t4106 160.672
R17277 VGND.t4047 VGND.t1381 160.672
R17278 VGND.t1381 VGND.t3931 160.672
R17279 VGND.t3931 VGND.t1097 160.672
R17280 VGND.t6020 VGND.t3219 160.672
R17281 VGND.t3219 VGND.t5815 160.672
R17282 VGND.t5815 VGND.t2658 160.672
R17283 VGND.t5018 VGND.t4321 160.672
R17284 VGND.t5079 VGND.t5018 160.672
R17285 VGND.t5251 VGND.t5079 160.672
R17286 VGND.t3554 VGND.t5251 160.672
R17287 VGND.t6536 VGND 160.494
R17288 VGND.t1663 VGND 156.96
R17289 VGND VGND.t3567 156.96
R17290 VGND.t5461 VGND 156.96
R17291 VGND VGND.t4223 156.96
R17292 VGND.n891 VGND.t1860 156.96
R17293 VGND.t3709 VGND.t881 156.96
R17294 VGND.t4117 VGND 156.96
R17295 VGND.t4684 VGND.t1622 156.96
R17296 VGND.t5912 VGND.t5025 156.96
R17297 VGND.t1607 VGND.n1123 156.96
R17298 VGND.t274 VGND.t4836 156.96
R17299 VGND.t2956 VGND 156.96
R17300 VGND.t3989 VGND 156.96
R17301 VGND.t1001 VGND.t5896 156.96
R17302 VGND.t1655 VGND.t2890 156.96
R17303 VGND VGND.t5163 156.96
R17304 VGND.t2475 VGND 156.96
R17305 VGND.t5721 VGND 156.96
R17306 VGND.t2100 VGND.t5624 156.96
R17307 VGND VGND.t5755 156.96
R17308 VGND.t2098 VGND 156.96
R17309 VGND.t4974 VGND 156.96
R17310 VGND.t3420 VGND.t4480 156.96
R17311 VGND VGND.t5743 156.96
R17312 VGND.t2249 VGND 156.96
R17313 VGND.n573 VGND.t2725 156.96
R17314 VGND.t5056 VGND.t3684 152.345
R17315 VGND.n1349 VGND.t6507 152.345
R17316 VGND.t4068 VGND.t1783 152.345
R17317 VGND.t5131 VGND.t1015 152.345
R17318 VGND.t3770 VGND.t3679 152.345
R17319 VGND.t1182 VGND.t1178 147.727
R17320 VGND VGND.t5790 147.727
R17321 VGND.t4848 VGND.t6679 147.727
R17322 VGND.t2130 VGND.t317 147.727
R17323 VGND.t6744 VGND.t3530 147.727
R17324 VGND.t3972 VGND 147.727
R17325 VGND.t6724 VGND.t3690 147.727
R17326 VGND.t1927 VGND.t468 147.727
R17327 VGND.t6488 VGND.t6790 147.727
R17328 VGND.t1929 VGND.t106 147.727
R17329 VGND.t3480 VGND.t100 147.727
R17330 VGND.t393 VGND.t3303 147.727
R17331 VGND.t6701 VGND.t1028 147.727
R17332 VGND.t6274 VGND.t3134 147.727
R17333 VGND.t6032 VGND 147.727
R17334 VGND.t3767 VGND.t479 147.727
R17335 VGND.t5954 VGND.t30 147.727
R17336 VGND.t4264 VGND 147.727
R17337 VGND.t6524 VGND.t869 147.727
R17338 VGND VGND.t3698 147.727
R17339 VGND.t234 VGND.t6622 147.727
R17340 VGND.t236 VGND.t6614 147.727
R17341 VGND VGND.t1218 147.727
R17342 VGND.t5570 VGND.t2861 147.727
R17343 VGND.t135 VGND.t2761 147.727
R17344 VGND.t223 VGND.t6518 147.727
R17345 VGND.t221 VGND.t85 147.727
R17346 VGND.t3788 VGND.t44 147.727
R17347 VGND.t2962 VGND.t4459 147.727
R17348 VGND.t1807 VGND.t4994 147.727
R17349 VGND.t6424 VGND.t6361 147.727
R17350 VGND.t4671 VGND.t950 143.112
R17351 VGND.t915 VGND.t1404 143.112
R17352 VGND.t6556 VGND.t6140 142.661
R17353 VGND.t6348 VGND.t4722 133.879
R17354 VGND VGND.t3677 133.879
R17355 VGND.t4198 VGND 133.879
R17356 VGND.t190 VGND.t4310 133.879
R17357 VGND VGND.t3937 129.262
R17358 VGND.t1464 VGND 129.262
R17359 VGND.t1858 VGND 129.262
R17360 VGND VGND.t2045 129.262
R17361 VGND.t6016 VGND 129.262
R17362 VGND VGND.t5046 129.262
R17363 VGND.t195 VGND 129.262
R17364 VGND.t6438 VGND 129.262
R17365 VGND.t6721 VGND 129.262
R17366 VGND.t6739 VGND.t6250 129.262
R17367 VGND VGND.t5533 129.262
R17368 VGND VGND.t6695 129.262
R17369 VGND VGND.t888 129.262
R17370 VGND.t6463 VGND.t6431 129.262
R17371 VGND.t212 VGND.t6326 129.262
R17372 VGND.t6549 VGND.t5297 129.262
R17373 VGND.t6539 VGND 129.262
R17374 VGND.t883 VGND 129.262
R17375 VGND VGND.t4561 129.262
R17376 VGND VGND.t4682 129.262
R17377 VGND.t759 VGND 129.262
R17378 VGND VGND.t200 129.262
R17379 VGND.t6668 VGND.t4688 129.262
R17380 VGND.t6472 VGND.t4053 129.262
R17381 VGND.t6028 VGND.t4054 129.262
R17382 VGND VGND.t6208 129.262
R17383 VGND.t2815 VGND 129.262
R17384 VGND VGND.t5914 129.262
R17385 VGND.t6784 VGND 129.262
R17386 VGND VGND.t1245 129.262
R17387 VGND.t539 VGND 129.262
R17388 VGND.t1696 VGND.t6315 129.262
R17389 VGND.t1212 VGND 129.262
R17390 VGND VGND.t4964 129.262
R17391 VGND.t5605 VGND 129.262
R17392 VGND.t219 VGND.t6108 129.262
R17393 VGND VGND.t2687 129.262
R17394 VGND.t3596 VGND 129.262
R17395 VGND VGND.t5165 129.262
R17396 VGND.t6450 VGND 129.262
R17397 VGND.t4648 VGND 129.262
R17398 VGND VGND.t3630 129.262
R17399 VGND.t181 VGND 129.262
R17400 VGND VGND.t260 129.262
R17401 VGND VGND.t262 129.262
R17402 VGND VGND.t2916 129.262
R17403 VGND.t5300 VGND 129.262
R17404 VGND VGND.t5494 129.262
R17405 VGND.t2914 VGND 129.262
R17406 VGND.t6336 VGND.t921 129.262
R17407 VGND.t2510 VGND.t427 129.262
R17408 VGND.t4317 VGND.t6715 129.262
R17409 VGND.t6025 VGND.t2470 129.262
R17410 VGND.t197 VGND.t1820 129.262
R17411 VGND VGND.t6711 129.262
R17412 VGND.t6189 VGND 129.262
R17413 VGND.t6125 VGND.t5366 129.262
R17414 VGND VGND.t5365 129.262
R17415 VGND.t5264 VGND.t1262 129.262
R17416 VGND.t6123 VGND.t1611 129.262
R17417 VGND VGND.t3015 129.262
R17418 VGND.t5870 VGND 129.262
R17419 VGND VGND.t5741 129.262
R17420 VGND.t2227 VGND.t3858 129.262
R17421 VGND VGND.t4160 129.262
R17422 VGND.t5215 VGND 129.262
R17423 VGND.t1105 VGND.t6141 127.007
R17424 VGND.t3058 VGND.t2945 124.645
R17425 VGND.t6555 VGND.t6666 124.645
R17426 VGND.t6560 VGND.t1147 124.645
R17427 VGND.t6510 VGND.t2413 124.645
R17428 VGND.t5749 VGND.t1975 124.645
R17429 VGND.t3905 VGND.t3556 121.072
R17430 VGND.t3556 VGND.t688 121.072
R17431 VGND.t688 VGND.t438 121.072
R17432 VGND.t438 VGND.t4911 121.072
R17433 VGND.t4911 VGND.t3497 121.072
R17434 VGND.t1335 VGND.t2508 121.072
R17435 VGND.t4887 VGND.t1335 121.072
R17436 VGND.t2705 VGND.t4887 121.072
R17437 VGND.t811 VGND.t2705 121.072
R17438 VGND.t1228 VGND.t811 121.072
R17439 VGND.t5207 VGND.t1228 121.072
R17440 VGND.t5005 VGND.t5207 121.072
R17441 VGND.t307 VGND.t4754 121.072
R17442 VGND.t4235 VGND.t307 121.072
R17443 VGND.t4774 VGND.t4235 121.072
R17444 VGND.t2709 VGND.t4774 121.072
R17445 VGND.t1468 VGND.t2709 121.072
R17446 VGND.t3562 VGND.t1468 121.072
R17447 VGND.t4949 VGND.t3562 121.072
R17448 VGND.t3285 VGND.t3448 121.072
R17449 VGND.t1875 VGND.t3285 121.072
R17450 VGND.t3804 VGND.t1875 121.072
R17451 VGND.t1881 VGND.t3804 121.072
R17452 VGND.t6817 VGND.t1881 121.072
R17453 VGND.t1499 VGND.t6817 121.072
R17454 VGND.t2027 VGND.t1499 121.072
R17455 VGND.n356 VGND.t4047 120.504
R17456 VGND.n3699 VGND.t1097 120.504
R17457 VGND.n3698 VGND.t4321 120.504
R17458 VGND.t6398 VGND.t6540 120.028
R17459 VGND.t1770 VGND.t1026 120.028
R17460 VGND.t3960 VGND.t26 117.934
R17461 VGND.t2875 VGND.t6624 117.934
R17462 VGND VGND.t1688 110.796
R17463 VGND.t6134 VGND.t6558 110.796
R17464 VGND VGND.t2818 110.796
R17465 VGND VGND.t4861 110.796
R17466 VGND VGND.t3267 110.796
R17467 VGND.t5578 VGND.t6281 110.796
R17468 VGND VGND.t6710 110.796
R17469 VGND.t4643 VGND.t6530 110.796
R17470 VGND.t4646 VGND.t6526 110.796
R17471 VGND.n737 VGND.t3773 110.796
R17472 VGND.t3753 VGND 110.796
R17473 VGND.t6110 VGND.t2136 110.796
R17474 VGND VGND.t96 110.796
R17475 VGND.t3829 VGND.t3102 110.796
R17476 VGND.t5621 VGND.t3145 110.796
R17477 VGND VGND.t456 110.796
R17478 VGND.t1264 VGND.t2569 110.796
R17479 VGND.t5502 VGND.t1906 110.796
R17480 VGND VGND.t47 110.796
R17481 VGND.t4864 VGND 110.796
R17482 VGND VGND.t6630 110.796
R17483 VGND.t3023 VGND.t3802 106.18
R17484 VGND.t4073 VGND.t1965 106.18
R17485 VGND.t4893 VGND.t6641 98.0801
R17486 VGND.n2952 VGND.t3905 97.8302
R17487 VGND.t2434 VGND 92.33
R17488 VGND.t6233 VGND.t6338 92.33
R17489 VGND.t5958 VGND 92.33
R17490 VGND.t3325 VGND.t425 92.33
R17491 VGND.t1955 VGND.n665 92.33
R17492 VGND.t5286 VGND 92.33
R17493 VGND.t1745 VGND.n529 92.33
R17494 VGND.t6042 VGND 92.33
R17495 VGND.n2951 VGND.t2508 90.8038
R17496 VGND.t4754 VGND.n2920 90.8038
R17497 VGND.t3448 VGND.n2921 90.8038
R17498 VGND.n3669 VGND.t3554 89.6606
R17499 VGND.t4965 VGND.t6024 87.7136
R17500 VGND.t4980 VGND.t3056 81.6474
R17501 VGND.t6620 VGND.t2874 81.6474
R17502 VGND.t6352 VGND 73.8641
R17503 VGND.t2392 VGND.t6069 73.8641
R17504 VGND.t1161 VGND.t6700 73.8641
R17505 VGND.t6132 VGND.t682 73.8641
R17506 VGND.t3945 VGND.t5506 73.8641
R17507 VGND.t6103 VGND.t3197 73.8641
R17508 VGND.t6301 VGND.t3892 73.8641
R17509 VGND.t6314 VGND 69.2477
R17510 VGND.t2415 VGND.t286 64.6312
R17511 VGND.t1698 VGND.t292 64.6312
R17512 VGND.t4854 VGND.t917 64.6312
R17513 VGND VGND.n356 64.5558
R17514 VGND VGND.n3698 64.5558
R17515 VGND.t6565 VGND.t4703 60.0147
R17516 VGND.t644 VGND.t4151 60.0147
R17517 VGND.t2417 VGND.t3121 60.0147
R17518 VGND.t4106 VGND 55.9484
R17519 VGND.t2658 VGND 55.9484
R17520 VGND.t3375 VGND 55.3982
R17521 VGND.t5435 VGND.t4296 55.3982
R17522 VGND VGND.t664 55.3982
R17523 VGND.t6436 VGND.t2863 55.3982
R17524 VGND.t984 VGND 55.3982
R17525 VGND.t6260 VGND 55.3982
R17526 VGND VGND.t3509 55.3982
R17527 VGND VGND.t387 55.3982
R17528 VGND.t1268 VGND 55.3982
R17529 VGND.n1731 VGND.t3852 55.3982
R17530 VGND.t1102 VGND.t6665 55.3982
R17531 VGND.t2178 VGND 55.3982
R17532 VGND VGND.t327 55.3982
R17533 VGND.t6160 VGND 55.3982
R17534 VGND.t6513 VGND.t4940 55.3982
R17535 VGND.n2922 VGND.n39 52.4286
R17536 VGND VGND.t114 50.7817
R17537 VGND.t2814 VGND.t5255 49.8958
R17538 VGND.n2922 VGND 49.7261
R17539 VGND VGND.n2951 48.6451
R17540 VGND.n2920 VGND 48.6451
R17541 VGND.n2921 VGND 48.6451
R17542 VGND VGND.t3746 46.1653
R17543 VGND VGND.t5908 46.1653
R17544 VGND VGND.t4359 46.1653
R17545 VGND VGND.t1032 46.1653
R17546 VGND VGND.t5662 46.1653
R17547 VGND VGND.t4917 46.1653
R17548 VGND VGND.t2859 46.1653
R17549 VGND.t5572 VGND 46.1653
R17550 VGND.t27 VGND.t2514 45.3599
R17551 VGND.t3497 VGND 42.1592
R17552 VGND VGND.t5005 42.1592
R17553 VGND VGND.t4949 42.1592
R17554 VGND VGND.t2027 42.1592
R17555 VGND.t5523 VGND.t1837 41.5488
R17556 VGND.t6468 VGND.t1532 41.5488
R17557 VGND.t2857 VGND 41.5488
R17558 VGND.t6575 VGND.n659 41.5488
R17559 VGND.t1007 VGND.t3041 41.5488
R17560 VGND.n3699 VGND.t6020 40.1682
R17561 VGND.t2436 VGND.t2437 36.9323
R17562 VGND.t4731 VGND.t3939 36.9323
R17563 VGND VGND.t4909 36.9323
R17564 VGND.t3302 VGND.t2457 36.9323
R17565 VGND.t6535 VGND.t1345 36.9323
R17566 VGND.t6210 VGND.t6659 36.9323
R17567 VGND.t3327 VGND.n144 36.9323
R17568 VGND.t3381 VGND.t6677 36.9323
R17569 VGND.t776 VGND.t89 36.9323
R17570 VGND.t780 VGND.t3138 36.9323
R17571 VGND.t988 VGND.t6329 36.9323
R17572 VGND.t3333 VGND.t1931 36.9323
R17573 VGND.t97 VGND.n206 36.9323
R17574 VGND.t6206 VGND.t6534 36.9323
R17575 VGND.t4374 VGND 36.9323
R17576 VGND.t6261 VGND.t2157 36.9323
R17577 VGND.t2155 VGND.t6289 36.9323
R17578 VGND.t171 VGND.t2786 36.9323
R17579 VGND.t948 VGND 36.9323
R17580 VGND.t4411 VGND.t6389 36.9323
R17581 VGND VGND.t6650 36.9323
R17582 VGND.t6708 VGND.t2296 36.9323
R17583 VGND.t4758 VGND.t716 36.9323
R17584 VGND.t3157 VGND.t6497 36.9323
R17585 VGND.t6663 VGND.t6511 36.9323
R17586 VGND.t4595 VGND.t153 36.9323
R17587 VGND.t4842 VGND.t6117 36.9323
R17588 VGND.t6610 VGND.t4847 36.9323
R17589 VGND.t6608 VGND.t4845 36.9323
R17590 VGND.t6144 VGND.t4273 36.9323
R17591 VGND.t3249 VGND.t5465 36.9323
R17592 VGND.t42 VGND.t4559 36.9323
R17593 VGND.t28 VGND.t3958 35.6658
R17594 VGND.t4522 VGND.t6616 35.6658
R17595 VGND.t4523 VGND.t6600 35.6658
R17596 VGND.t2876 VGND.t6606 35.6658
R17597 VGND.t2873 VGND.t6602 35.6658
R17598 VGND.t4525 VGND.t6604 35.6658
R17599 VGND.t4535 VGND.t6626 35.6658
R17600 VGND.t19 VGND.t2321 32.3158
R17601 VGND.t3642 VGND.t4718 27.6994
R17602 VGND.t3357 VGND.t2047 27.6994
R17603 VGND.t329 VGND.t4281 27.6994
R17604 VGND.t6786 VGND.t5684 27.6994
R17605 VGND.t1501 VGND.t4004 27.6994
R17606 VGND.t5902 VGND.t1243 27.6994
R17607 VGND.t2400 VGND.t2685 27.6994
R17608 VGND.t3594 VGND.t2689 27.6994
R17609 VGND.t5688 VGND.t1555 27.6994
R17610 VGND.t4959 VGND.t2918 27.6994
R17611 VGND.t2912 VGND.t4254 27.6994
R17612 VGND.t1312 VGND.t3017 27.6994
R17613 VGND.t5872 VGND.t1323 27.6994
R17614 VGND.t5991 VGND.t4382 27.6994
R17615 VGND.t1296 VGND.t1520 27.6994
R17616 VGND.t3277 VGND.t5014 27.6994
R17617 VGND.t2244 VGND.t663 27.2161
R17618 VGND VGND.t401 23.0829
R17619 VGND VGND.t4192 23.0829
R17620 VGND.t6792 VGND 23.0829
R17621 VGND VGND.t6306 23.0829
R17622 VGND.t938 VGND 23.0829
R17623 VGND.n2952 VGND.t5135 21.9565
R17624 VGND.t5096 VGND.n42 18.4664
R17625 VGND VGND.t6653 18.4664
R17626 VGND VGND.t1462 18.4664
R17627 VGND.t6008 VGND.t4903 18.4664
R17628 VGND VGND.t3614 18.4664
R17629 VGND.t5673 VGND 18.4664
R17630 VGND.t6746 VGND 18.4664
R17631 VGND VGND.t6719 18.4664
R17632 VGND.t6777 VGND.t6728 18.4664
R17633 VGND.t1454 VGND.t6204 18.4664
R17634 VGND VGND.t2361 18.4664
R17635 VGND.t2116 VGND 18.4664
R17636 VGND.t3941 VGND.t5054 18.4664
R17637 VGND VGND.t6350 18.4664
R17638 VGND VGND.t37 18.4664
R17639 VGND VGND.t6788 18.4664
R17640 VGND.n1499 VGND.t6295 18.4664
R17641 VGND.t4055 VGND.t3430 18.4664
R17642 VGND.t3426 VGND 18.4664
R17643 VGND.t6067 VGND.t611 18.4664
R17644 VGND VGND.t825 18.4664
R17645 VGND.t1055 VGND 18.4664
R17646 VGND VGND.t5229 18.4664
R17647 VGND VGND.t119 18.4664
R17648 VGND VGND.t3477 18.4664
R17649 VGND.t3726 VGND.t3211 18.4664
R17650 VGND VGND.t2279 18.4664
R17651 VGND VGND.t4006 18.4664
R17652 VGND VGND.t1239 18.4664
R17653 VGND.n605 VGND.t270 18.4664
R17654 VGND.t1679 VGND 18.4664
R17655 VGND.t5472 VGND.t6129 18.4664
R17656 VGND.t6379 VGND 18.4664
R17657 VGND VGND.t6642 18.4664
R17658 VGND VGND.t2512 18.4664
R17659 VGND VGND.t4323 18.4664
R17660 VGND.t246 VGND.t3124 18.4664
R17661 VGND VGND.t4692 18.4664
R17662 VGND VGND.t5734 18.4664
R17663 VGND.t428 VGND.t184 18.4664
R17664 VGND.t1827 VGND.t3232 18.4664
R17665 VGND.t6120 VGND.t3751 18.4664
R17666 VGND VGND.t637 18.4664
R17667 VGND VGND.t1074 18.4664
R17668 VGND VGND.t4493 18.4664
R17669 VGND.t5401 VGND 18.4664
R17670 VGND.t3245 VGND 18.4664
R17671 VGND.t6304 VGND 18.4664
R17672 VGND.t1673 VGND.t2094 18.4664
R17673 VGND.t2764 VGND.t206 18.4664
R17674 VGND VGND.t5029 18.4664
R17675 VGND.t1683 VGND 18.4664
R17676 VGND VGND.t723 18.4664
R17677 VGND VGND.t3189 18.4664
R17678 VGND.t1629 VGND 18.4664
R17679 VGND.t3812 VGND 18.4664
R17680 VGND.t305 VGND 18.4664
R17681 VGND VGND.t5980 18.4664
R17682 VGND.t6737 VGND.t2240 18.1443
R17683 VGND.n151 VGND.t4977 17.8331
R17684 VGND.t662 VGND.t6253 17.8331
R17685 VGND.t6588 VGND.t5796 13.8499
R17686 VGND.t6586 VGND.t5794 13.8499
R17687 VGND.n2165 VGND.n551 12.033
R17688 VGND.n2055 VGND.n562 12.033
R17689 VGND.n241 VGND.n227 12.033
R17690 VGND.n189 VGND.n181 12.033
R17691 VGND.n169 VGND.n160 12.033
R17692 VGND.n1410 VGND.n1402 12.033
R17693 VGND.n880 VGND.n870 12.033
R17694 VGND.n1567 VGND.n1357 12.033
R17695 VGND.n1375 VGND.n1373 12.033
R17696 VGND.n3422 VGND.n148 12.033
R17697 VGND.n3412 VGND.n155 12.033
R17698 VGND.n322 VGND.n275 12.033
R17699 VGND.n1397 VGND.n1361 12.033
R17700 VGND.n1540 VGND.n1489 12.033
R17701 VGND.n3390 VGND.n204 12.033
R17702 VGND.n262 VGND.n248 12.033
R17703 VGND.n3396 VGND.n201 12.033
R17704 VGND.n1549 VGND.n1486 12.033
R17705 VGND.n1476 VGND.n1474 12.033
R17706 VGND.n1657 VGND.n792 12.033
R17707 VGND.n1685 VGND.n775 12.033
R17708 VGND.n1739 VGND.n1732 12.033
R17709 VGND.n1751 VGND.n1728 12.033
R17710 VGND.n1764 VGND.n1723 12.033
R17711 VGND.n1781 VGND.n1717 12.033
R17712 VGND.n763 VGND.n730 12.033
R17713 VGND.n1808 VGND.n723 12.033
R17714 VGND.n1797 VGND.n727 12.033
R17715 VGND.n1982 VGND.n582 12.033
R17716 VGND.n1906 VGND.n664 12.033
R17717 VGND.n1985 VGND.n580 12.033
R17718 VGND.n954 VGND.n946 12.033
R17719 VGND.n2394 VGND.n477 12.033
R17720 VGND.n2199 VGND.n2197 12.033
R17721 VGND.n2385 VGND.n481 12.033
R17722 VGND.n2408 VGND.n471 12.033
R17723 VGND.n510 VGND.n509 12.033
R17724 VGND.n2363 VGND.n528 12.033
R17725 VGND.n2374 VGND.n524 12.033
R17726 VGND.n2163 VGND.t43 11.0292
R17727 VGND.n2057 VGND.t194 11.0292
R17728 VGND.n238 VGND.t138 11.0292
R17729 VGND.n187 VGND.t157 11.0292
R17730 VGND.n172 VGND.t6094 11.0292
R17731 VGND.n1407 VGND.t6743 11.0292
R17732 VGND.n883 VGND.t6634 11.0292
R17733 VGND.n1400 VGND.t6727 11.0292
R17734 VGND.n1374 VGND.t6738 11.0292
R17735 VGND.n3420 VGND.t91 11.0292
R17736 VGND.n3411 VGND.t6559 11.0292
R17737 VGND.n325 VGND.t6592 11.0292
R17738 VGND.n1394 VGND.t6776 11.0292
R17739 VGND.n1537 VGND.t6325 11.0292
R17740 VGND.n3387 VGND.t98 11.0292
R17741 VGND.n265 VGND.t6102 11.0292
R17742 VGND.n3393 VGND.t6068 11.0292
R17743 VGND.n1546 VGND.t228 11.0292
R17744 VGND.n1559 VGND.t142 11.0292
R17745 VGND.n1652 VGND.t6100 11.0292
R17746 VGND.n1682 VGND.t172 11.0292
R17747 VGND.n1736 VGND.t6681 11.0292
R17748 VGND.n1750 VGND.t6709 11.0292
R17749 VGND.n1760 VGND.t6474 11.0292
R17750 VGND.n1780 VGND.t31 11.0292
R17751 VGND.n767 VGND.t6130 11.0292
R17752 VGND.n1811 VGND.t6118 11.0292
R17753 VGND.n1800 VGND.t154 11.0292
R17754 VGND.n1984 VGND.t25 11.0292
R17755 VGND.n1903 VGND.t95 11.0292
R17756 VGND.n1988 VGND.t6313 11.0292
R17757 VGND.n956 VGND.t6145 11.0292
R17758 VGND.n2392 VGND.t6714 11.0292
R17759 VGND.n2169 VGND.t83 11.0292
R17760 VGND.n2388 VGND.t6192 11.0292
R17761 VGND.n950 VGND.t118 11.0292
R17762 VGND.n2380 VGND.t6731 11.0292
R17763 VGND.n2360 VGND.t6629 11.0292
R17764 VGND.n2377 VGND.t159 11.0292
R17765 VGND.n1578 VGND.t6722 10.9914
R17766 VGND.n1581 VGND.t645 10.9914
R17767 VGND.n1583 VGND.t17 10.9914
R17768 VGND.n1586 VGND.t886 10.9914
R17769 VGND.n1464 VGND.t6725 10.9914
R17770 VGND.n1468 VGND.t643 10.9914
R17771 VGND.n755 VGND.t1213 10.9914
R17772 VGND.n752 VGND.t4966 10.9914
R17773 VGND.n751 VGND.t1680 10.9914
R17774 VGND.n747 VGND.t231 10.9914
R17775 VGND.n1930 VGND.t6519 10.9914
R17776 VGND.n1928 VGND.t2513 10.9914
R17777 VGND.n819 VGND.t1078 10.9855
R17778 VGND.n815 VGND.t6564 10.9855
R17779 VGND.n316 VGND.t6587 10.9855
R17780 VGND.n1675 VGND.t4645 10.9855
R17781 VGND.n632 VGND.t4860 10.9855
R17782 VGND.n2039 VGND.t4313 10.9418
R17783 VGND.n320 VGND.t2599 10.9418
R17784 VGND.n1379 VGND.t6554 10.9418
R17785 VGND.n1669 VGND.t111 10.9418
R17786 VGND.n1953 VGND.t11 10.9418
R17787 VGND.n1973 VGND.t918 10.9418
R17788 VGND.n2401 VGND.t132 10.9418
R17789 VGND.n1420 VGND.t6411 10.5091
R17790 VGND.n1438 VGND.t6403 10.2792
R17791 VGND.n1432 VGND.t6405 10.2607
R17792 VGND.n925 VGND.t5882 10.0514
R17793 VGND.n921 VGND.t5884 10.0514
R17794 VGND.n851 VGND.t4517 10.0514
R17795 VGND.n855 VGND.t4518 10.0514
R17796 VGND.n3444 VGND.t4816 10.0514
R17797 VGND.n3448 VGND.t4813 10.0514
R17798 VGND.n928 VGND.t1063 10.0514
R17799 VGND.n933 VGND.t1061 10.0514
R17800 VGND.n1395 VGND.t4029 10.0514
R17801 VGND.n1391 VGND.t4033 10.0514
R17802 VGND.n1460 VGND.t2868 10.0514
R17803 VGND.n1457 VGND.t2866 10.0514
R17804 VGND.n2070 VGND.t3246 9.93604
R17805 VGND.n2083 VGND.t6581 9.93604
R17806 VGND.n2068 VGND.t6517 9.93604
R17807 VGND.n2031 VGND.t4161 9.93604
R17808 VGND.n827 VGND.t3210 9.93604
R17809 VGND.n859 VGND.t6458 9.93604
R17810 VGND.n824 VGND.t6698 9.93604
R17811 VGND.n1316 VGND.t324 9.93604
R17812 VGND.n1588 VGND.t6439 9.93604
R17813 VGND.n310 VGND.t6382 9.93604
R17814 VGND.n1566 VGND.t6499 9.93604
R17815 VGND.n1568 VGND.t6505 9.93604
R17816 VGND.n1592 VGND.t6720 9.93604
R17817 VGND.n1314 VGND.t3685 9.93604
R17818 VGND.n1311 VGND.t6570 9.93604
R17819 VGND.n1310 VGND.t2131 9.93604
R17820 VGND.n1470 VGND.t4064 9.93604
R17821 VGND.n1548 VGND.t5646 9.93604
R17822 VGND.n1514 VGND.t6789 9.93604
R17823 VGND.n255 VGND.t3061 9.93604
R17824 VGND.n1603 VGND.t15 9.93604
R17825 VGND.n838 VGND.t6351 9.93604
R17826 VGND.n1779 VGND.t5955 9.93604
R17827 VGND.n1149 VGND.t5903 9.93604
R17828 VGND.n640 VGND.t6417 9.93604
R17829 VGND.n626 VGND.t3146 9.93604
R17830 VGND.n2409 VGND.t4657 9.93604
R17831 VGND.n2166 VGND.t2228 9.93029
R17832 VGND.n128 VGND.t39 9.93029
R17833 VGND.n1343 VGND.t3342 9.93029
R17834 VGND.n301 VGND.t1183 9.93029
R17835 VGND.n1577 VGND.t2322 9.93029
R17836 VGND.n3406 VGND.t955 9.93029
R17837 VGND.n3391 VGND.t3486 9.93029
R17838 VGND.n1753 VGND.t6674 9.93029
R17839 VGND.n1774 VGND.t474 9.93029
R17840 VGND.n1707 VGND.t2057 9.93029
R17841 VGND.n1702 VGND.t5657 9.93029
R17842 VGND.n1929 VGND.t6640 9.93029
R17843 VGND.n1913 VGND.t5345 9.93029
R17844 VGND.n627 VGND.t182 9.93029
R17845 VGND.n2183 VGND.t5367 9.93029
R17846 VGND.n2201 VGND.t5265 9.93029
R17847 VGND.n2198 VGND.t2572 9.93029
R17848 VGND.n2396 VGND.t4318 9.93029
R17849 VGND.n2373 VGND.t4890 9.93029
R17850 VGND.n1655 VGND.t6275 9.8287
R17851 VGND.n1943 VGND.t275 9.8287
R17852 VGND.n1932 VGND.t6599 9.8287
R17853 VGND.n1670 VGND.t6268 9.82208
R17854 VGND.n1956 VGND.t297 9.82208
R17855 VGND.n644 VGND.t6619 9.82208
R17856 VGND.n909 VGND.t1304 9.80518
R17857 VGND.n802 VGND.t335 9.80518
R17858 VGND.n800 VGND.t2788 9.80518
R17859 VGND.n847 VGND.t3985 9.80518
R17860 VGND.n1504 VGND.t3433 9.74705
R17861 VGND.n2049 VGND.t4995 9.6277
R17862 VGND.n162 VGND.t6794 9.6277
R17863 VGND.n1249 VGND.t3942 9.6277
R17864 VGND.n3397 VGND.t6143 9.6277
R17865 VGND.n3384 VGND.t4375 9.6277
R17866 VGND.n1506 VGND.t4056 9.6277
R17867 VGND.n1523 VGND.t6255 9.6277
R17868 VGND.n1786 VGND.t6467 9.6277
R17869 VGND.n1771 VGND.t6651 9.6277
R17870 VGND.n1698 VGND.t949 9.6277
R17871 VGND.n643 VGND.t3125 9.6277
R17872 VGND.n636 VGND.t4858 9.6277
R17873 VGND.n2387 VGND.t3251 9.6277
R17874 VGND.n2187 VGND.t6645 9.6277
R17875 VGND.n485 VGND.t2627 9.6277
R17876 VGND.n1965 VGND.t5388 9.56913
R17877 VGND.n2045 VGND.t129 9.38548
R17878 VGND.n2047 VGND.t6414 9.38548
R17879 VGND.n2084 VGND.t2452 9.38548
R17880 VGND.n2082 VGND.t6305 9.38548
R17881 VGND.n831 VGND.t6699 9.38548
R17882 VGND.n829 VGND.t6454 9.38548
R17883 VGND.n3443 VGND.t2239 9.38548
R17884 VGND.n3441 VGND.t5705 9.38548
R17885 VGND.n3440 VGND.t5708 9.38548
R17886 VGND.n3439 VGND.t6340 9.38548
R17887 VGND.n3437 VGND.t6470 9.38548
R17888 VGND.n3435 VGND.t3409 9.38548
R17889 VGND.n167 VGND.t103 9.38548
R17890 VGND.n168 VGND.t6652 9.38548
R17891 VGND.n174 VGND.t6339 9.38548
R17892 VGND.n175 VGND.t5613 9.38548
R17893 VGND.n226 VGND.t6391 9.38548
R17894 VGND.n242 VGND.t6585 9.38548
R17895 VGND.n139 VGND.t3326 9.38548
R17896 VGND.n3434 VGND.t109 9.38548
R17897 VGND.n863 VGND.t6462 9.38548
R17898 VGND.n862 VGND.t6445 9.38548
R17899 VGND.n886 VGND.t2630 9.38548
R17900 VGND.n1593 VGND.t196 9.38548
R17901 VGND.n291 VGND.t1106 9.38548
R17902 VGND.n292 VGND.t6399 9.38548
R17903 VGND.n294 VGND.t4730 9.38548
R17904 VGND.n295 VGND.t2429 9.38548
R17905 VGND.n324 VGND.t2458 9.38548
R17906 VGND.n326 VGND.t6393 9.38548
R17907 VGND.n302 VGND.t3938 9.38548
R17908 VGND.n300 VGND.t1179 9.38548
R17909 VGND.n1601 VGND.t889 9.38548
R17910 VGND.n1529 VGND.t105 9.38548
R17911 VGND.n1527 VGND.t6252 9.38548
R17912 VGND.n1507 VGND.t953 9.38548
R17913 VGND.n1509 VGND.t6234 9.38548
R17914 VGND.n1517 VGND.t107 9.38548
R17915 VGND.n1519 VGND.t6791 9.38548
R17916 VGND.n1541 VGND.t6550 9.38548
R17917 VGND.n1542 VGND.t213 9.38548
R17918 VGND.n1465 VGND.t3691 9.38548
R17919 VGND.n1463 VGND.t116 9.38548
R17920 VGND.n1599 VGND.t5623 9.38548
R17921 VGND.n1708 VGND.t4963 9.38548
R17922 VGND.n1710 VGND.t6546 9.38548
R17923 VGND.n1758 VGND.t2816 9.38548
R17924 VGND.n1757 VGND.t6386 9.38548
R17925 VGND.n1697 VGND.t4533 9.38548
R17926 VGND.n1695 VGND.t6156 9.38548
R17927 VGND.n1681 VGND.t3154 9.38548
R17928 VGND.n1679 VGND.t120 9.38548
R17929 VGND.n799 VGND.t6688 9.38548
R17930 VGND.n1209 VGND.t4562 9.38548
R17931 VGND.n1925 VGND.t6322 9.38548
R17932 VGND.n1923 VGND.t3198 9.38548
R17933 VGND.n1920 VGND.t6544 9.38548
R17934 VGND.n1918 VGND.t6303 9.38548
R17935 VGND.n1908 VGND.t6105 9.38548
R17936 VGND.n1907 VGND.t6317 9.38548
R17937 VGND.n1917 VGND.t4324 9.38548
R17938 VGND.n1919 VGND.t3204 9.38548
R17939 VGND.n2193 VGND.t6572 9.38548
R17940 VGND.n2205 VGND.t2568 9.38548
R17941 VGND.n2364 VGND.t215 9.38548
R17942 VGND.n2365 VGND.t4404 9.38548
R17943 VGND.n744 VGND.t2330 9.31505
R17944 VGND.n635 VGND.t6423 9.31505
R17945 VGND.n1431 VGND.t3516 9.25462
R17946 VGND.n3447 VGND.t3513 9.25462
R17947 VGND.n134 VGND.t1139 9.25462
R17948 VGND.n125 VGND.t1142 9.25462
R17949 VGND.n129 VGND.t147 9.25462
R17950 VGND.n138 VGND.t150 9.25462
R17951 VGND.n3436 VGND.t6063 9.25462
R17952 VGND.n3442 VGND.t6064 9.25462
R17953 VGND.n1390 VGND.t5704 9.25462
R17954 VGND.n1383 VGND.t5699 9.25462
R17955 VGND.n1525 VGND.t1926 9.25462
R17956 VGND.n1516 VGND.t1930 9.25462
R17957 VGND.n857 VGND.t7 9.17206
R17958 VGND.n1461 VGND.t6464 9.17206
R17959 VGND.n808 VGND.t6736 9.15882
R17960 VGND.n3450 VGND.t6242 9.15882
R17961 VGND.n926 VGND.t6072 9.15882
R17962 VGND.n1396 VGND.t1610 9.15882
R17963 VGND.n801 VGND.t3683 8.76488
R17964 VGND.n1493 VGND.t472 8.76488
R17965 VGND.n1719 VGND.t6669 8.76488
R17966 VGND.n661 VGND.t6109 8.76488
R17967 VGND.n2173 VGND.t6126 8.76488
R17968 VGND.n525 VGND.t5369 8.76488
R17969 VGND.n2053 VGND.t4311 8.76406
R17970 VGND.n1579 VGND.t1784 8.76406
R17971 VGND.n3414 VGND.t2946 8.76406
R17972 VGND.n1300 VGND.t4704 8.76406
R17973 VGND.n1208 VGND.t4199 8.76406
R17974 VGND.n750 VGND.t4681 8.76406
R17975 VGND.n1819 VGND.t6672 8.76406
R17976 VGND.n832 VGND.t5102 8.71342
R17977 VGND.n1298 VGND.t6561 8.71342
R17978 VGND.n3358 VGND.t5542 8.65297
R17979 VGND.n559 VGND.t3680 8.63064
R17980 VGND.n740 VGND.t3215 8.63064
R17981 VGND.n611 VGND.t3470 8.52948
R17982 VGND.n631 VGND.t1405 8.52948
R17983 VGND.n1959 VGND.t870 8.51593
R17984 VGND.n1020 VGND.t5222 8.51132
R17985 VGND.n2006 VGND.t3944 8.51132
R17986 VGND.n2023 VGND.t5987 8.51132
R17987 VGND.n2025 VGND.t5002 8.51132
R17988 VGND.n2027 VGND.t1852 8.51132
R17989 VGND.n2029 VGND.t1759 8.51132
R17990 VGND.n2032 VGND.t1670 8.51132
R17991 VGND.n2041 VGND.t2902 8.51132
R17992 VGND.n2043 VGND.t4506 8.51132
R17993 VGND.n2072 VGND.t4109 8.51132
R17994 VGND.n2074 VGND.t4701 8.51132
R17995 VGND.n2085 VGND.t5583 8.51132
R17996 VGND.n2090 VGND.t5418 8.51132
R17997 VGND.n2088 VGND.t2095 8.51132
R17998 VGND.n2162 VGND.t4560 8.51132
R17999 VGND.n2159 VGND.t4396 8.51132
R18000 VGND.n2157 VGND.t5068 8.51132
R18001 VGND.n2155 VGND.t5554 8.51132
R18002 VGND.n2153 VGND.t3588 8.51132
R18003 VGND.n2151 VGND.t6035 8.51132
R18004 VGND.n2149 VGND.t3926 8.51132
R18005 VGND.n2147 VGND.t971 8.51132
R18006 VGND.n2145 VGND.t3697 8.51132
R18007 VGND.n2143 VGND.t5950 8.51132
R18008 VGND.n2140 VGND.t2742 8.51132
R18009 VGND.n2138 VGND.t1299 8.51132
R18010 VGND.n2136 VGND.t3878 8.51132
R18011 VGND.n2134 VGND.t5927 8.51132
R18012 VGND.n2131 VGND.t2062 8.51132
R18013 VGND.n2129 VGND.t2893 8.51132
R18014 VGND.n2127 VGND.t4807 8.51132
R18015 VGND.n2125 VGND.t2967 8.51132
R18016 VGND.n2122 VGND.t2113 8.51132
R18017 VGND.n2120 VGND.t1790 8.51132
R18018 VGND.n2118 VGND.t4167 8.51132
R18019 VGND.n2116 VGND.t2135 8.51132
R18020 VGND.n2114 VGND.t4268 8.51132
R18021 VGND.n2112 VGND.t4025 8.51132
R18022 VGND.n2110 VGND.t4569 8.51132
R18023 VGND.n2108 VGND.t1707 8.51132
R18024 VGND.n2106 VGND.t3051 8.51132
R18025 VGND.n2104 VGND.t2539 8.51132
R18026 VGND.n2102 VGND.t3407 8.51132
R18027 VGND.n2100 VGND.t2423 8.51132
R18028 VGND.n2098 VGND.t3775 8.51132
R18029 VGND.n3339 VGND.t5526 8.51132
R18030 VGND.n3341 VGND.t973 8.51132
R18031 VGND.n3343 VGND.t4452 8.51132
R18032 VGND.n3345 VGND.t3346 8.51132
R18033 VGND.n3349 VGND.t3374 8.51132
R18034 VGND.n3349 VGND.t370 8.51132
R18035 VGND.n3350 VGND.t3541 8.51132
R18036 VGND.n3350 VGND.t5840 8.51132
R18037 VGND.n3351 VGND.t2026 8.51132
R18038 VGND.n3351 VGND.t2882 8.51132
R18039 VGND.n3352 VGND.t1006 8.51132
R18040 VGND.n3352 VGND.t1079 8.51132
R18041 VGND.n3353 VGND.t2201 8.51132
R18042 VGND.n3353 VGND.t2846 8.51132
R18043 VGND.n3354 VGND.t4116 8.51132
R18044 VGND.n3354 VGND.t3166 8.51132
R18045 VGND.n3355 VGND.t1042 8.51132
R18046 VGND.n3355 VGND.t5729 8.51132
R18047 VGND.n3356 VGND.t3781 8.51132
R18048 VGND.n3356 VGND.t1579 8.51132
R18049 VGND.n3346 VGND.t1391 8.51132
R18050 VGND.n3344 VGND.t975 8.51132
R18051 VGND.n3342 VGND.t2346 8.51132
R18052 VGND.n3340 VGND.t1727 8.51132
R18053 VGND.n2097 VGND.t2427 8.51132
R18054 VGND.n2099 VGND.t2750 8.51132
R18055 VGND.n2101 VGND.t1717 8.51132
R18056 VGND.n2103 VGND.t4441 8.51132
R18057 VGND.n2107 VGND.t996 8.51132
R18058 VGND.n2109 VGND.t4902 8.51132
R18059 VGND.n2111 VGND.t5921 8.51132
R18060 VGND.n2113 VGND.t5200 8.51132
R18061 VGND.n2115 VGND.t3695 8.51132
R18062 VGND.n2117 VGND.t1792 8.51132
R18063 VGND.n2119 VGND.t3605 8.51132
R18064 VGND.n2121 VGND.t1435 8.51132
R18065 VGND.n2123 VGND.t3601 8.51132
R18066 VGND.n2126 VGND.t2872 8.51132
R18067 VGND.n2128 VGND.t5976 8.51132
R18068 VGND.n2130 VGND.t3539 8.51132
R18069 VGND.n2133 VGND.t3091 8.51132
R18070 VGND.n2135 VGND.t4368 8.51132
R18071 VGND.n2137 VGND.t1744 8.51132
R18072 VGND.n2139 VGND.t567 8.51132
R18073 VGND.n2142 VGND.t4736 8.51132
R18074 VGND.n2144 VGND.t4353 8.51132
R18075 VGND.n2146 VGND.t2184 8.51132
R18076 VGND.n2148 VGND.t2224 8.51132
R18077 VGND.n2150 VGND.t5482 8.51132
R18078 VGND.n2152 VGND.t2848 8.51132
R18079 VGND.n2154 VGND.t5398 8.51132
R18080 VGND.n2156 VGND.t4464 8.51132
R18081 VGND.n2081 VGND.t5905 8.51132
R18082 VGND.n2080 VGND.t3040 8.51132
R18083 VGND.n2076 VGND.t1411 8.51132
R18084 VGND.n2075 VGND.t486 8.51132
R18085 VGND.n2073 VGND.t1742 8.51132
R18086 VGND.n2042 VGND.t2150 8.51132
R18087 VGND.n2030 VGND.t2328 8.51132
R18088 VGND.n2028 VGND.t3257 8.51132
R18089 VGND.n2026 VGND.t5373 8.51132
R18090 VGND.n2024 VGND.t5390 8.51132
R18091 VGND.n2009 VGND.t2387 8.51132
R18092 VGND.n2007 VGND.t1870 8.51132
R18093 VGND.n1035 VGND.t5176 8.51132
R18094 VGND.n1037 VGND.t544 8.51132
R18095 VGND.n1040 VGND.t5142 8.51132
R18096 VGND.n1047 VGND.t2214 8.51132
R18097 VGND.n1063 VGND.t4434 8.51132
R18098 VGND.n1065 VGND.t4661 8.51132
R18099 VGND.n1018 VGND.t3653 8.51132
R18100 VGND.n1016 VGND.t994 8.51132
R18101 VGND.n3672 VGND.t3655 8.51132
R18102 VGND.n3670 VGND.t5333 8.51132
R18103 VGND.n3681 VGND.t3109 8.51132
R18104 VGND.n3681 VGND.t1575 8.51132
R18105 VGND.n3680 VGND.t3457 8.51132
R18106 VGND.n3680 VGND.t3010 8.51132
R18107 VGND.n3679 VGND.t4402 8.51132
R18108 VGND.n3679 VGND.t2752 8.51132
R18109 VGND.n3678 VGND.t3832 8.51132
R18110 VGND.n3678 VGND.t2684 8.51132
R18111 VGND.n3677 VGND.t4205 8.51132
R18112 VGND.n3677 VGND.t5767 8.51132
R18113 VGND.n3676 VGND.t1261 8.51132
R18114 VGND.n3676 VGND.t3123 8.51132
R18115 VGND.n3675 VGND.t5932 8.51132
R18116 VGND.n3675 VGND.t5799 8.51132
R18117 VGND.n3674 VGND.t5276 8.51132
R18118 VGND.n3674 VGND.t4713 8.51132
R18119 VGND.n3682 VGND.t3415 8.51132
R18120 VGND.n3671 VGND.t4753 8.51132
R18121 VGND.n3483 VGND.t6807 8.51132
R18122 VGND.n3485 VGND.t421 8.51132
R18123 VGND.n3493 VGND.t5655 8.51132
R18124 VGND.n3493 VGND.t4833 8.51132
R18125 VGND.n3492 VGND.t5040 8.51132
R18126 VGND.n3492 VGND.t4408 8.51132
R18127 VGND.n3491 VGND.t409 8.51132
R18128 VGND.n3491 VGND.t6087 8.51132
R18129 VGND.n3490 VGND.t3408 8.51132
R18130 VGND.n3490 VGND.t1399 8.51132
R18131 VGND.n3489 VGND.t4760 8.51132
R18132 VGND.n3489 VGND.t620 8.51132
R18133 VGND.n3488 VGND.t2534 8.51132
R18134 VGND.n3488 VGND.t2282 8.51132
R18135 VGND.n3487 VGND.t3344 8.51132
R18136 VGND.n3487 VGND.t5969 8.51132
R18137 VGND.n3486 VGND.t1802 8.51132
R18138 VGND.n3486 VGND.t767 8.51132
R18139 VGND.n3494 VGND.t2009 8.51132
R18140 VGND.n3484 VGND.t4472 8.51132
R18141 VGND.n3635 VGND.t1457 8.51132
R18142 VGND.n3637 VGND.t1748 8.51132
R18143 VGND.n3646 VGND.t3055 8.51132
R18144 VGND.n3646 VGND.t5879 8.51132
R18145 VGND.n3645 VGND.t2884 8.51132
R18146 VGND.n3645 VGND.t4629 8.51132
R18147 VGND.n3644 VGND.t5443 8.51132
R18148 VGND.n3644 VGND.t3669 8.51132
R18149 VGND.n3643 VGND.t4097 8.51132
R18150 VGND.n3643 VGND.t2209 8.51132
R18151 VGND.n3642 VGND.t3849 8.51132
R18152 VGND.n3642 VGND.t641 8.51132
R18153 VGND.n3641 VGND.t1315 8.51132
R18154 VGND.n3641 VGND.t4001 8.51132
R18155 VGND.n3640 VGND.t2188 8.51132
R18156 VGND.n3640 VGND.t5814 8.51132
R18157 VGND.n3639 VGND.t3840 8.51132
R18158 VGND.n3639 VGND.t4976 8.51132
R18159 VGND.n3647 VGND.t2647 8.51132
R18160 VGND.n3636 VGND.t3963 8.51132
R18161 VGND.n3650 VGND.t4545 8.51132
R18162 VGND.n3652 VGND.t3137 8.51132
R18163 VGND.n3661 VGND.t1911 8.51132
R18164 VGND.n3661 VGND.t1366 8.51132
R18165 VGND.n3660 VGND.t2936 8.51132
R18166 VGND.n3660 VGND.t6764 8.51132
R18167 VGND.n3659 VGND.t2193 8.51132
R18168 VGND.n3659 VGND.t2564 8.51132
R18169 VGND.n3658 VGND.t3393 8.51132
R18170 VGND.n3658 VGND.t2944 8.51132
R18171 VGND.n3657 VGND.t4954 8.51132
R18172 VGND.n3657 VGND.t2978 8.51132
R18173 VGND.n3656 VGND.t4473 8.51132
R18174 VGND.n3656 VGND.t4186 8.51132
R18175 VGND.n3655 VGND.t4609 8.51132
R18176 VGND.n3655 VGND.t417 8.51132
R18177 VGND.n3654 VGND.t3831 8.51132
R18178 VGND.n3654 VGND.t2682 8.51132
R18179 VGND.n3662 VGND.t2536 8.51132
R18180 VGND.n3651 VGND.t4344 8.51132
R18181 VGND.n3466 VGND.t1267 8.51132
R18182 VGND.n3468 VGND.t1903 8.51132
R18183 VGND.n3476 VGND.t556 8.51132
R18184 VGND.n3476 VGND.t1364 8.51132
R18185 VGND.n3475 VGND.t1087 8.51132
R18186 VGND.n3475 VGND.t64 8.51132
R18187 VGND.n3474 VGND.t5715 8.51132
R18188 VGND.n3474 VGND.t2589 8.51132
R18189 VGND.n3473 VGND.t1290 8.51132
R18190 VGND.n3473 VGND.t2881 8.51132
R18191 VGND.n3472 VGND.t5476 8.51132
R18192 VGND.n3472 VGND.t5331 8.51132
R18193 VGND.n3471 VGND.t1317 8.51132
R18194 VGND.n3471 VGND.t3000 8.51132
R18195 VGND.n3470 VGND.t4260 8.51132
R18196 VGND.n3470 VGND.t651 8.51132
R18197 VGND.n3469 VGND.t5171 8.51132
R18198 VGND.n3469 VGND.t2176 8.51132
R18199 VGND.n3477 VGND.t2268 8.51132
R18200 VGND.n3467 VGND.t4228 8.51132
R18201 VGND.n3574 VGND.t518 8.51132
R18202 VGND.n3572 VGND.t5196 8.51132
R18203 VGND.n3583 VGND.t3445 8.51132
R18204 VGND.n3583 VGND.t5972 8.51132
R18205 VGND.n3582 VGND.t3827 8.51132
R18206 VGND.n3582 VGND.t3543 8.51132
R18207 VGND.n3581 VGND.t3618 8.51132
R18208 VGND.n3581 VGND.t855 8.51132
R18209 VGND.n3580 VGND.t3762 8.51132
R18210 VGND.n3580 VGND.t2462 8.51132
R18211 VGND.n3579 VGND.t743 8.51132
R18212 VGND.n3579 VGND.t1040 8.51132
R18213 VGND.n3578 VGND.t4154 8.51132
R18214 VGND.n3578 VGND.t5197 8.51132
R18215 VGND.n3577 VGND.t2107 8.51132
R18216 VGND.n3577 VGND.t5527 8.51132
R18217 VGND.n3576 VGND.t4618 8.51132
R18218 VGND.n3576 VGND.t3194 8.51132
R18219 VGND.n3584 VGND.t2607 8.51132
R18220 VGND.n3573 VGND.t3320 8.51132
R18221 VGND.n3606 VGND.t4262 8.51132
R18222 VGND.n3604 VGND.t3504 8.51132
R18223 VGND.n3615 VGND.t2195 8.51132
R18224 VGND.n3615 VGND.t5158 8.51132
R18225 VGND.n3614 VGND.t5499 8.51132
R18226 VGND.n3614 VGND.t5780 8.51132
R18227 VGND.n3613 VGND.t4180 8.51132
R18228 VGND.n3613 VGND.t1723 8.51132
R18229 VGND.n3612 VGND.t4251 8.51132
R18230 VGND.n3612 VGND.t355 8.51132
R18231 VGND.n3611 VGND.t1803 8.51132
R18232 VGND.n3611 VGND.t490 8.51132
R18233 VGND.n3610 VGND.t5837 8.51132
R18234 VGND.n3610 VGND.t2850 8.51132
R18235 VGND.n3609 VGND.t5536 8.51132
R18236 VGND.n3609 VGND.t3508 8.51132
R18237 VGND.n3608 VGND.t1021 8.51132
R18238 VGND.n3608 VGND.t62 8.51132
R18239 VGND.n3616 VGND.t4827 8.51132
R18240 VGND.n3605 VGND.t1668 8.51132
R18241 VGND.n3622 VGND.t6756 8.51132
R18242 VGND.n3620 VGND.t1084 8.51132
R18243 VGND.n3631 VGND.t1031 8.51132
R18244 VGND.n3631 VGND.t2231 8.51132
R18245 VGND.n3630 VGND.t5584 8.51132
R18246 VGND.n3630 VGND.t4128 8.51132
R18247 VGND.n3629 VGND.t5214 8.51132
R18248 VGND.n3629 VGND.t6762 8.51132
R18249 VGND.n3628 VGND.t3077 8.51132
R18250 VGND.n3628 VGND.t6163 8.51132
R18251 VGND.n3627 VGND.t3848 8.51132
R18252 VGND.n3627 VGND.t558 8.51132
R18253 VGND.n3626 VGND.t4157 8.51132
R18254 VGND.n3626 VGND.t1089 8.51132
R18255 VGND.n3625 VGND.t2712 8.51132
R18256 VGND.n3625 VGND.t4935 8.51132
R18257 VGND.n3624 VGND.t623 8.51132
R18258 VGND.n3624 VGND.t5066 8.51132
R18259 VGND.n3632 VGND.t2226 8.51132
R18260 VGND.n3621 VGND.t2529 8.51132
R18261 VGND.n3590 VGND.t2089 8.51132
R18262 VGND.n3588 VGND.t2716 8.51132
R18263 VGND.n3599 VGND.t2014 8.51132
R18264 VGND.n3599 VGND.t906 8.51132
R18265 VGND.n3598 VGND.t1878 8.51132
R18266 VGND.n3598 VGND.t6769 8.51132
R18267 VGND.n3597 VGND.t4442 8.51132
R18268 VGND.n3597 VGND.t2081 8.51132
R18269 VGND.n3596 VGND.t1498 8.51132
R18270 VGND.n3596 VGND.t3008 8.51132
R18271 VGND.n3595 VGND.t4082 8.51132
R18272 VGND.n3595 VGND.t3512 8.51132
R18273 VGND.n3594 VGND.t1938 8.51132
R18274 VGND.n3594 VGND.t2822 8.51132
R18275 VGND.n3593 VGND.t1170 8.51132
R18276 VGND.n3593 VGND.t2291 8.51132
R18277 VGND.n3592 VGND.t4043 8.51132
R18278 VGND.n3592 VGND.t3971 8.51132
R18279 VGND.n3600 VGND.t1660 8.51132
R18280 VGND.n3589 VGND.t2488 8.51132
R18281 VGND.n3558 VGND.t5283 8.51132
R18282 VGND.n3556 VGND.t5120 8.51132
R18283 VGND.n3567 VGND.t2127 8.51132
R18284 VGND.n3567 VGND.t5052 8.51132
R18285 VGND.n3566 VGND.t3778 8.51132
R18286 VGND.n3566 VGND.t783 8.51132
R18287 VGND.n3565 VGND.t4900 8.51132
R18288 VGND.n3565 VGND.t5577 8.51132
R18289 VGND.n3564 VGND.t2925 8.51132
R18290 VGND.n3564 VGND.t4504 8.51132
R18291 VGND.n3563 VGND.t3722 8.51132
R18292 VGND.n3563 VGND.t1840 8.51132
R18293 VGND.n3562 VGND.t2563 8.51132
R18294 VGND.n3562 VGND.t1215 8.51132
R18295 VGND.n3561 VGND.t1765 8.51132
R18296 VGND.n3561 VGND.t3723 8.51132
R18297 VGND.n3560 VGND.t4438 8.51132
R18298 VGND.n3560 VGND.t2007 8.51132
R18299 VGND.n3568 VGND.t6783 8.51132
R18300 VGND.n3557 VGND.t1695 8.51132
R18301 VGND.n3540 VGND.t1543 8.51132
R18302 VGND.n3542 VGND.t5811 8.51132
R18303 VGND.n3551 VGND.t4009 8.51132
R18304 VGND.n3551 VGND.t5953 8.51132
R18305 VGND.n3550 VGND.t3043 8.51132
R18306 VGND.n3550 VGND.t2730 8.51132
R18307 VGND.n3549 VGND.t3221 8.51132
R18308 VGND.n3549 VGND.t2708 8.51132
R18309 VGND.n3548 VGND.t3808 8.51132
R18310 VGND.n3548 VGND.t2897 8.51132
R18311 VGND.n3547 VGND.t5614 8.51132
R18312 VGND.n3547 VGND.t1050 8.51132
R18313 VGND.n3546 VGND.t1709 8.51132
R18314 VGND.n3546 VGND.t5233 8.51132
R18315 VGND.n3545 VGND.t1909 8.51132
R18316 VGND.n3545 VGND.t5111 8.51132
R18317 VGND.n3544 VGND.t4373 8.51132
R18318 VGND.n3544 VGND.t5237 8.51132
R18319 VGND.n3552 VGND.t4364 8.51132
R18320 VGND.n3541 VGND.t4042 8.51132
R18321 VGND.n3703 VGND.t3687 8.51132
R18322 VGND.n3701 VGND.t2060 8.51132
R18323 VGND.n3712 VGND.t2541 8.51132
R18324 VGND.n3712 VGND.t5860 8.51132
R18325 VGND.n3711 VGND.t4939 8.51132
R18326 VGND.n3711 VGND.t5281 8.51132
R18327 VGND.n3710 VGND.t3295 8.51132
R18328 VGND.n3710 VGND.t4014 8.51132
R18329 VGND.n3709 VGND.t4501 8.51132
R18330 VGND.n3709 VGND.t4201 8.51132
R18331 VGND.n3708 VGND.t1473 8.51132
R18332 VGND.n3708 VGND.t372 8.51132
R18333 VGND.n3707 VGND.t5675 8.51132
R18334 VGND.n3707 VGND.t3500 8.51132
R18335 VGND.n3706 VGND.t3021 8.51132
R18336 VGND.n3706 VGND.t502 8.51132
R18337 VGND.n3705 VGND.t321 8.51132
R18338 VGND.n3705 VGND.t1675 8.51132
R18339 VGND.n3713 VGND.t4214 8.51132
R18340 VGND.n3702 VGND.t5118 8.51132
R18341 VGND.n22 VGND.t4062 8.51132
R18342 VGND.n24 VGND.t3580 8.51132
R18343 VGND.n32 VGND.t1376 8.51132
R18344 VGND.n32 VGND.t3299 8.51132
R18345 VGND.n31 VGND.t5946 8.51132
R18346 VGND.n31 VGND.t1131 8.51132
R18347 VGND.n30 VGND.t5676 8.51132
R18348 VGND.n30 VGND.t2714 8.51132
R18349 VGND.n29 VGND.t2889 8.51132
R18350 VGND.n29 VGND.t763 8.51132
R18351 VGND.n28 VGND.t449 8.51132
R18352 VGND.n28 VGND.t4070 8.51132
R18353 VGND.n27 VGND.t5765 8.51132
R18354 VGND.n27 VGND.t2143 8.51132
R18355 VGND.n26 VGND.t2773 8.51132
R18356 VGND.n26 VGND.t3603 8.51132
R18357 VGND.n25 VGND.t1407 8.51132
R18358 VGND.n25 VGND.t2482 8.51132
R18359 VGND.n33 VGND.t4179 8.51132
R18360 VGND.n23 VGND.t5354 8.51132
R18361 VGND.n3495 VGND.t3451 8.51132
R18362 VGND.n3497 VGND.t5140 8.51132
R18363 VGND.n3506 VGND.t5152 8.51132
R18364 VGND.n3506 VGND.t731 8.51132
R18365 VGND.n3505 VGND.t5750 8.51132
R18366 VGND.n3505 VGND.t4081 8.51132
R18367 VGND.n3504 VGND.t2621 8.51132
R18368 VGND.n3504 VGND.t363 8.51132
R18369 VGND.n3503 VGND.t2087 8.51132
R18370 VGND.n3503 VGND.t5172 8.51132
R18371 VGND.n3502 VGND.t3756 8.51132
R18372 VGND.n3502 VGND.t4386 8.51132
R18373 VGND.n3501 VGND.t734 8.51132
R18374 VGND.n3501 VGND.t1 8.51132
R18375 VGND.n3500 VGND.t3063 8.51132
R18376 VGND.n3500 VGND.t5856 8.51132
R18377 VGND.n3499 VGND.t353 8.51132
R18378 VGND.n3499 VGND.t4439 8.51132
R18379 VGND.n3507 VGND.t3582 8.51132
R18380 VGND.n3496 VGND.t5339 8.51132
R18381 VGND.n3510 VGND.t1874 8.51132
R18382 VGND.n3512 VGND.t3965 8.51132
R18383 VGND.n3521 VGND.t3106 8.51132
R18384 VGND.n3521 VGND.t3032 8.51132
R18385 VGND.n3520 VGND.t5640 8.51132
R18386 VGND.n3520 VGND.t6073 8.51132
R18387 VGND.n3519 VGND.t3254 8.51132
R18388 VGND.n3519 VGND.t2270 8.51132
R18389 VGND.n3518 VGND.t6084 8.51132
R18390 VGND.n3518 VGND.t4075 8.51132
R18391 VGND.n3517 VGND.t608 8.51132
R18392 VGND.n3517 VGND.t3933 8.51132
R18393 VGND.n3516 VGND.t653 8.51132
R18394 VGND.n3516 VGND.t1889 8.51132
R18395 VGND.n3515 VGND.t6183 8.51132
R18396 VGND.n3515 VGND.t2440 8.51132
R18397 VGND.n3514 VGND.t476 8.51132
R18398 VGND.n3514 VGND.t4733 8.51132
R18399 VGND.n3522 VGND.t74 8.51132
R18400 VGND.n3511 VGND.t5821 8.51132
R18401 VGND.n3525 VGND.t1231 8.51132
R18402 VGND.n3527 VGND.t4637 8.51132
R18403 VGND.n3536 VGND.t4921 8.51132
R18404 VGND.n3536 VGND.t1642 8.51132
R18405 VGND.n3535 VGND.t3874 8.51132
R18406 VGND.n3535 VGND.t998 8.51132
R18407 VGND.n3534 VGND.t647 8.51132
R18408 VGND.n3534 VGND.t1894 8.51132
R18409 VGND.n3533 VGND.t2587 8.51132
R18410 VGND.n3533 VGND.t6080 8.51132
R18411 VGND.n3532 VGND.t3846 8.51132
R18412 VGND.n3532 VGND.t4486 8.51132
R18413 VGND.n3531 VGND.t3340 8.51132
R18414 VGND.n3531 VGND.t4638 8.51132
R18415 VGND.n3530 VGND.t4187 8.51132
R18416 VGND.n3530 VGND.t1800 8.51132
R18417 VGND.n3529 VGND.t5576 8.51132
R18418 VGND.n3529 VGND.t3891 8.51132
R18419 VGND.n3537 VGND.t3780 8.51132
R18420 VGND.n3526 VGND.t2285 8.51132
R18421 VGND.n927 VGND.t5115 8.51132
R18422 VGND.n828 VGND.t4679 8.51132
R18423 VGND.n827 VGND.t5599 8.51132
R18424 VGND.n867 VGND.t2628 8.51132
R18425 VGND.n879 VGND.t1096 8.51132
R18426 VGND.n878 VGND.t2911 8.51132
R18427 VGND.n877 VGND.t2829 8.51132
R18428 VGND.n874 VGND.t2455 8.51132
R18429 VGND.n872 VGND.t5250 8.51132
R18430 VGND.n1404 VGND.t5124 8.51132
R18431 VGND.n1406 VGND.t1857 8.51132
R18432 VGND.n1408 VGND.t5352 8.51132
R18433 VGND.n1411 VGND.t6805 8.51132
R18434 VGND.n1412 VGND.t621 8.51132
R18435 VGND.n1414 VGND.t4123 8.51132
R18436 VGND.n1416 VGND.t3132 8.51132
R18437 VGND.n1417 VGND.t1385 8.51132
R18438 VGND.n1419 VGND.t6004 8.51132
R18439 VGND.n1441 VGND.t709 8.51132
R18440 VGND.n1439 VGND.t5304 8.51132
R18441 VGND.n140 VGND.t2625 8.51132
R18442 VGND.n137 VGND.t1358 8.51132
R18443 VGND.n164 VGND.t2180 8.51132
R18444 VGND.n170 VGND.t1160 8.51132
R18445 VGND.n193 VGND.t761 8.51132
R18446 VGND.n191 VGND.t2408 8.51132
R18447 VGND.n190 VGND.t3255 8.51132
R18448 VGND.n186 VGND.t5937 8.51132
R18449 VGND.n184 VGND.t1582 8.51132
R18450 VGND.n216 VGND.t5143 8.51132
R18451 VGND.n218 VGND.t546 8.51132
R18452 VGND.n220 VGND.t5177 8.51132
R18453 VGND.n222 VGND.t5130 8.51132
R18454 VGND.n224 VGND.t1236 8.51132
R18455 VGND.n239 VGND.t4435 8.51132
R18456 VGND.n237 VGND.t1982 8.51132
R18457 VGND.n236 VGND.t2182 8.51132
R18458 VGND.n234 VGND.t2949 8.51132
R18459 VGND.n232 VGND.t1804 8.51132
R18460 VGND.n62 VGND.t2210 8.51132
R18461 VGND.n68 VGND.t1751 8.51132
R18462 VGND.n70 VGND.t545 8.51132
R18463 VGND.n74 VGND.t2320 8.51132
R18464 VGND.n76 VGND.t1318 8.51132
R18465 VGND.n83 VGND.t1173 8.51132
R18466 VGND.n83 VGND.t2495 8.51132
R18467 VGND.n87 VGND.t1111 8.51132
R18468 VGND.n89 VGND.t1080 8.51132
R18469 VGND.n93 VGND.t2624 8.51132
R18470 VGND.n107 VGND.t1626 8.51132
R18471 VGND.n105 VGND.t999 8.51132
R18472 VGND.n101 VGND.t4176 8.51132
R18473 VGND.n99 VGND.t3625 8.51132
R18474 VGND.n97 VGND.t842 8.51132
R18475 VGND.n54 VGND.t3527 8.51132
R18476 VGND.n3460 VGND.t5555 8.51132
R18477 VGND.n3460 VGND.t5857 8.51132
R18478 VGND.n3459 VGND.t4821 8.51132
R18479 VGND.n3459 VGND.t5033 8.51132
R18480 VGND.n3458 VGND.t4946 8.51132
R18481 VGND.n3458 VGND.t336 8.51132
R18482 VGND.n3457 VGND.t6169 8.51132
R18483 VGND.n3457 VGND.t3112 8.51132
R18484 VGND.n3456 VGND.t5236 8.51132
R18485 VGND.n3456 VGND.t4742 8.51132
R18486 VGND.n3455 VGND.t4467 8.51132
R18487 VGND.n3455 VGND.t648 8.51132
R18488 VGND.n3454 VGND.t1866 8.51132
R18489 VGND.n3454 VGND.t2695 8.51132
R18490 VGND.n3453 VGND.t79 8.51132
R18491 VGND.n3453 VGND.t4079 8.51132
R18492 VGND.n3461 VGND.t744 8.51132
R18493 VGND.n96 VGND.t4358 8.51132
R18494 VGND.n98 VGND.t6759 8.51132
R18495 VGND.n100 VGND.t2633 8.51132
R18496 VGND.n102 VGND.t4443 8.51132
R18497 VGND.n103 VGND.t5581 8.51132
R18498 VGND.n106 VGND.t2421 8.51132
R18499 VGND.n108 VGND.t364 8.51132
R18500 VGND.n109 VGND.t6172 8.51132
R18501 VGND.n95 VGND.t3085 8.51132
R18502 VGND.n92 VGND.t431 8.51132
R18503 VGND.n91 VGND.t737 8.51132
R18504 VGND.n88 VGND.t2373 8.51132
R18505 VGND.n86 VGND.t1104 8.51132
R18506 VGND.n85 VGND.t3167 8.51132
R18507 VGND.n82 VGND.t696 8.51132
R18508 VGND.n79 VGND.t6179 8.51132
R18509 VGND.n77 VGND.t6752 8.51132
R18510 VGND.n75 VGND.t5374 8.51132
R18511 VGND.n73 VGND.t3133 8.51132
R18512 VGND.n72 VGND.t1479 8.51132
R18513 VGND.n69 VGND.t649 8.51132
R18514 VGND.n67 VGND.t6763 8.51132
R18515 VGND.n66 VGND.t72 8.51132
R18516 VGND.n64 VGND.t4096 8.51132
R18517 VGND.n229 VGND.t2283 8.51132
R18518 VGND.n230 VGND.t6810 8.51132
R18519 VGND.n233 VGND.t6091 8.51132
R18520 VGND.n235 VGND.t3966 8.51132
R18521 VGND.n215 VGND.t4345 8.51132
R18522 VGND.n214 VGND.t6175 8.51132
R18523 VGND.n1418 VGND.t3323 8.51132
R18524 VGND.n923 VGND.t1617 8.51132
R18525 VGND.n1324 VGND.t4113 8.51132
R18526 VGND.n1330 VGND.t5697 8.51132
R18527 VGND.n1589 VGND.t4093 8.51132
R18528 VGND.n304 VGND.t492 8.51132
R18529 VGND.n304 VGND.t790 8.51132
R18530 VGND.n305 VGND.t2618 8.51132
R18531 VGND.n305 VGND.t5095 8.51132
R18532 VGND.n307 VGND.t5929 8.51132
R18533 VGND.n308 VGND.t2064 8.51132
R18534 VGND.n328 VGND.t2921 8.51132
R18535 VGND.n329 VGND.t2736 8.51132
R18536 VGND.n331 VGND.t5235 8.51132
R18537 VGND.n335 VGND.t3706 8.51132
R18538 VGND.n337 VGND.t3883 8.51132
R18539 VGND.n339 VGND.t4270 8.51132
R18540 VGND.n341 VGND.t5543 8.51132
R18541 VGND.n342 VGND.t4571 8.51132
R18542 VGND.n343 VGND.t5974 8.51132
R18543 VGND.n344 VGND.t1149 8.51132
R18544 VGND.n345 VGND.t4107 8.51132
R18545 VGND.n354 VGND.t4048 8.51132
R18546 VGND.n353 VGND.t1382 8.51132
R18547 VGND.n352 VGND.t3932 8.51132
R18548 VGND.n351 VGND.t1098 8.51132
R18549 VGND.n350 VGND.t6021 8.51132
R18550 VGND.n349 VGND.t3220 8.51132
R18551 VGND.n348 VGND.t5816 8.51132
R18552 VGND.n347 VGND.t2659 8.51132
R18553 VGND.n3696 VGND.t4322 8.51132
R18554 VGND.n3695 VGND.t5019 8.51132
R18555 VGND.n3694 VGND.t5080 8.51132
R18556 VGND.n3693 VGND.t5252 8.51132
R18557 VGND.n3692 VGND.t3555 8.51132
R18558 VGND.n3690 VGND.t5097 8.51132
R18559 VGND.n3689 VGND.t5907 8.51132
R18560 VGND.n3687 VGND.t3049 8.51132
R18561 VGND.n51 VGND.t484 8.51132
R18562 VGND.n51 VGND.t3287 8.51132
R18563 VGND.n50 VGND.t3502 8.51132
R18564 VGND.n50 VGND.t4124 8.51132
R18565 VGND.n49 VGND.t2768 8.51132
R18566 VGND.n49 VGND.t3602 8.51132
R18567 VGND.n48 VGND.t5936 8.51132
R18568 VGND.n48 VGND.t459 8.51132
R18569 VGND.n47 VGND.t2507 8.51132
R18570 VGND.n47 VGND.t1824 8.51132
R18571 VGND.n46 VGND.t4913 8.51132
R18572 VGND.n46 VGND.t1905 8.51132
R18573 VGND.n45 VGND.t3673 8.51132
R18574 VGND.n45 VGND.t3809 8.51132
R18575 VGND.n44 VGND.t687 8.51132
R18576 VGND.n44 VGND.t5322 8.51132
R18577 VGND.n52 VGND.t1238 8.51132
R18578 VGND.n3688 VGND.t1750 8.51132
R18579 VGND.n338 VGND.t4023 8.51132
R18580 VGND.n336 VGND.t1380 8.51132
R18581 VGND.n334 VGND.t300 8.51132
R18582 VGND.n332 VGND.t2738 8.51132
R18583 VGND.n330 VGND.t2077 8.51132
R18584 VGND.n309 VGND.t1619 8.51132
R18585 VGND.n1569 VGND.t5436 8.51132
R18586 VGND.n1571 VGND.t4072 8.51132
R18587 VGND.n1594 VGND.t5037 8.51132
R18588 VGND.n1340 VGND.t2632 8.51132
R18589 VGND.n1342 VGND.t3531 8.51132
R18590 VGND.n1346 VGND.t3529 8.51132
R18591 VGND.n1328 VGND.t2395 8.51132
R18592 VGND.n1326 VGND.t3549 8.51132
R18593 VGND.n1308 VGND.t4904 8.51132
R18594 VGND.n1306 VGND.t3169 8.51132
R18595 VGND.n1275 VGND.t5777 8.51132
R18596 VGND.n1267 VGND.t5210 8.51132
R18597 VGND.n1261 VGND.t2372 8.51132
R18598 VGND.n1259 VGND.t1737 8.51132
R18599 VGND.n1257 VGND.t1836 8.51132
R18600 VGND.n1254 VGND.t4377 8.51132
R18601 VGND.n1253 VGND.t5460 8.51132
R18602 VGND.n1251 VGND.t2766 8.51132
R18603 VGND.n1250 VGND.t344 8.51132
R18604 VGND.n1247 VGND.t5285 8.51132
R18605 VGND.n1623 VGND.t3659 8.51132
R18606 VGND.n1618 VGND.t3312 8.51132
R18607 VGND.n1616 VGND.t5396 8.51132
R18608 VGND.n1614 VGND.t983 8.51132
R18609 VGND.n1606 VGND.t4320 8.51132
R18610 VGND.n1605 VGND.t3609 8.51132
R18611 VGND.n1602 VGND.t5261 8.51132
R18612 VGND.n1601 VGND.t5589 8.51132
R18613 VGND.n1477 VGND.t5220 8.51132
R18614 VGND.n1475 VGND.t920 8.51132
R18615 VGND.n1443 VGND.t3607 8.51132
R18616 VGND.n1558 VGND.t2987 8.51132
R18617 VGND.n1556 VGND.t5866 8.51132
R18618 VGND.n1555 VGND.t3272 8.51132
R18619 VGND.n1551 VGND.t5306 8.51132
R18620 VGND.n1550 VGND.t5008 8.51132
R18621 VGND.n1547 VGND.t5183 8.51132
R18622 VGND.n3403 VGND.t1564 8.51132
R18623 VGND.n3401 VGND.t862 8.51132
R18624 VGND.n3398 VGND.t4230 8.51132
R18625 VGND.n3381 VGND.t2655 8.51132
R18626 VGND.n3381 VGND.t5596 8.51132
R18627 VGND.n208 VGND.t1095 8.51132
R18628 VGND.n208 VGND.t351 8.51132
R18629 VGND.n254 VGND.t3304 8.51132
R18630 VGND.n260 VGND.t3263 8.51132
R18631 VGND.n261 VGND.t5351 8.51132
R18632 VGND.n263 VGND.t2222 8.51132
R18633 VGND.n264 VGND.t451 8.51132
R18634 VGND.n266 VGND.t5695 8.51132
R18635 VGND.n267 VGND.t4602 8.51132
R18636 VGND.n268 VGND.t2342 8.51132
R18637 VGND.n268 VGND.t4476 8.51132
R18638 VGND.n269 VGND.t2066 8.51132
R18639 VGND.n269 VGND.t5561 8.51132
R18640 VGND.n3382 VGND.t3476 8.51132
R18641 VGND.n3404 VGND.t5567 8.51132
R18642 VGND.n3405 VGND.t3186 8.51132
R18643 VGND.n198 VGND.t1786 8.51132
R18644 VGND.n1515 VGND.t3496 8.51132
R18645 VGND.n1533 VGND.t2197 8.51132
R18646 VGND.n1534 VGND.t5017 8.51132
R18647 VGND.n1536 VGND.t386 8.51132
R18648 VGND.n1538 VGND.t5887 8.51132
R18649 VGND.n1604 VGND.t4835 8.51132
R18650 VGND.n1608 VGND.t3930 8.51132
R18651 VGND.n1610 VGND.t6058 8.51132
R18652 VGND.n1612 VGND.t3114 8.51132
R18653 VGND.n1615 VGND.t594 8.51132
R18654 VGND.n1627 VGND.t4169 8.51132
R18655 VGND.n1252 VGND.t5179 8.51132
R18656 VGND.n1256 VGND.t1778 8.51132
R18657 VGND.n1258 VGND.t3005 8.51132
R18658 VGND.n1260 VGND.t3291 8.51132
R18659 VGND.n1262 VGND.t4820 8.51132
R18660 VGND.n1271 VGND.t2306 8.51132
R18661 VGND.n1233 VGND.t3710 8.51132
R18662 VGND.n1229 VGND.t695 8.51132
R18663 VGND.n1221 VGND.t1162 8.51132
R18664 VGND.n1219 VGND.t4875 8.51132
R18665 VGND.n1216 VGND.t3761 8.51132
R18666 VGND.n1214 VGND.t478 8.51132
R18667 VGND.n1212 VGND.t706 8.51132
R18668 VGND.n1633 VGND.t2460 8.51132
R18669 VGND.n1634 VGND.t902 8.51132
R18670 VGND.n1637 VGND.t433 8.51132
R18671 VGND.n1649 VGND.t4421 8.51132
R18672 VGND.n1696 VGND.t4937 8.51132
R18673 VGND.n1699 VGND.t3537 8.51132
R18674 VGND.n1700 VGND.t480 8.51132
R18675 VGND.n1703 VGND.t6799 8.51132
R18676 VGND.n1705 VGND.t3996 8.51132
R18677 VGND.n1706 VGND.t3821 8.51132
R18678 VGND.n1715 VGND.t3014 8.51132
R18679 VGND.n1714 VGND.t1701 8.51132
R18680 VGND.n1714 VGND.t494 8.51132
R18681 VGND.n1713 VGND.t1796 8.51132
R18682 VGND.n1713 VGND.t5999 8.51132
R18683 VGND.n1712 VGND.t5961 8.51132
R18684 VGND.n1712 VGND.t5241 8.51132
R18685 VGND.n1711 VGND.t1472 8.51132
R18686 VGND.n1711 VGND.t908 8.51132
R18687 VGND.n1790 VGND.t4727 8.51132
R18688 VGND.n1790 VGND.t1992 8.51132
R18689 VGND.n1788 VGND.t3212 8.51132
R18690 VGND.n1777 VGND.t5996 8.51132
R18691 VGND.n1776 VGND.t3634 8.51132
R18692 VGND.n1761 VGND.t4782 8.51132
R18693 VGND.n1759 VGND.t681 8.51132
R18694 VGND.n1749 VGND.t2297 8.51132
R18695 VGND.n1747 VGND.t5060 8.51132
R18696 VGND.n1746 VGND.t5836 8.51132
R18697 VGND.n3374 VGND.t3034 8.51132
R18698 VGND.n3372 VGND.t3306 8.51132
R18699 VGND.n3370 VGND.t5998 8.51132
R18700 VGND.n3367 VGND.t2024 8.51132
R18701 VGND.n3367 VGND.t4751 8.51132
R18702 VGND.n3366 VGND.t1409 8.51132
R18703 VGND.n3366 VGND.t2071 8.51132
R18704 VGND.n3365 VGND.t5679 8.51132
R18705 VGND.n3365 VGND.t2125 8.51132
R18706 VGND.n3364 VGND.t2550 8.51132
R18707 VGND.n3364 VGND.t2492 8.51132
R18708 VGND.n3363 VGND.t3462 8.51132
R18709 VGND.n3363 VGND.t2295 8.51132
R18710 VGND.n3362 VGND.t4829 8.51132
R18711 VGND.n3362 VGND.t5058 8.51132
R18712 VGND.n3361 VGND.t661 8.51132
R18713 VGND.n3361 VGND.t3363 8.51132
R18714 VGND.n3360 VGND.t2218 8.51132
R18715 VGND.n3360 VGND.t5480 8.51132
R18716 VGND.n3368 VGND.t2653 8.51132
R18717 VGND.n3371 VGND.t5952 8.51132
R18718 VGND.n3373 VGND.t3975 8.51132
R18719 VGND.n3375 VGND.t5114 8.51132
R18720 VGND.n3376 VGND.t600 8.51132
R18721 VGND.n1735 VGND.t5563 8.51132
R18722 VGND.n1737 VGND.t5377 8.51132
R18723 VGND.n1738 VGND.t5254 8.51132
R18724 VGND.n1740 VGND.t5308 8.51132
R18725 VGND.n1743 VGND.t2145 8.51132
R18726 VGND.n1745 VGND.t5317 8.51132
R18727 VGND.n1770 VGND.t346 8.51132
R18728 VGND.n1775 VGND.t1554 8.51132
R18729 VGND.n1683 VGND.t2787 8.51132
R18730 VGND.n1653 VGND.t5505 8.51132
R18731 VGND.n1650 VGND.t3108 8.51132
R18732 VGND.n1648 VGND.t2055 8.51132
R18733 VGND.n1647 VGND.t1623 8.51132
R18734 VGND.n1645 VGND.t4392 8.51132
R18735 VGND.n1636 VGND.t677 8.51132
R18736 VGND.n1120 VGND.t5026 8.51132
R18737 VGND.n1152 VGND.t2704 8.51132
R18738 VGND.n1137 VGND.t3238 8.51132
R18739 VGND.n1137 VGND.t4916 8.51132
R18740 VGND.n1136 VGND.t2075 8.51132
R18741 VGND.n1136 VGND.t4942 8.51132
R18742 VGND.n1135 VGND.t2407 8.51132
R18743 VGND.n1135 VGND.t1330 8.51132
R18744 VGND.n1134 VGND.t2005 8.51132
R18745 VGND.n1134 VGND.t1091 8.51132
R18746 VGND.n1133 VGND.t552 8.51132
R18747 VGND.n1133 VGND.t1363 8.51132
R18748 VGND.n1131 VGND.t5869 8.51132
R18749 VGND.n1129 VGND.t5224 8.51132
R18750 VGND.n746 VGND.t1697 8.51132
R18751 VGND.n1796 VGND.t2490 8.51132
R18752 VGND.n1798 VGND.t4551 8.51132
R18753 VGND.n1801 VGND.t4596 8.51132
R18754 VGND.n1803 VGND.t3885 8.51132
R18755 VGND.n721 VGND.t571 8.51132
R18756 VGND.n721 VGND.t361 8.51132
R18757 VGND.n1868 VGND.t1899 8.51132
R18758 VGND.n1866 VGND.t1307 8.51132
R18759 VGND.n1864 VGND.t4165 8.51132
R18760 VGND.n1862 VGND.t2661 8.51132
R18761 VGND.n1860 VGND.t6093 8.51132
R18762 VGND.n1858 VGND.t1901 8.51132
R18763 VGND.n1856 VGND.t4556 8.51132
R18764 VGND.n1854 VGND.t2293 8.51132
R18765 VGND.n1851 VGND.t2266 8.51132
R18766 VGND.n1849 VGND.t2486 8.51132
R18767 VGND.n1847 VGND.t3797 8.51132
R18768 VGND.n1845 VGND.t312 8.51132
R18769 VGND.n1843 VGND.t6187 8.51132
R18770 VGND.n1840 VGND.t2310 8.51132
R18771 VGND.n1838 VGND.t5337 8.51132
R18772 VGND.n1836 VGND.t4448 8.51132
R18773 VGND.n1834 VGND.t659 8.51132
R18774 VGND.n1831 VGND.t2368 8.51132
R18775 VGND.n1831 VGND.t5740 8.51132
R18776 VGND.n1830 VGND.t524 8.51132
R18777 VGND.n1830 VGND.t6170 8.51132
R18778 VGND.n1829 VGND.t403 8.51132
R18779 VGND.n1829 VGND.t6083 8.51132
R18780 VGND.n1828 VGND.t4477 8.51132
R18781 VGND.n1828 VGND.t1166 8.51132
R18782 VGND.n1827 VGND.t720 8.51132
R18783 VGND.n1827 VGND.t3222 8.51132
R18784 VGND.n1826 VGND.t2744 8.51132
R18785 VGND.n1826 VGND.t4606 8.51132
R18786 VGND.n1825 VGND.t5941 8.51132
R18787 VGND.n1825 VGND.t1250 8.51132
R18788 VGND.n1824 VGND.t1880 8.51132
R18789 VGND.n1824 VGND.t6771 8.51132
R18790 VGND.n1832 VGND.t3390 8.51132
R18791 VGND.n1835 VGND.t1998 8.51132
R18792 VGND.n1837 VGND.t4797 8.51132
R18793 VGND.n1839 VGND.t1739 8.51132
R18794 VGND.n1841 VGND.t1441 8.51132
R18795 VGND.n1844 VGND.t698 8.51132
R18796 VGND.n1846 VGND.t711 8.51132
R18797 VGND.n1848 VGND.t3559 8.51132
R18798 VGND.n1850 VGND.t2406 8.51132
R18799 VGND.n1853 VGND.t54 8.51132
R18800 VGND.n1855 VGND.t5569 8.51132
R18801 VGND.n1857 VGND.t334 8.51132
R18802 VGND.n1859 VGND.t4340 8.51132
R18803 VGND.n1861 VGND.t5440 8.51132
R18804 VGND.n1863 VGND.t3494 8.51132
R18805 VGND.n1865 VGND.t5126 8.51132
R18806 VGND.n1867 VGND.t437 8.51132
R18807 VGND.n1869 VGND.t2955 8.51132
R18808 VGND.n1871 VGND.t1517 8.51132
R18809 VGND.n1872 VGND.t3946 8.51132
R18810 VGND.n1874 VGND.t1103 8.51132
R18811 VGND.n1816 VGND.t1484 8.51132
R18812 VGND.n1820 VGND.t4738 8.51132
R18813 VGND.n1812 VGND.t4843 8.51132
R18814 VGND.n1810 VGND.t4810 8.51132
R18815 VGND.n1809 VGND.t2811 8.51132
R18816 VGND.n1807 VGND.t693 8.51132
R18817 VGND.n1806 VGND.t708 8.51132
R18818 VGND.n765 VGND.t5032 8.51132
R18819 VGND.n764 VGND.t1374 8.51132
R18820 VGND.n762 VGND.t5192 8.51132
R18821 VGND.n761 VGND.t3441 8.51132
R18822 VGND.n1132 VGND.t914 8.51132
R18823 VGND.n1138 VGND.t5586 8.51132
R18824 VGND.n1140 VGND.t4871 8.51132
R18825 VGND.n1142 VGND.t1152 8.51132
R18826 VGND.n1165 VGND.t2620 8.51132
R18827 VGND.n1167 VGND.t1320 8.51132
R18828 VGND.n1174 VGND.t5035 8.51132
R18829 VGND.n1176 VGND.t3270 8.51132
R18830 VGND.n1178 VGND.t4253 8.51132
R18831 VGND.n1180 VGND.t4825 8.51132
R18832 VGND.n1182 VGND.t1471 8.51132
R18833 VGND.n1184 VGND.t750 8.51132
R18834 VGND.n1106 VGND.t3348 8.51132
R18835 VGND.n1101 VGND.t56 8.51132
R18836 VGND.n1098 VGND.t4695 8.51132
R18837 VGND.n1096 VGND.t1002 8.51132
R18838 VGND.n1094 VGND.t5122 8.51132
R18839 VGND.n1092 VGND.t3651 8.51132
R18840 VGND.n1091 VGND.t5155 8.51132
R18841 VGND.n1091 VGND.t2639 8.51132
R18842 VGND.n1089 VGND.t2891 8.51132
R18843 VGND.n1086 VGND.t4990 8.51132
R18844 VGND.n1085 VGND.t5295 8.51132
R18845 VGND.n1078 VGND.t4956 8.51132
R18846 VGND.n576 VGND.t4932 8.51132
R18847 VGND.n576 VGND.t824 8.51132
R18848 VGND.n1991 VGND.t5509 8.51132
R18849 VGND.n1989 VGND.t857 8.51132
R18850 VGND.n1987 VGND.t516 8.51132
R18851 VGND.n637 VGND.t3405 8.51132
R18852 VGND.n1916 VGND.t1586 8.51132
R18853 VGND.n1904 VGND.t2938 8.51132
R18854 VGND.n1902 VGND.t4511 8.51132
R18855 VGND.n1900 VGND.t582 8.51132
R18856 VGND.n1899 VGND.t1856 8.51132
R18857 VGND.n1897 VGND.t2356 8.51132
R18858 VGND.n1895 VGND.t5636 8.51132
R18859 VGND.n1893 VGND.t963 8.51132
R18860 VGND.n1891 VGND.t4787 8.51132
R18861 VGND.n1888 VGND.t4175 8.51132
R18862 VGND.n1886 VGND.t4288 8.51132
R18863 VGND.n1884 VGND.t4381 8.51132
R18864 VGND.n1882 VGND.t1568 8.51132
R18865 VGND.n1880 VGND.t1634 8.51132
R18866 VGND.n720 VGND.t4091 8.51132
R18867 VGND.n718 VGND.t808 8.51132
R18868 VGND.n716 VGND.t1309 8.51132
R18869 VGND.n714 VGND.t5206 8.51132
R18870 VGND.n711 VGND.t3764 8.51132
R18871 VGND.n709 VGND.t4513 8.51132
R18872 VGND.n707 VGND.t6079 8.51132
R18873 VGND.n705 VGND.t4234 8.51132
R18874 VGND.n703 VGND.t1342 8.51132
R18875 VGND.n701 VGND.t1248 8.51132
R18876 VGND.n699 VGND.t3352 8.51132
R18877 VGND.n697 VGND.t3908 8.51132
R18878 VGND.n694 VGND.t4945 8.51132
R18879 VGND.n692 VGND.t3842 8.51132
R18880 VGND.n690 VGND.t5138 8.51132
R18881 VGND.n688 VGND.t5901 8.51132
R18882 VGND.n686 VGND.t1865 8.51132
R18883 VGND.n683 VGND.t691 8.51132
R18884 VGND.n681 VGND.t3535 8.51132
R18885 VGND.n679 VGND.t1529 8.51132
R18886 VGND.n677 VGND.t5099 8.51132
R18887 VGND.n674 VGND.t3412 8.51132
R18888 VGND.n674 VGND.t4446 8.51132
R18889 VGND.n673 VGND.t1614 8.51132
R18890 VGND.n673 VGND.t2826 8.51132
R18891 VGND.n672 VGND.t2364 8.51132
R18892 VGND.n672 VGND.t2696 8.51132
R18893 VGND.n671 VGND.t4597 8.51132
R18894 VGND.n671 VGND.t1562 8.51132
R18895 VGND.n670 VGND.t3213 8.51132
R18896 VGND.n670 VGND.t2301 8.51132
R18897 VGND.n669 VGND.t5878 8.51132
R18898 VGND.n669 VGND.t5063 8.51132
R18899 VGND.n668 VGND.t2344 8.51132
R18900 VGND.n668 VGND.t3661 8.51132
R18901 VGND.n667 VGND.t3978 8.51132
R18902 VGND.n667 VGND.t6033 8.51132
R18903 VGND.n675 VGND.t2258 8.51132
R18904 VGND.n678 VGND.t598 8.51132
R18905 VGND.n680 VGND.t4479 8.51132
R18906 VGND.n682 VGND.t5545 8.51132
R18907 VGND.n684 VGND.t2070 8.51132
R18908 VGND.n687 VGND.t4750 8.51132
R18909 VGND.n689 VGND.t3308 8.51132
R18910 VGND.n691 VGND.t5325 8.51132
R18911 VGND.n693 VGND.t1636 8.51132
R18912 VGND.n696 VGND.t4425 8.51132
R18913 VGND.n698 VGND.t2680 8.51132
R18914 VGND.n700 VGND.t1571 8.51132
R18915 VGND.n702 VGND.t2585 8.51132
R18916 VGND.n704 VGND.t2319 8.51132
R18917 VGND.n706 VGND.t3360 8.51132
R18918 VGND.n708 VGND.t5162 8.51132
R18919 VGND.n710 VGND.t4677 8.51132
R18920 VGND.n712 VGND.t1924 8.51132
R18921 VGND.n715 VGND.t413 8.51132
R18922 VGND.n717 VGND.t5448 8.51132
R18923 VGND.n719 VGND.t3095 8.51132
R18924 VGND.n1879 VGND.t4553 8.51132
R18925 VGND.n1881 VGND.t3461 8.51132
R18926 VGND.n1883 VGND.t2806 8.51132
R18927 VGND.n1885 VGND.t5363 8.51132
R18928 VGND.n1887 VGND.t4492 8.51132
R18929 VGND.n1890 VGND.t1123 8.51132
R18930 VGND.n1892 VGND.t2775 8.51132
R18931 VGND.n1894 VGND.t1981 8.51132
R18932 VGND.n1896 VGND.t4744 8.51132
R18933 VGND.n1898 VGND.t3636 8.51132
R18934 VGND.n1074 VGND.t5263 8.51132
R18935 VGND.n940 VGND.t4246 8.51132
R18936 VGND.n938 VGND.t4675 8.51132
R18937 VGND.n936 VGND.t5842 8.51132
R18938 VGND.n1011 VGND.t876 8.51132
R18939 VGND.n1009 VGND.t1018 8.51132
R18940 VGND.n1006 VGND.t2904 8.51132
R18941 VGND.n1006 VGND.t6804 8.51132
R18942 VGND.n1005 VGND.t5895 8.51132
R18943 VGND.n1005 VGND.t3301 8.51132
R18944 VGND.n1004 VGND.t2900 8.51132
R18945 VGND.n1004 VGND.t2740 8.51132
R18946 VGND.n1003 VGND.t50 8.51132
R18947 VGND.n1003 VGND.t1067 8.51132
R18948 VGND.n1002 VGND.t4135 8.51132
R18949 VGND.n1002 VGND.t2843 8.51132
R18950 VGND.n1001 VGND.t1569 8.51132
R18951 VGND.n1001 VGND.t1023 8.51132
R18952 VGND.n1000 VGND.t5268 8.51132
R18953 VGND.n1000 VGND.t4740 8.51132
R18954 VGND.n999 VGND.t5151 8.51132
R18955 VGND.n999 VGND.t5467 8.51132
R18956 VGND.n997 VGND.t1640 8.51132
R18957 VGND.n995 VGND.t6758 8.51132
R18958 VGND.n963 VGND.t773 8.51132
R18959 VGND.n962 VGND.t2675 8.51132
R18960 VGND.n960 VGND.t3397 8.51132
R18961 VGND.n2186 VGND.t2678 8.51132
R18962 VGND.n2188 VGND.t5157 8.51132
R18963 VGND.n2189 VGND.t6165 8.51132
R18964 VGND.n2191 VGND.t6075 8.51132
R18965 VGND.n2192 VGND.t866 8.51132
R18966 VGND.n2217 VGND.t76 8.51132
R18967 VGND.n2215 VGND.t1979 8.51132
R18968 VGND.n2215 VGND.t1884 8.51132
R18969 VGND.n2214 VGND.t3593 8.51132
R18970 VGND.n2214 VGND.t5874 8.51132
R18971 VGND.n2213 VGND.t4554 8.51132
R18972 VGND.n2213 VGND.t3354 8.51132
R18973 VGND.n2212 VGND.t5379 8.51132
R18974 VGND.n2212 VGND.t2583 8.51132
R18975 VGND.n2211 VGND.t5181 8.51132
R18976 VGND.n2211 VGND.t6088 8.51132
R18977 VGND.n2210 VGND.t3361 8.51132
R18978 VGND.n2210 VGND.t78 8.51132
R18979 VGND.n2209 VGND.t5537 8.51132
R18980 VGND.n2209 VGND.t3867 8.51132
R18981 VGND.n2208 VGND.t1037 8.51132
R18982 VGND.n2208 VGND.t2236 8.51132
R18983 VGND.n2216 VGND.t3889 8.51132
R18984 VGND.n2391 VGND.t2389 8.51132
R18985 VGND.n2397 VGND.t4587 8.51132
R18986 VGND.n2399 VGND.t3233 8.51132
R18987 VGND.n955 VGND.t4274 8.51132
R18988 VGND.n959 VGND.t4543 8.51132
R18989 VGND.n961 VGND.t1970 8.51132
R18990 VGND.n975 VGND.t5819 8.51132
R18991 VGND.n977 VGND.t5620 8.51132
R18992 VGND.n979 VGND.t1547 8.51132
R18993 VGND.n981 VGND.t2141 8.51132
R18994 VGND.n1007 VGND.t5823 8.51132
R18995 VGND.n1010 VGND.t1990 8.51132
R18996 VGND.n1012 VGND.t630 8.51132
R18997 VGND.n937 VGND.t1594 8.51132
R18998 VGND.n939 VGND.t1185 8.51132
R18999 VGND.n941 VGND.t3708 8.51132
R19000 VGND.n2564 VGND.t5000 8.51132
R19001 VGND.n2562 VGND.t1782 8.51132
R19002 VGND.n2560 VGND.t4757 8.51132
R19003 VGND.n2598 VGND.t1368 8.51132
R19004 VGND.n2596 VGND.t1199 8.51132
R19005 VGND.n2594 VGND.t4191 8.51132
R19006 VGND.n2592 VGND.t2623 8.51132
R19007 VGND.n2590 VGND.t3029 8.51132
R19008 VGND.n2587 VGND.t713 8.51132
R19009 VGND.n2585 VGND.t4699 8.51132
R19010 VGND.n2583 VGND.t4203 8.51132
R19011 VGND.n2581 VGND.t2308 8.51132
R19012 VGND.n2579 VGND.t5931 8.51132
R19013 VGND.n2577 VGND.t746 8.51132
R19014 VGND.n2575 VGND.t1082 8.51132
R19015 VGND.n2573 VGND.t4823 8.51132
R19016 VGND.n2570 VGND.t5918 8.51132
R19017 VGND.n2568 VGND.t590 8.51132
R19018 VGND.n2566 VGND.t4615 8.51132
R19019 VGND.n410 VGND.t4143 8.51132
R19020 VGND.n2829 VGND.t1693 8.51132
R19021 VGND.n2831 VGND.t3259 8.51132
R19022 VGND.n2833 VGND.t5772 8.51132
R19023 VGND.n2835 VGND.t5603 8.51132
R19024 VGND.n2837 VGND.t3075 8.51132
R19025 VGND.n2840 VGND.t2577 8.51132
R19026 VGND.n2842 VGND.t2166 8.51132
R19027 VGND.n2844 VGND.t1370 8.51132
R19028 VGND.n2846 VGND.t1201 8.51132
R19029 VGND.n2848 VGND.t4195 8.51132
R19030 VGND.n2850 VGND.t3093 8.51132
R19031 VGND.n2852 VGND.t3261 8.51132
R19032 VGND.n2854 VGND.t3116 8.51132
R19033 VGND.n2861 VGND.t419 8.51132
R19034 VGND.n2859 VGND.t1481 8.51132
R19035 VGND.n2857 VGND.t2527 8.51132
R19036 VGND.n409 VGND.t6019 8.51132
R19037 VGND.n2881 VGND.t3395 8.51132
R19038 VGND.n2879 VGND.t4184 8.51132
R19039 VGND.n2877 VGND.t675 8.51132
R19040 VGND.n2875 VGND.t1757 8.51132
R19041 VGND.n2873 VGND.t4238 8.51132
R19042 VGND.n2870 VGND.t580 8.51132
R19043 VGND.n2870 VGND.t1153 8.51132
R19044 VGND.n2869 VGND.t3949 8.51132
R19045 VGND.n2869 VGND.t3572 8.51132
R19046 VGND.n2868 VGND.t2951 8.51132
R19047 VGND.n2868 VGND.t5275 8.51132
R19048 VGND.n2867 VGND.t1733 8.51132
R19049 VGND.n2867 VGND.t1822 8.51132
R19050 VGND.n2866 VGND.t5471 8.51132
R19051 VGND.n2866 VGND.t342 8.51132
R19052 VGND.n2865 VGND.t4430 8.51132
R19053 VGND.n2865 VGND.t382 8.51132
R19054 VGND.n2864 VGND.t3826 8.51132
R19055 VGND.n2864 VGND.t3045 8.51132
R19056 VGND.n2863 VGND.t5451 8.51132
R19057 VGND.n2863 VGND.t614 8.51132
R19058 VGND.n2871 VGND.t1492 8.51132
R19059 VGND.n2874 VGND.t1761 8.51132
R19060 VGND.n2876 VGND.t3998 8.51132
R19061 VGND.n2878 VGND.t4462 8.51132
R19062 VGND.n2880 VGND.t5957 8.51132
R19063 VGND.n2882 VGND.t3526 8.51132
R19064 VGND.n2856 VGND.t2989 8.51132
R19065 VGND.n2858 VGND.t488 8.51132
R19066 VGND.n2860 VGND.t3667 8.51132
R19067 VGND.n2855 VGND.t1387 8.51132
R19068 VGND.n2853 VGND.t3869 8.51132
R19069 VGND.n2851 VGND.t3657 8.51132
R19070 VGND.n2849 VGND.t5948 8.51132
R19071 VGND.n2847 VGND.t4301 8.51132
R19072 VGND.n2845 VGND.t4445 8.51132
R19073 VGND.n2843 VGND.t3443 8.51132
R19074 VGND.n2841 VGND.t5438 8.51132
R19075 VGND.n2839 VGND.t3474 8.51132
R19076 VGND.n2836 VGND.t4908 8.51132
R19077 VGND.n2834 VGND.t5852 8.51132
R19078 VGND.n2832 VGND.t733 8.51132
R19079 VGND.n2830 VGND.t2105 8.51132
R19080 VGND.n2828 VGND.t3871 8.51132
R19081 VGND.n2565 VGND.t4717 8.51132
R19082 VGND.n2567 VGND.t4134 8.51132
R19083 VGND.n2569 VGND.t2403 8.51132
R19084 VGND.n2572 VGND.t3881 8.51132
R19085 VGND.n2574 VGND.t4666 8.51132
R19086 VGND.n2576 VGND.t3745 8.51132
R19087 VGND.n2578 VGND.t1535 8.51132
R19088 VGND.n2580 VGND.t2370 8.51132
R19089 VGND.n2582 VGND.t2348 8.51132
R19090 VGND.n2584 VGND.t3665 8.51132
R19091 VGND.n2586 VGND.t4293 8.51132
R19092 VGND.n2588 VGND.t2825 8.51132
R19093 VGND.n2591 VGND.t4611 8.51132
R19094 VGND.n2593 VGND.t2651 8.51132
R19095 VGND.n2595 VGND.t4608 8.51132
R19096 VGND.n2597 VGND.t4882 8.51132
R19097 VGND.n2559 VGND.t1157 8.51132
R19098 VGND.n2561 VGND.t1628 8.51132
R19099 VGND.n2563 VGND.t1566 8.51132
R19100 VGND.n2613 VGND.t3079 8.51132
R19101 VGND.n2613 VGND.t4139 8.51132
R19102 VGND.n2614 VGND.t4880 8.51132
R19103 VGND.n2614 VGND.t4943 8.51132
R19104 VGND.n2620 VGND.t4678 8.51132
R19105 VGND.n2620 VGND.t578 8.51132
R19106 VGND.n2619 VGND.t4206 8.51132
R19107 VGND.n2619 VGND.t864 8.51132
R19108 VGND.n2618 VGND.t5601 8.51132
R19109 VGND.n2618 VGND.t5021 8.51132
R19110 VGND.n2617 VGND.t3310 8.51132
R19111 VGND.n2617 VGND.t4102 8.51132
R19112 VGND.n2616 VGND.t3289 8.51132
R19113 VGND.n2616 VGND.t4600 8.51132
R19114 VGND.n2615 VGND.t2233 8.51132
R19115 VGND.n2615 VGND.t4922 8.51132
R19116 VGND.n2612 VGND.t5939 8.51132
R19117 VGND.n2602 VGND.t4058 8.51132
R19118 VGND.n2602 VGND.t1322 8.51132
R19119 VGND.n2603 VGND.t1117 8.51132
R19120 VGND.n2603 VGND.t5477 8.51132
R19121 VGND.n2609 VGND.t5315 8.51132
R19122 VGND.n2609 VGND.t2595 8.51132
R19123 VGND.n2608 VGND.t5925 8.51132
R19124 VGND.n2608 VGND.t5990 8.51132
R19125 VGND.n2607 VGND.t4035 8.51132
R19126 VGND.n2607 VGND.t6171 8.51132
R19127 VGND.n2606 VGND.t2948 8.51132
R19128 VGND.n2606 VGND.t6795 8.51132
R19129 VGND.n2605 VGND.t2700 8.51132
R19130 VGND.n2605 VGND.t5979 8.51132
R19131 VGND.n2604 VGND.t5855 8.51132
R19132 VGND.n2604 VGND.t3472 8.51132
R19133 VGND.n2601 VGND.t3371 8.51132
R19134 VGND.n391 VGND.t4588 8.51132
R19135 VGND.n391 VGND.t4291 8.51132
R19136 VGND.n392 VGND.t3899 8.51132
R19137 VGND.n392 VGND.t3386 8.51132
R19138 VGND.n394 VGND.t2472 8.51132
R19139 VGND.n394 VGND.t5773 8.51132
R19140 VGND.n395 VGND.t1257 8.51132
R19141 VGND.n395 VGND.t834 8.51132
R19142 VGND.n396 VGND.t967 8.51132
R19143 VGND.n396 VGND.t5022 8.51132
R19144 VGND.n397 VGND.t3097 8.51132
R19145 VGND.n397 VGND.t3362 8.51132
R19146 VGND.n398 VGND.t5919 8.51132
R19147 VGND.n398 VGND.t4605 8.51132
R19148 VGND.n399 VGND.t2796 8.51132
R19149 VGND.n399 VGND.t5133 8.51132
R19150 VGND.n390 VGND.t3492 8.51132
R19151 VGND.n386 VGND.t3524 8.51132
R19152 VGND.n386 VGND.t3700 8.51132
R19153 VGND.n385 VGND.t5659 8.51132
R19154 VGND.n385 VGND.t5877 8.51132
R19155 VGND.n2960 VGND.t1794 8.51132
R19156 VGND.n2960 VGND.t3717 8.51132
R19157 VGND.n2959 VGND.t5812 8.51132
R19158 VGND.n2959 VGND.t2641 8.51132
R19159 VGND.n2958 VGND.t4038 8.51132
R19160 VGND.n2958 VGND.t465 8.51132
R19161 VGND.n2957 VGND.t3750 8.51132
R19162 VGND.n2957 VGND.t671 8.51132
R19163 VGND.n2956 VGND.t5611 8.51132
R19164 VGND.n2956 VGND.t2961 8.51132
R19165 VGND.n2955 VGND.t5885 8.51132
R19166 VGND.n2955 VGND.t4549 8.51132
R19167 VGND.n387 VGND.t3702 8.51132
R19168 VGND.n413 VGND.t3173 8.51132
R19169 VGND.n415 VGND.t4037 8.51132
R19170 VGND.n417 VGND.t2030 8.51132
R19171 VGND.n2733 VGND.t979 8.51132
R19172 VGND.n2735 VGND.t1175 8.51132
R19173 VGND.n2737 VGND.t2756 8.51132
R19174 VGND.n2739 VGND.t1044 8.51132
R19175 VGND.n2741 VGND.t5627 8.51132
R19176 VGND.n2744 VGND.t5327 8.51132
R19177 VGND.n2746 VGND.t3713 8.51132
R19178 VGND.n2748 VGND.t4272 8.51132
R19179 VGND.n2750 VGND.t1531 8.51132
R19180 VGND.n2752 VGND.t5381 8.51132
R19181 VGND.n2754 VGND.t4793 8.51132
R19182 VGND.n2756 VGND.t2366 8.51132
R19183 VGND.n2758 VGND.t4089 8.51132
R19184 VGND.n2765 VGND.t5347 8.51132
R19185 VGND.n2763 VGND.t5011 8.51132
R19186 VGND.n2761 VGND.t5889 8.51132
R19187 VGND.n412 VGND.t3844 8.51132
R19188 VGND.n2822 VGND.t3120 8.51132
R19189 VGND.n2820 VGND.t1344 8.51132
R19190 VGND.n2818 VGND.t3439 8.51132
R19191 VGND.n2816 VGND.t3551 8.51132
R19192 VGND.n2814 VGND.t3392 8.51132
R19193 VGND.n2811 VGND.t3855 8.51132
R19194 VGND.n2809 VGND.t5830 8.51132
R19195 VGND.n2807 VGND.t5247 8.51132
R19196 VGND.n2805 VGND.t4892 8.51132
R19197 VGND.n2803 VGND.t5960 8.51132
R19198 VGND.n2801 VGND.t52 8.51132
R19199 VGND.n2799 VGND.t3586 8.51132
R19200 VGND.n2797 VGND.t1577 8.51132
R19201 VGND.n2794 VGND.t4379 8.51132
R19202 VGND.n2792 VGND.t4764 8.51132
R19203 VGND.n2790 VGND.t669 8.51132
R19204 VGND.n2788 VGND.t4726 8.51132
R19205 VGND.n2785 VGND.t3206 8.51132
R19206 VGND.n2783 VGND.t5801 8.51132
R19207 VGND.n2781 VGND.t3012 8.51132
R19208 VGND.n2779 VGND.t5104 8.51132
R19209 VGND.n2777 VGND.t2702 8.51132
R19210 VGND.n2774 VGND.t4567 8.51132
R19211 VGND.n2774 VGND.t1815 8.51132
R19212 VGND.n2773 VGND.t5039 8.51132
R19213 VGND.n2773 VGND.t5271 8.51132
R19214 VGND.n2772 VGND.t4369 8.51132
R19215 VGND.n2772 VGND.t1525 8.51132
R19216 VGND.n2771 VGND.t3896 8.51132
R19217 VGND.n2771 VGND.t2928 8.51132
R19218 VGND.n2770 VGND.t1340 8.51132
R19219 VGND.n2770 VGND.t6059 8.51132
R19220 VGND.n2769 VGND.t2340 8.51132
R19221 VGND.n2769 VGND.t3236 8.51132
R19222 VGND.n2768 VGND.t3038 8.51132
R19223 VGND.n2768 VGND.t5535 8.51132
R19224 VGND.n2767 VGND.t3218 8.51132
R19225 VGND.n2767 VGND.t3757 8.51132
R19226 VGND.n2775 VGND.t548 8.51132
R19227 VGND.n2778 VGND.t1332 8.51132
R19228 VGND.n2780 VGND.t1211 8.51132
R19229 VGND.n2782 VGND.t4357 8.51132
R19230 VGND.n2784 VGND.t1223 8.51132
R19231 VGND.n2786 VGND.t1658 8.51132
R19232 VGND.n2789 VGND.t5408 8.51132
R19233 VGND.n2791 VGND.t2190 8.51132
R19234 VGND.n2793 VGND.t2350 8.51132
R19235 VGND.n2796 VGND.t3570 8.51132
R19236 VGND.n2798 VGND.t534 8.51132
R19237 VGND.n2800 VGND.t5718 8.51132
R19238 VGND.n2802 VGND.t2326 8.51132
R19239 VGND.n2804 VGND.t673 8.51132
R19240 VGND.n2806 VGND.t4771 8.51132
R19241 VGND.n2808 VGND.t3036 8.51132
R19242 VGND.n2810 VGND.t5075 8.51132
R19243 VGND.n2812 VGND.t1819 8.51132
R19244 VGND.n2815 VGND.t5839 8.51132
R19245 VGND.n2817 VGND.t2886 8.51132
R19246 VGND.n2819 VGND.t4450 8.51132
R19247 VGND.n2821 VGND.t5187 8.51132
R19248 VGND.n2823 VGND.t4659 8.51132
R19249 VGND.n2760 VGND.t3994 8.51132
R19250 VGND.n2762 VGND.t3020 8.51132
R19251 VGND.n2764 VGND.t1338 8.51132
R19252 VGND.n2759 VGND.t5803 8.51132
R19253 VGND.n2757 VGND.t4398 8.51132
R19254 VGND.n2755 VGND.t2091 8.51132
R19255 VGND.n2753 VGND.t1834 8.51132
R19256 VGND.n2751 VGND.t785 8.51132
R19257 VGND.n2749 VGND.t3715 8.51132
R19258 VGND.n2747 VGND.t496 8.51132
R19259 VGND.n2745 VGND.t4711 8.51132
R19260 VGND.n2743 VGND.t2324 8.51132
R19261 VGND.n2740 VGND.t1958 8.51132
R19262 VGND.n2738 VGND.t3799 8.51132
R19263 VGND.n2736 VGND.t5648 8.51132
R19264 VGND.n2734 VGND.t1357 8.51132
R19265 VGND.n418 VGND.t1467 8.51132
R19266 VGND.n416 VGND.t5826 8.51132
R19267 VGND.n414 VGND.t3171 8.51132
R19268 VGND.n2624 VGND.t3399 8.51132
R19269 VGND.n2627 VGND.t5106 8.51132
R19270 VGND.n2625 VGND.t2790 8.51132
R19271 VGND.n2728 VGND.t5469 8.51132
R19272 VGND.n2726 VGND.t3231 8.51132
R19273 VGND.n2724 VGND.t814 8.51132
R19274 VGND.n2722 VGND.t5004 8.51132
R19275 VGND.n2720 VGND.t2899 8.51132
R19276 VGND.n2716 VGND.t463 8.51132
R19277 VGND.n2714 VGND.t6816 8.51132
R19278 VGND.n2712 VGND.t6768 8.51132
R19279 VGND.n2710 VGND.t380 8.51132
R19280 VGND.n2708 VGND.t4780 8.51132
R19281 VGND.n2706 VGND.t4212 8.51132
R19282 VGND.n2704 VGND.t2123 8.51132
R19283 VGND.n2702 VGND.t2287 8.51132
R19284 VGND.n2700 VGND.t4953 8.51132
R19285 VGND.n2697 VGND.t2657 8.51132
R19286 VGND.n2695 VGND.t6803 8.51132
R19287 VGND.n2693 VGND.t3184 8.51132
R19288 VGND.n2690 VGND.t4305 8.51132
R19289 VGND.n2688 VGND.t4483 8.51132
R19290 VGND.n2686 VGND.t2148 8.51132
R19291 VGND.n2684 VGND.t2304 8.51132
R19292 VGND.n2682 VGND.t1996 8.51132
R19293 VGND.n2679 VGND.t5557 8.51132
R19294 VGND.n2677 VGND.t1677 8.51132
R19295 VGND.n2675 VGND.t1598 8.51132
R19296 VGND.n2673 VGND.t1197 8.51132
R19297 VGND.n2671 VGND.t792 8.51132
R19298 VGND.n2669 VGND.t4488 8.51132
R19299 VGND.n2667 VGND.t1916 8.51132
R19300 VGND.n2665 VGND.t3384 8.51132
R19301 VGND.n2663 VGND.t3188 8.51132
R19302 VGND.n2661 VGND.t3638 8.51132
R19303 VGND.n2659 VGND.t5270 8.51132
R19304 VGND.n2657 VGND.t5319 8.51132
R19305 VGND.n2654 VGND.t5731 8.51132
R19306 VGND.n2652 VGND.t1600 8.51132
R19307 VGND.n2650 VGND.t66 8.51132
R19308 VGND.n2648 VGND.t6041 8.51132
R19309 VGND.n2646 VGND.t6174 8.51132
R19310 VGND.n2642 VGND.t5513 8.51132
R19311 VGND.n2642 VGND.t5867 8.51132
R19312 VGND.n2641 VGND.t2334 8.51132
R19313 VGND.n2641 VGND.t4015 8.51132
R19314 VGND.n2640 VGND.t1288 8.51132
R19315 VGND.n2640 VGND.t4728 8.51132
R19316 VGND.n2639 VGND.t5112 8.51132
R19317 VGND.n2639 VGND.t3704 8.51132
R19318 VGND.n2638 VGND.t2558 8.51132
R19319 VGND.n2638 VGND.t3976 8.51132
R19320 VGND.n2637 VGND.t3898 8.51132
R19321 VGND.n2637 VGND.t6178 8.51132
R19322 VGND.n2636 VGND.t5116 8.51132
R19323 VGND.n2636 VGND.t1155 8.51132
R19324 VGND.n2635 VGND.t1740 8.51132
R19325 VGND.n2635 VGND.t340 8.51132
R19326 VGND.n2645 VGND.t5145 8.51132
R19327 VGND.n2647 VGND.t500 8.51132
R19328 VGND.n2649 VGND.t5978 8.51132
R19329 VGND.n2651 VGND.t3143 8.51132
R19330 VGND.n2653 VGND.t1711 8.51132
R19331 VGND.n2656 VGND.t5453 8.51132
R19332 VGND.n2658 VGND.t4503 8.51132
R19333 VGND.n2660 VGND.t1844 8.51132
R19334 VGND.n2664 VGND.t3793 8.51132
R19335 VGND.n2666 VGND.t1433 8.51132
R19336 VGND.n2668 VGND.t5862 8.51132
R19337 VGND.n2670 VGND.t5575 8.51132
R19338 VGND.n2672 VGND.t5202 8.51132
R19339 VGND.n2674 VGND.t4831 8.51132
R19340 VGND.n2676 VGND.t3928 8.51132
R19341 VGND.n2678 VGND.t1048 8.51132
R19342 VGND.n2680 VGND.t3369 8.51132
R19343 VGND.n2683 VGND.t435 8.51132
R19344 VGND.n2685 VGND.t1478 8.51132
R19345 VGND.n2687 VGND.t4715 8.51132
R19346 VGND.n2689 VGND.t1988 8.51132
R19347 VGND.n2691 VGND.t1282 8.51132
R19348 VGND.n2694 VGND.t5065 8.51132
R19349 VGND.n2696 VGND.t4216 8.51132
R19350 VGND.n2699 VGND.t5595 8.51132
R19351 VGND.n2701 VGND.t2216 8.51132
R19352 VGND.n2703 VGND.t4928 8.51132
R19353 VGND.n2705 VGND.t3647 8.51132
R19354 VGND.n2707 VGND.t1108 8.51132
R19355 VGND.n2709 VGND.t4250 8.51132
R19356 VGND.n2711 VGND.t2720 8.51132
R19357 VGND.n2713 VGND.t4851 8.51132
R19358 VGND.n2717 VGND.t5450 8.51132
R19359 VGND.n2719 VGND.t1389 8.51132
R19360 VGND.n2721 VGND.t1277 8.51132
R19361 VGND.n2723 VGND.t959 8.51132
R19362 VGND.n2725 VGND.t5739 8.51132
R19363 VGND.n2727 VGND.t1798 8.51132
R19364 VGND.n2623 VGND.t4475 8.51132
R19365 VGND.n2626 VGND.t3857 8.51132
R19366 VGND.n430 VGND.t1592 8.51132
R19367 VGND.n432 VGND.t1638 8.51132
R19368 VGND.n434 VGND.t2410 8.51132
R19369 VGND.n437 VGND.t1893 8.51132
R19370 VGND.n439 VGND.t3918 8.51132
R19371 VGND.n442 VGND.t3968 8.51132
R19372 VGND.n442 VGND.t5154 8.51132
R19373 VGND.n443 VGND.t1763 8.51132
R19374 VGND.n443 VGND.t2146 8.51132
R19375 VGND.n444 VGND.t2926 8.51132
R19376 VGND.n444 VGND.t1644 8.51132
R19377 VGND.n445 VGND.t554 8.51132
R19378 VGND.n445 VGND.t4951 8.51132
R19379 VGND.n446 VGND.t702 8.51132
R19380 VGND.n446 VGND.t1895 8.51132
R19381 VGND.n447 VGND.t5548 8.51132
R19382 VGND.n447 VGND.t3920 8.51132
R19383 VGND.n448 VGND.t5712 8.51132
R19384 VGND.n448 VGND.t3719 8.51132
R19385 VGND.n449 VGND.t965 8.51132
R19386 VGND.n449 VGND.t6180 8.51132
R19387 VGND.n464 VGND.t3916 8.51132
R19388 VGND.n2443 VGND.t4266 8.51132
R19389 VGND.n2440 VGND.t3240 8.51132
R19390 VGND.n2440 VGND.t4776 8.51132
R19391 VGND.n2439 VGND.t3649 8.51132
R19392 VGND.n2439 VGND.t5153 8.51132
R19393 VGND.n2438 VGND.t2036 8.51132
R19394 VGND.n2438 VGND.t6060 8.51132
R19395 VGND.n2430 VGND.t5239 8.51132
R19396 VGND.n2428 VGND.t4490 8.51132
R19397 VGND.n2426 VGND.t1918 8.51132
R19398 VGND.n2424 VGND.t3388 8.51132
R19399 VGND.n2422 VGND.t1527 8.51132
R19400 VGND.n2420 VGND.t1203 8.51132
R19401 VGND.n2418 VGND.t2501 8.51132
R19402 VGND.n2416 VGND.t5321 8.51132
R19403 VGND.n2414 VGND.t4101 8.51132
R19404 VGND.n488 VGND.t1360 8.51132
R19405 VGND.n490 VGND.t4197 8.51132
R19406 VGND.n494 VGND.t3777 8.51132
R19407 VGND.n496 VGND.t2841 8.51132
R19408 VGND.n498 VGND.t6182 8.51132
R19409 VGND.n500 VGND.t2718 8.51132
R19410 VGND.n502 VGND.t4812 8.51132
R19411 VGND.n504 VGND.t4371 8.51132
R19412 VGND.n506 VGND.t3490 8.51132
R19413 VGND.n519 VGND.t1235 8.51132
R19414 VGND.n518 VGND.t4642 8.51132
R19415 VGND.n2355 VGND.t2235 8.51132
R19416 VGND.n2353 VGND.t765 8.51132
R19417 VGND.n546 VGND.t5110 8.51132
R19418 VGND.n544 VGND.t4138 8.51132
R19419 VGND.n542 VGND.t561 8.51132
R19420 VGND.n539 VGND.t5442 8.51132
R19421 VGND.n539 VGND.t5565 8.51132
R19422 VGND.n538 VGND.t977 8.51132
R19423 VGND.n538 VGND.t2616 8.51132
R19424 VGND.n537 VGND.t4884 8.51132
R19425 VGND.n537 VGND.t6770 8.51132
R19426 VGND.n536 VGND.t4984 8.51132
R19427 VGND.n536 VGND.t5612 8.51132
R19428 VGND.n535 VGND.t2771 8.51132
R19429 VGND.n535 VGND.t4289 8.51132
R19430 VGND.n534 VGND.t5940 8.51132
R19431 VGND.n534 VGND.t5650 8.51132
R19432 VGND.n533 VGND.t1940 8.51132
R19433 VGND.n533 VGND.t2823 8.51132
R19434 VGND.n532 VGND.t2198 8.51132
R19435 VGND.n532 VGND.t1401 8.51132
R19436 VGND.n540 VGND.t3244 8.51132
R19437 VGND.n543 VGND.t5128 8.51132
R19438 VGND.n545 VGND.t4427 8.51132
R19439 VGND.n547 VGND.t1417 8.51132
R19440 VGND.n2354 VGND.t2043 8.51132
R19441 VGND.n2356 VGND.t592 8.51132
R19442 VGND.n2357 VGND.t2317 8.51132
R19443 VGND.n2359 VGND.t573 8.51132
R19444 VGND.n2361 VGND.t1486 8.51132
R19445 VGND.n2366 VGND.t4104 8.51132
R19446 VGND.n512 VGND.t679 8.51132
R19447 VGND.n513 VGND.t5714 8.51132
R19448 VGND.n515 VGND.t5174 8.51132
R19449 VGND.n517 VGND.t576 8.51132
R19450 VGND.n507 VGND.t5249 8.51132
R19451 VGND.n505 VGND.t5846 8.51132
R19452 VGND.n503 VGND.t2694 8.51132
R19453 VGND.n501 VGND.t2910 8.51132
R19454 VGND.n499 VGND.t5343 8.51132
R19455 VGND.n497 VGND.t756 8.51132
R19456 VGND.n495 VGND.t5160 8.51132
R19457 VGND.n493 VGND.t5724 8.51132
R19458 VGND.n492 VGND.t4171 8.51132
R19459 VGND.n489 VGND.t3819 8.51132
R19460 VGND.n468 VGND.t1437 8.51132
R19461 VGND.n2415 VGND.t3561 8.51132
R19462 VGND.n2417 VGND.t5848 8.51132
R19463 VGND.n2419 VGND.t729 8.51132
R19464 VGND.n2421 VGND.t563 8.51132
R19465 VGND.n2423 VGND.t2068 8.51132
R19466 VGND.n2425 VGND.t2581 8.51132
R19467 VGND.n2441 VGND.t6044 8.51132
R19468 VGND.n2444 VGND.t3901 8.51132
R19469 VGND.n2445 VGND.t3629 8.51132
R19470 VGND.n462 VGND.t359 8.51132
R19471 VGND.n441 VGND.t3242 8.51132
R19472 VGND.n438 VGND.t655 8.51132
R19473 VGND.n436 VGND.t4873 8.51132
R19474 VGND.n433 VGND.t1974 8.51132
R19475 VGND.n431 VGND.t2637 8.51132
R19476 VGND.n429 VGND.t4785 8.51132
R19477 VGND.n424 VGND.t6185 8.51132
R19478 VGND.n422 VGND.t6167 8.51132
R19479 VGND.n420 VGND.t1725 8.51132
R19480 VGND.n2485 VGND.t3099 8.51132
R19481 VGND.n2483 VGND.t1826 8.51132
R19482 VGND.n2480 VGND.t5078 8.51132
R19483 VGND.n2478 VGND.t1279 8.51132
R19484 VGND.n2476 VGND.t2290 8.51132
R19485 VGND.n2474 VGND.t2051 8.51132
R19486 VGND.n2472 VGND.t2264 8.51132
R19487 VGND.n2470 VGND.t851 8.51132
R19488 VGND.n2468 VGND.t319 8.51132
R19489 VGND.n2466 VGND.t4697 8.51132
R19490 VGND.n2463 VGND.t5194 8.51132
R19491 VGND.n2462 VGND.t3025 8.51132
R19492 VGND.n2462 VGND.t5123 8.51132
R19493 VGND.n2224 VGND.t6749 8.51132
R19494 VGND.n2226 VGND.t4481 8.51132
R19495 VGND.n2230 VGND.t3624 8.51132
R19496 VGND.n2243 VGND.t1832 8.51132
R19497 VGND.n2245 VGND.t992 8.51132
R19498 VGND.n2248 VGND.t6809 8.51132
R19499 VGND.n2250 VGND.t6766 8.51132
R19500 VGND.n2252 VGND.t4508 8.51132
R19501 VGND.n2254 VGND.t3274 8.51132
R19502 VGND.n2256 VGND.t5681 8.51132
R19503 VGND.n2258 VGND.t2566 8.51132
R19504 VGND.n2260 VGND.t504 8.51132
R19505 VGND.n2263 VGND.t5314 8.51132
R19506 VGND.n2265 VGND.t4429 8.51132
R19507 VGND.n2268 VGND.t1020 8.51132
R19508 VGND.n2270 VGND.t3622 8.51132
R19509 VGND.n2272 VGND.t3807 8.51132
R19510 VGND.n2274 VGND.t1581 8.51132
R19511 VGND.n2276 VGND.t1560 8.51132
R19512 VGND.n2278 VGND.t6751 8.51132
R19513 VGND.n2280 VGND.t4622 8.51132
R19514 VGND.n2282 VGND.t602 8.51132
R19515 VGND.n2285 VGND.t2205 8.51132
R19516 VGND.n2287 VGND.t1125 8.51132
R19517 VGND.n2289 VGND.t1886 8.51132
R19518 VGND.n2291 VGND.t6077 8.51132
R19519 VGND.n2293 VGND.t4330 8.51132
R19520 VGND.n2295 VGND.t4432 8.51132
R19521 VGND.n2298 VGND.t2152 8.51132
R19522 VGND.n2300 VGND.t1004 8.51132
R19523 VGND.n2302 VGND.t1284 8.51132
R19524 VGND.n2305 VGND.t1494 8.51132
R19525 VGND.n2307 VGND.t3671 8.51132
R19526 VGND.n2309 VGND.t5541 8.51132
R19527 VGND.n2311 VGND.t1964 8.51132
R19528 VGND.n2313 VGND.t1439 8.51132
R19529 VGND.n2315 VGND.t4613 8.51132
R19530 VGND.n2317 VGND.t1393 8.51132
R19531 VGND.n2319 VGND.t6797 8.51132
R19532 VGND.n2330 VGND.t853 8.51132
R19533 VGND.n2328 VGND.t4115 8.51132
R19534 VGND.n2326 VGND.t5550 8.51132
R19535 VGND.n2324 VGND.t2186 8.51132
R19536 VGND.n2322 VGND.t3574 8.51132
R19537 VGND.n2222 VGND.t2004 8.51132
R19538 VGND.n2347 VGND.t800 8.51132
R19539 VGND.n2345 VGND.t1942 8.51132
R19540 VGND.n2343 VGND.t3914 8.51132
R19541 VGND.n2340 VGND.t1914 8.51132
R19542 VGND.n2340 VGND.t1133 8.51132
R19543 VGND.n2339 VGND.t1280 8.51132
R19544 VGND.n2339 VGND.t405 8.51132
R19545 VGND.n2338 VGND.t3830 8.51132
R19546 VGND.n2338 VGND.t3547 8.51132
R19547 VGND.n2337 VGND.t4095 8.51132
R19548 VGND.n2337 VGND.t4149 8.51132
R19549 VGND.n2336 VGND.t2878 8.51132
R19550 VGND.n2336 VGND.t4011 8.51132
R19551 VGND.n2335 VGND.t1431 8.51132
R19552 VGND.n2335 VGND.t1842 8.51132
R19553 VGND.n2334 VGND.t4111 8.51132
R19554 VGND.n2334 VGND.t5198 8.51132
R19555 VGND.n2333 VGND.t1476 8.51132
R19556 VGND.n2333 VGND.t910 8.51132
R19557 VGND.n2341 VGND.t4040 8.51132
R19558 VGND.n2344 VGND.t1872 8.51132
R19559 VGND.n2346 VGND.t3721 8.51132
R19560 VGND.n2348 VGND.t4915 8.51132
R19561 VGND.n2321 VGND.t1496 8.51132
R19562 VGND.n2323 VGND.t1648 8.51132
R19563 VGND.n2325 VGND.t3743 8.51132
R19564 VGND.n2327 VGND.t5360 8.51132
R19565 VGND.n2329 VGND.t3627 8.51132
R19566 VGND.n2320 VGND.t2499 8.51132
R19567 VGND.n2318 VGND.t2256 8.51132
R19568 VGND.n2316 VGND.t2575 8.51132
R19569 VGND.n2314 VGND.t1952 8.51132
R19570 VGND.n2312 VGND.t3578 8.51132
R19571 VGND.n2310 VGND.t2312 8.51132
R19572 VGND.n2308 VGND.t4156 8.51132
R19573 VGND.n2306 VGND.t2792 8.51132
R19574 VGND.n2304 VGND.t415 8.51132
R19575 VGND.n2301 VGND.t4877 8.51132
R19576 VGND.n2299 VGND.t2111 8.51132
R19577 VGND.n2296 VGND.t2079 8.51132
R19578 VGND.n2294 VGND.t4189 8.51132
R19579 VGND.n2292 VGND.t5876 8.51132
R19580 VGND.n2290 VGND.t4351 8.51132
R19581 VGND.n2288 VGND.t1094 8.51132
R19582 VGND.n2286 VGND.t5434 8.51132
R19583 VGND.n2283 VGND.t3988 8.51132
R19584 VGND.n2281 VGND.t4795 8.51132
R19585 VGND.n2279 VGND.t1490 8.51132
R19586 VGND.n2277 VGND.t1445 8.51132
R19587 VGND.n2275 VGND.t1550 8.51132
R19588 VGND.n2273 VGND.t5358 8.51132
R19589 VGND.n2271 VGND.t1715 8.51132
R19590 VGND.n2269 VGND.t941 8.51132
R19591 VGND.n2267 VGND.t1397 8.51132
R19592 VGND.n2264 VGND.t4988 8.51132
R19593 VGND.n2262 VGND.t4766 8.51132
R19594 VGND.n2259 VGND.t796 8.51132
R19595 VGND.n2257 VGND.t5522 8.51132
R19596 VGND.n2255 VGND.t1415 8.51132
R19597 VGND.n2253 VGND.t5669 8.51132
R19598 VGND.n2251 VGND.t4220 8.51132
R19599 VGND.n2249 VGND.t4581 8.51132
R19600 VGND.n2246 VGND.t4547 8.51132
R19601 VGND.n2244 VGND.t2635 8.51132
R19602 VGND.n2242 VGND.t5226 8.51132
R19603 VGND.n2460 VGND.t5625 8.51132
R19604 VGND.n2465 VGND.t3663 8.51132
R19605 VGND.n2467 VGND.t794 8.51132
R19606 VGND.n2469 VGND.t2543 8.51132
R19607 VGND.n2471 VGND.t5094 8.51132
R19608 VGND.n2473 VGND.t5654 8.51132
R19609 VGND.n2475 VGND.t4218 8.51132
R19610 VGND.n2477 VGND.t4470 8.51132
R19611 VGND.n2479 VGND.t4141 8.51132
R19612 VGND.n2481 VGND.t398 8.51132
R19613 VGND.n2484 VGND.t5971 8.51132
R19614 VGND.n2486 VGND.t2934 8.51132
R19615 VGND.n421 VGND.t618 8.51132
R19616 VGND.n423 VGND.t5678 8.51132
R19617 VGND.n425 VGND.t6052 8.51132
R19618 VGND.n2491 VGND.t4044 8.51132
R19619 VGND.n2491 VGND.t3922 8.51132
R19620 VGND.n2490 VGND.t2037 8.51132
R19621 VGND.n2490 VGND.t969 8.51132
R19622 VGND.n2489 VGND.t880 8.51132
R19623 VGND.n2489 VGND.t2985 8.51132
R19624 VGND.n2556 VGND.t5024 8.51132
R19625 VGND.n2556 VGND.t5328 8.51132
R19626 VGND.n2555 VGND.t1687 8.51132
R19627 VGND.n2555 VGND.t727 8.51132
R19628 VGND.n2554 VGND.t3617 8.51132
R19629 VGND.n2554 VGND.t5491 8.51132
R19630 VGND.n2553 VGND.t5479 8.51132
R19631 VGND.n2553 VGND.t5716 8.51132
R19632 VGND.n2550 VGND.t1846 8.51132
R19633 VGND.n2548 VGND.t5108 8.51132
R19634 VGND.n2546 VGND.t3904 8.51132
R19635 VGND.n2544 VGND.t4248 8.51132
R19636 VGND.n2542 VGND.t5486 8.51132
R19637 VGND.n2540 VGND.t704 8.51132
R19638 VGND.n2538 VGND.t5458 8.51132
R19639 VGND.n2536 VGND.t2671 8.51132
R19640 VGND.n2512 VGND.t1806 8.51132
R19641 VGND.n2512 VGND.t4509 8.51132
R19642 VGND.n2511 VGND.t1066 8.51132
R19643 VGND.n2511 VGND.t5296 8.51132
R19644 VGND.n2510 VGND.t3067 8.51132
R19645 VGND.n2510 VGND.t5892 8.51132
R19646 VGND.n2509 VGND.t4769 8.51132
R19647 VGND.n2509 VGND.t2160 8.51132
R19648 VGND.n2508 VGND.t447 8.51132
R19649 VGND.n2508 VGND.t5069 8.51132
R19650 VGND.n2507 VGND.t5560 8.51132
R19651 VGND.n2507 VGND.t961 8.51132
R19652 VGND.n2506 VGND.t4010 8.51132
R19653 VGND.n2506 VGND.t1372 8.51132
R19654 VGND.n2505 VGND.t5604 8.51132
R19655 VGND.n2505 VGND.t376 8.51132
R19656 VGND.n2501 VGND.t2856 8.51132
R19657 VGND.n2500 VGND.t498 8.51132
R19658 VGND.n2500 VGND.t6801 8.51132
R19659 VGND.n2499 VGND.t3452 8.51132
R19660 VGND.n2499 VGND.t3182 8.51132
R19661 VGND.n2498 VGND.t4741 8.51132
R19662 VGND.n2498 VGND.t4303 8.51132
R19663 VGND.n2887 VGND.t4078 8.51132
R19664 VGND.n2887 VGND.t2556 8.51132
R19665 VGND.n2888 VGND.t3030 8.51132
R19666 VGND.n2888 VGND.t2880 8.51132
R19667 VGND.n2889 VGND.t4399 8.51132
R19668 VGND.n2889 VGND.t374 8.51132
R19669 VGND.n2890 VGND.t5518 8.51132
R19670 VGND.n2890 VGND.t2352 8.51132
R19671 VGND.n2893 VGND.t1209 8.51132
R19672 VGND.n2895 VGND.t4706 8.51132
R19673 VGND.n2897 VGND.t4575 8.51132
R19674 VGND.n2899 VGND.t2299 8.51132
R19675 VGND.n2901 VGND.t5349 8.51132
R19676 VGND.n2903 VGND.t2397 8.51132
R19677 VGND.n2905 VGND.t60 8.51132
R19678 VGND.n2907 VGND.t522 8.51132
R19679 VGND.n2910 VGND.t2888 8.51132
R19680 VGND.n2910 VGND.t3847 8.51132
R19681 VGND.n2912 VGND.t5136 8.51132
R19682 VGND.n2913 VGND.t3906 8.51132
R19683 VGND.n2914 VGND.t3557 8.51132
R19684 VGND.n2915 VGND.t689 8.51132
R19685 VGND.n2917 VGND.t439 8.51132
R19686 VGND.n2918 VGND.t4912 8.51132
R19687 VGND.n2919 VGND.t3498 8.51132
R19688 VGND.n2949 VGND.t2509 8.51132
R19689 VGND.n2948 VGND.t1336 8.51132
R19690 VGND.n2947 VGND.t4888 8.51132
R19691 VGND.n2946 VGND.t2706 8.51132
R19692 VGND.n2945 VGND.t812 8.51132
R19693 VGND.n2944 VGND.t1229 8.51132
R19694 VGND.n2943 VGND.t5208 8.51132
R19695 VGND.n2942 VGND.t5006 8.51132
R19696 VGND.n2940 VGND.t4755 8.51132
R19697 VGND.n2939 VGND.t308 8.51132
R19698 VGND.n2938 VGND.t4236 8.51132
R19699 VGND.n2937 VGND.t4775 8.51132
R19700 VGND.n2936 VGND.t2710 8.51132
R19701 VGND.n2934 VGND.t1469 8.51132
R19702 VGND.n2933 VGND.t3563 8.51132
R19703 VGND.n2932 VGND.t4950 8.51132
R19704 VGND.n2930 VGND.t3449 8.51132
R19705 VGND.n2929 VGND.t3286 8.51132
R19706 VGND.n2928 VGND.t1876 8.51132
R19707 VGND.n2927 VGND.t3805 8.51132
R19708 VGND.n2926 VGND.t1882 8.51132
R19709 VGND.n2925 VGND.t6818 8.51132
R19710 VGND.n2924 VGND.t1500 8.51132
R19711 VGND.n2923 VGND.t2028 8.51132
R19712 VGND.n2909 VGND.t3069 8.51132
R19713 VGND.n2906 VGND.t2336 8.51132
R19714 VGND.n2904 VGND.t2613 8.51132
R19715 VGND.n2902 VGND.t5168 8.51132
R19716 VGND.n2900 VGND.t1541 8.51132
R19717 VGND.n2898 VGND.t3876 8.51132
R19718 VGND.n2896 VGND.t4558 8.51132
R19719 VGND.n2894 VGND.t3464 8.51132
R19720 VGND.n2892 VGND.t4818 8.51132
R19721 VGND.n2503 VGND.t3783 8.51132
R19722 VGND.n2513 VGND.t2039 8.51132
R19723 VGND.n2516 VGND.t3863 8.51132
R19724 VGND.n2523 VGND.t5082 8.51132
R19725 VGND.n2526 VGND.t1519 8.51132
R19726 VGND.n2528 VGND.t3641 8.51132
R19727 VGND.n2531 VGND.t3454 8.51132
R19728 VGND.n2534 VGND.t2109 8.51132
R19729 VGND.n2537 VGND.t4394 8.51132
R19730 VGND.n2539 VGND.t1913 8.51132
R19731 VGND.n2541 VGND.t5752 8.51132
R19732 VGND.n2543 VGND.t5432 8.51132
R19733 VGND.n2545 VGND.t2212 8.51132
R19734 VGND.n2547 VGND.t2391 8.51132
R19735 VGND.n2549 VGND.t4148 8.51132
R19736 VGND.n2551 VGND.t5559 8.51132
R19737 VGND.n2968 VGND.t5754 8.51132
R19738 VGND.n2966 VGND.t6090 8.51132
R19739 VGND.n2964 VGND.t685 8.51132
R19740 VGND.n2997 VGND.t5204 8.51132
R19741 VGND.n2995 VGND.t822 8.51132
R19742 VGND.n2993 VGND.t846 8.51132
R19743 VGND.n2990 VGND.t5188 8.51132
R19744 VGND.n2990 VGND.t565 8.51132
R19745 VGND.n2989 VGND.t1054 8.51132
R19746 VGND.n2989 VGND.t4878 8.51132
R19747 VGND.n2988 VGND.t981 8.51132
R19748 VGND.n2988 VGND.t5735 8.51132
R19749 VGND.n2987 VGND.t1205 8.51132
R19750 VGND.n2987 VGND.t2834 8.51132
R19751 VGND.n2985 VGND.t4046 8.51132
R19752 VGND.n2983 VGND.t2533 8.51132
R19753 VGND.n2981 VGND.t58 8.51132
R19754 VGND.n2979 VGND.t3235 8.51132
R19755 VGND.n2976 VGND.t1999 8.51132
R19756 VGND.n2976 VGND.t957 8.51132
R19757 VGND.n2975 VGND.t1686 8.51132
R19758 VGND.n2975 VGND.t4808 8.51132
R19759 VGND.n2974 VGND.t806 8.51132
R19760 VGND.n2974 VGND.t6800 8.51132
R19761 VGND.n2973 VGND.t4328 8.51132
R19762 VGND.n2973 VGND.t4468 8.51132
R19763 VGND.n2972 VGND.t1025 8.51132
R19764 VGND.n2972 VGND.t5634 8.51132
R19765 VGND.n3044 VGND.t752 8.51132
R19766 VGND.n3044 VGND.t1362 8.51132
R19767 VGND.n3045 VGND.t445 8.51132
R19768 VGND.n3045 VGND.t624 8.51132
R19769 VGND.n3046 VGND.t894 8.51132
R19770 VGND.n3046 VGND.t849 8.51132
R19771 VGND.n3049 VGND.t4208 8.51132
R19772 VGND.n3051 VGND.t1233 8.51132
R19773 VGND.n3053 VGND.t1168 8.51132
R19774 VGND.n3055 VGND.t4299 8.51132
R19775 VGND.n3058 VGND.t2794 8.51132
R19776 VGND.n3059 VGND.t2754 8.51132
R19777 VGND.n3059 VGND.t5041 8.51132
R19778 VGND.n3060 VGND.t5287 8.51132
R19779 VGND.n3060 VGND.t441 8.51132
R19780 VGND.n3061 VGND.t3459 8.51132
R19781 VGND.n3061 VGND.t5009 8.51132
R19782 VGND.n3071 VGND.t4500 8.51132
R19783 VGND.n3069 VGND.t3599 8.51132
R19784 VGND.n3067 VGND.t5671 8.51132
R19785 VGND.n3065 VGND.t2562 8.51132
R19786 VGND.n3063 VGND.t5406 8.51132
R19787 VGND.n375 VGND.t2802 8.51132
R19788 VGND.n3101 VGND.t2615 8.51132
R19789 VGND.n3099 VGND.t6056 8.51132
R19790 VGND.n3096 VGND.t3322 8.51132
R19791 VGND.n3096 VGND.t5766 8.51132
R19792 VGND.n3095 VGND.t3815 8.51132
R19793 VGND.n3095 VGND.t1868 8.51132
R19794 VGND.n3094 VGND.t1801 8.51132
R19795 VGND.n3094 VGND.t1355 8.51132
R19796 VGND.n3093 VGND.t2093 8.51132
R19797 VGND.n3093 VGND.t4125 8.51132
R19798 VGND.n3092 VGND.t2970 8.51132
R19799 VGND.n3092 VGND.t3174 8.51132
R19800 VGND.n3090 VGND.t1135 8.51132
R19801 VGND.n3088 VGND.t5629 8.51132
R19802 VGND.n3086 VGND.t482 8.51132
R19803 VGND.n3083 VGND.t4707 8.51132
R19804 VGND.n3083 VGND.t639 8.51132
R19805 VGND.n3082 VGND.t5652 8.51132
R19806 VGND.n3082 VGND.t5430 8.51132
R19807 VGND.n3081 VGND.t4783 8.51132
R19808 VGND.n3081 VGND.t3518 8.51132
R19809 VGND.n3080 VGND.t3264 8.51132
R19810 VGND.n3080 VGND.t924 8.51132
R19811 VGND.n3079 VGND.t1177 8.51132
R19812 VGND.n3079 VGND.t2974 8.51132
R19813 VGND.n3078 VGND.t2288 8.51132
R19814 VGND.n3078 VGND.t810 8.51132
R19815 VGND.n3148 VGND.t1972 8.51132
R19816 VGND.n3148 VGND.t5378 8.51132
R19817 VGND.n3149 VGND.t5134 8.51132
R19818 VGND.n3149 VGND.t4640 8.51132
R19819 VGND.n3152 VGND.t310 8.51132
R19820 VGND.n3154 VGND.t844 8.51132
R19821 VGND.n3156 VGND.t3817 8.51132
R19822 VGND.n3158 VGND.t6082 8.51132
R19823 VGND.n3160 VGND.t2669 8.51132
R19824 VGND.n3163 VGND.t3403 8.51132
R19825 VGND.n3164 VGND.t2002 8.51132
R19826 VGND.n3164 VGND.t1086 8.51132
R19827 VGND.n3165 VGND.t5361 8.51132
R19828 VGND.n3165 VGND.t3162 8.51132
R19829 VGND.n3177 VGND.t1984 8.51132
R19830 VGND.n3175 VGND.t2663 8.51132
R19831 VGND.n3173 VGND.t816 8.51132
R19832 VGND.n3171 VGND.t3873 8.51132
R19833 VGND.n3169 VGND.t4746 8.51132
R19834 VGND.n3167 VGND.t715 8.51132
R19835 VGND.n3207 VGND.t2001 8.51132
R19836 VGND.n3205 VGND.t6177 8.51132
R19837 VGND.n3202 VGND.t4132 8.51132
R19838 VGND.n3202 VGND.t4662 8.51132
R19839 VGND.n3201 VGND.t893 8.51132
R19840 VGND.n3201 VGND.t2676 8.51132
R19841 VGND.n3200 VGND.t667 8.51132
R19842 VGND.n3200 VGND.t3660 8.51132
R19843 VGND.n3199 VGND.t4136 8.51132
R19844 VGND.n3199 VGND.t736 8.51132
R19845 VGND.n3198 VGND.t1625 8.51132
R19846 VGND.n3198 VGND.t3902 8.51132
R19847 VGND.n3197 VGND.t574 8.51132
R19848 VGND.n3197 VGND.t368 8.51132
R19849 VGND.n3195 VGND.t3338 8.51132
R19850 VGND.n3193 VGND.t4390 8.51132
R19851 VGND.n3190 VGND.t3296 8.51132
R19852 VGND.n3190 VGND.t2230 8.51132
R19853 VGND.n3189 VGND.t3716 8.51132
R19854 VGND.n3189 VGND.t3178 8.51132
R19855 VGND.n3188 VGND.t4105 8.51132
R19856 VGND.n3188 VGND.t2162 8.51132
R19857 VGND.n3187 VGND.t3223 8.51132
R19858 VGND.n3187 VGND.t3127 8.51132
R19859 VGND.n3186 VGND.t4603 8.51132
R19860 VGND.n3186 VGND.t596 8.51132
R19861 VGND.n3185 VGND.t3053 8.51132
R19862 VGND.n3185 VGND.t4177 8.51132
R19863 VGND.n3184 VGND.t3948 8.51132
R19864 VGND.n3184 VGND.t5580 8.51132
R19865 VGND.n3276 VGND.t1978 8.51132
R19866 VGND.n3276 VGND.t2049 8.51132
R19867 VGND.n3279 VGND.t4803 8.51132
R19868 VGND.n3281 VGND.t5963 8.51132
R19869 VGND.n3283 VGND.t2552 8.51132
R19870 VGND.n3285 VGND.t3620 8.51132
R19871 VGND.n3287 VGND.t6062 8.51132
R19872 VGND.n3289 VGND.t2444 8.51132
R19873 VGND.n3292 VGND.t3293 8.51132
R19874 VGND.n3293 VGND.t4126 8.51132
R19875 VGND.n3293 VGND.t3229 8.51132
R19876 VGND.n3307 VGND.t3533 8.51132
R19877 VGND.n3305 VGND.t1817 8.51132
R19878 VGND.n3303 VGND.t5267 8.51132
R19879 VGND.n3301 VGND.t3141 8.51132
R19880 VGND.n3299 VGND.t3725 8.51132
R19881 VGND.n3297 VGND.t6773 8.51132
R19882 VGND.n3295 VGND.t2831 8.51132
R19883 VGND.n3334 VGND.t3553 8.51132
R19884 VGND.n3331 VGND.t1944 8.51132
R19885 VGND.n3331 VGND.t5709 8.51132
R19886 VGND.n3330 VGND.t3164 8.51132
R19887 VGND.n3330 VGND.t3986 8.51132
R19888 VGND.n3329 VGND.t1121 8.51132
R19889 VGND.n3329 VGND.t5100 8.51132
R19890 VGND.n3328 VGND.t1129 8.51132
R19891 VGND.n3328 VGND.t5212 8.51132
R19892 VGND.n3327 VGND.t2494 8.51132
R19893 VGND.n3327 VGND.t6005 8.51132
R19894 VGND.n3326 VGND.t5375 8.51132
R19895 VGND.n3326 VGND.t1137 8.51132
R19896 VGND.n3325 VGND.t1092 8.51132
R19897 VGND.n3325 VGND.t68 8.51132
R19898 VGND.n3323 VGND.t5455 8.51132
R19899 VGND.n3320 VGND.t1548 8.51132
R19900 VGND.n3320 VGND.t1273 8.51132
R19901 VGND.n3319 VGND.t3298 8.51132
R19902 VGND.n3319 VGND.t3787 8.51132
R19903 VGND.n3318 VGND.t1888 8.51132
R19904 VGND.n3318 VGND.t6774 8.51132
R19905 VGND.n3317 VGND.t1207 8.51132
R19906 VGND.n3317 VGND.t2835 8.51132
R19907 VGND.n3316 VGND.t378 8.51132
R19908 VGND.n3316 VGND.t559 8.51132
R19909 VGND.n3315 VGND.t514 8.51132
R19910 VGND.n3315 VGND.t6168 8.51132
R19911 VGND.n3314 VGND.t1482 8.51132
R19912 VGND.n3314 VGND.t896 8.51132
R19913 VGND.n4 VGND.t550 8.51132
R19914 VGND.n4 VGND.t2302 8.51132
R19915 VGND.n3751 VGND.t934 8.51132
R19916 VGND.n3749 VGND.t1731 8.51132
R19917 VGND.n3747 VGND.t4173 8.51132
R19918 VGND.n3745 VGND.t2852 8.51132
R19919 VGND.n3743 VGND.t841 8.51132
R19920 VGND.n3741 VGND.t1159 8.51132
R19921 VGND.n3739 VGND.t4624 8.51132
R19922 VGND.n3736 VGND.t1046 8.51132
R19923 VGND.n3733 VGND.t5312 8.51132
R19924 VGND.n3731 VGND.t5923 8.51132
R19925 VGND.n3729 VGND.t2497 8.51132
R19926 VGND.n3727 VGND.t4577 8.51132
R19927 VGND.n3725 VGND.t5638 8.51132
R19928 VGND.n3723 VGND.t5854 8.51132
R19929 VGND.n3721 VGND.t632 8.51132
R19930 VGND.n3719 VGND.t3196 8.51132
R19931 VGND.n16 VGND.t5587 8.51132
R19932 VGND.n16 VGND.t4130 8.51132
R19933 VGND.n15 VGND.t5768 8.51132
R19934 VGND.n15 VGND.t2953 8.51132
R19935 VGND.n14 VGND.t4734 8.51132
R19936 VGND.n14 VGND.t1172 8.51132
R19937 VGND.n13 VGND.t3564 8.51132
R19938 VGND.n13 VGND.t1221 8.51132
R19939 VGND.n12 VGND.t348 8.51132
R19940 VGND.n12 VGND.t2769 8.51132
R19941 VGND.n11 VGND.t1225 8.51132
R19942 VGND.n11 VGND.t4702 8.51132
R19943 VGND.n10 VGND.t1293 8.51132
R19944 VGND.n10 VGND.t5933 8.51132
R19945 VGND.n9 VGND.t2968 8.51132
R19946 VGND.n9 VGND.t2923 8.51132
R19947 VGND.n17 VGND.t5762 8.51132
R19948 VGND.n3720 VGND.t4924 8.51132
R19949 VGND.n3722 VGND.t3545 8.51132
R19950 VGND.n3724 VGND.t2649 8.51132
R19951 VGND.n3726 VGND.t4244 8.51132
R19952 VGND.n3728 VGND.t423 8.51132
R19953 VGND.n3730 VGND.t798 8.51132
R19954 VGND.n3732 VGND.t4355 8.51132
R19955 VGND.n3734 VGND.t657 8.51132
R19956 VGND.n3738 VGND.t1729 8.51132
R19957 VGND.n3740 VGND.t4182 8.51132
R19958 VGND.n3742 VGND.t4773 8.51132
R19959 VGND.n3744 VGND.t3365 8.51132
R19960 VGND.n3746 VGND.t4210 8.51132
R19961 VGND.n3748 VGND.t1475 8.51132
R19962 VGND.n3750 VGND.t5071 8.51132
R19963 VGND.n3752 VGND.t4592 8.51132
R19964 VGND.n3321 VGND.t830 8.51132
R19965 VGND.n3332 VGND.t520 8.51132
R19966 VGND.n3294 VGND.t3083 8.51132
R19967 VGND.n3296 VGND.t6007 8.51132
R19968 VGND.n3298 VGND.t4060 8.51132
R19969 VGND.n3300 VGND.t4948 8.51132
R19970 VGND.n3302 VGND.t1616 8.51132
R19971 VGND.n3304 VGND.t5274 8.51132
R19972 VGND.n3306 VGND.t3811 8.51132
R19973 VGND.n3308 VGND.t5775 8.51132
R19974 VGND.n3290 VGND.t1713 8.51132
R19975 VGND.n3288 VGND.t1227 8.51132
R19976 VGND.n3286 VGND.t5727 8.51132
R19977 VGND.n3284 VGND.t6054 8.51132
R19978 VGND.n3282 VGND.t5539 8.51132
R19979 VGND.n3280 VGND.t5832 8.51132
R19980 VGND.n3278 VGND.t1780 8.51132
R19981 VGND.n3191 VGND.t1994 8.51132
R19982 VGND.n3194 VGND.t1119 8.51132
R19983 VGND.n3203 VGND.t748 8.51132
R19984 VGND.n3206 VGND.t5073 8.51132
R19985 VGND.n3166 VGND.t4599 8.51132
R19986 VGND.n3168 VGND.t1721 8.51132
R19987 VGND.n3170 VGND.t1488 8.51132
R19988 VGND.n3172 VGND.t4620 8.51132
R19989 VGND.n3174 VGND.t384 8.51132
R19990 VGND.n3176 VGND.t634 8.51132
R19991 VGND.n3178 VGND.t1891 8.51132
R19992 VGND.n3161 VGND.t2845 8.51132
R19993 VGND.n3159 VGND.t1052 8.51132
R19994 VGND.n3157 VGND.t1897 8.51132
R19995 VGND.n3155 VGND.t4853 8.51132
R19996 VGND.n3153 VGND.t2164 8.51132
R19997 VGND.n3151 VGND.t1753 8.51132
R19998 VGND.n3084 VGND.t2579 8.51132
R19999 VGND.n3087 VGND.t4626 8.51132
R20000 VGND.n3089 VGND.t3089 8.51132
R20001 VGND.n3097 VGND.t1646 8.51132
R20002 VGND.n3100 VGND.t4485 8.51132
R20003 VGND.n3102 VGND.t3865 8.51132
R20004 VGND.n3062 VGND.t3735 8.51132
R20005 VGND.n3064 VGND.t4762 8.51132
R20006 VGND.n3066 VGND.t3007 8.51132
R20007 VGND.n3068 VGND.t4635 8.51132
R20008 VGND.n3070 VGND.t1954 8.51132
R20009 VGND.n3072 VGND.t1691 8.51132
R20010 VGND.n3056 VGND.t532 8.51132
R20011 VGND.n3054 VGND.t4805 8.51132
R20012 VGND.n3052 VGND.t3759 8.51132
R20013 VGND.n3050 VGND.t4286 8.51132
R20014 VGND.n3048 VGND.t4466 8.51132
R20015 VGND.n2977 VGND.t4633 8.51132
R20016 VGND.n2980 VGND.t3506 8.51132
R20017 VGND.n2982 VGND.t754 8.51132
R20018 VGND.n2984 VGND.t839 8.51132
R20019 VGND.n2991 VGND.t1110 8.51132
R20020 VGND.n2994 VGND.t4801 8.51132
R20021 VGND.n2996 VGND.t366 8.51132
R20022 VGND.n2963 VGND.t818 8.51132
R20023 VGND.n2965 VGND.t2999 8.51132
R20024 VGND.n2967 VGND.t2073 8.51132
R20025 VGND.n381 VGND.t4342 8.51132
R20026 VGND.n382 VGND.t2013 8.51132
R20027 VGND.n383 VGND.t2673 8.51132
R20028 VGND.n3002 VGND.t700 8.51132
R20029 VGND.n3003 VGND.t4406 8.51132
R20030 VGND.n3004 VGND.t5552 8.51132
R20031 VGND.n3006 VGND.t5859 8.51132
R20032 VGND.n3007 VGND.t3951 8.51132
R20033 VGND.n3008 VGND.t1275 8.51132
R20034 VGND.n3009 VGND.t4799 8.51132
R20035 VGND.n3010 VGND.t4617 8.51132
R20036 VGND.n3011 VGND.t4021 8.51132
R20037 VGND.n3012 VGND.t1962 8.51132
R20038 VGND.n3013 VGND.t2932 8.51132
R20039 VGND.n3017 VGND.t5764 8.51132
R20040 VGND.n3016 VGND.t2442 8.51132
R20041 VGND.n3015 VGND.t4926 8.51132
R20042 VGND.n3014 VGND.t2425 8.51132
R20043 VGND.n379 VGND.t1960 8.51132
R20044 VGND.n3039 VGND.t5310 8.51132
R20045 VGND.n3038 VGND.t5043 8.51132
R20046 VGND.n3037 VGND.t1164 8.51132
R20047 VGND.n3035 VGND.t1303 8.51132
R20048 VGND.n3034 VGND.t4768 8.51132
R20049 VGND.n3033 VGND.t4013 8.51132
R20050 VGND.n3032 VGND.t3953 8.51132
R20051 VGND.n3031 VGND.t2034 8.51132
R20052 VGND.n3030 VGND.t2549 8.51132
R20053 VGND.n3029 VGND.t2804 8.51132
R20054 VGND.n3028 VGND.t2809 8.51132
R20055 VGND.n3026 VGND.t5943 8.51132
R20056 VGND.n3025 VGND.t4585 8.51132
R20057 VGND.n3024 VGND.t1259 8.51132
R20058 VGND.n3023 VGND.t5834 8.51132
R20059 VGND.n3022 VGND.t2484 8.51132
R20060 VGND.n373 VGND.t3733 8.51132
R20061 VGND.n3107 VGND.t5642 8.51132
R20062 VGND.n3108 VGND.t4259 8.51132
R20063 VGND.n3110 VGND.t4594 8.51132
R20064 VGND.n3111 VGND.t2777 8.51132
R20065 VGND.n3112 VGND.t3160 8.51132
R20066 VGND.n3113 VGND.t2667 8.51132
R20067 VGND.n3114 VGND.t5547 8.51132
R20068 VGND.n3115 VGND.t628 8.51132
R20069 VGND.n3116 VGND.t4240 8.51132
R20070 VGND.n3117 VGND.t1968 8.51132
R20071 VGND.n3122 VGND.t2129 8.51132
R20072 VGND.n3121 VGND.t6754 8.51132
R20073 VGND.n3120 VGND.t6086 8.51132
R20074 VGND.n3119 VGND.t904 8.51132
R20075 VGND.n3118 VGND.t4986 8.51132
R20076 VGND.n371 VGND.t4401 8.51132
R20077 VGND.n3143 VGND.t2531 8.51132
R20078 VGND.n3142 VGND.t4000 8.51132
R20079 VGND.n3140 VGND.t2139 8.51132
R20080 VGND.n3139 VGND.t4583 8.51132
R20081 VGND.n3138 VGND.t407 8.51132
R20082 VGND.n3137 VGND.t1552 8.51132
R20083 VGND.n3136 VGND.t3367 8.51132
R20084 VGND.n3135 VGND.t4748 8.51132
R20085 VGND.n3134 VGND.t4388 8.51132
R20086 VGND.n3133 VGND.t626 8.51132
R20087 VGND.n3131 VGND.t3180 8.51132
R20088 VGND.n3130 VGND.t4664 8.51132
R20089 VGND.n3129 VGND.t5259 8.51132
R20090 VGND.n3128 VGND.t837 8.51132
R20091 VGND.n3127 VGND.t3208 8.51132
R20092 VGND.n366 VGND.t616 8.51132
R20093 VGND.n3212 VGND.t4631 8.51132
R20094 VGND.n3213 VGND.t2041 8.51132
R20095 VGND.n3215 VGND.t2207 8.51132
R20096 VGND.n3216 VGND.t3284 8.51132
R20097 VGND.n3217 VGND.t1719 8.51132
R20098 VGND.n3218 VGND.t5484 8.51132
R20099 VGND.n3219 VGND.t3087 8.51132
R20100 VGND.n3220 VGND.t4709 8.51132
R20101 VGND.n3221 VGND.t3791 8.51132
R20102 VGND.n3222 VGND.t3111 8.51132
R20103 VGND.n3228 VGND.t3766 8.51132
R20104 VGND.n3227 VGND.t1621 8.51132
R20105 VGND.n3226 VGND.t1735 8.51132
R20106 VGND.n3225 VGND.t2554 8.51132
R20107 VGND.n3224 VGND.t4099 8.51132
R20108 VGND.n3223 VGND.t5529 8.51132
R20109 VGND.n364 VGND.t2976 8.51132
R20110 VGND.n3271 VGND.t3350 8.51132
R20111 VGND.n3269 VGND.t1936 8.51132
R20112 VGND.n3268 VGND.t6162 8.51132
R20113 VGND.n3267 VGND.t6814 8.51132
R20114 VGND.n3266 VGND.t5989 8.51132
R20115 VGND.n3265 VGND.t5497 8.51132
R20116 VGND.n3264 VGND.t1584 8.51132
R20117 VGND.n3263 VGND.t6030 8.51132
R20118 VGND.n3262 VGND.t2833 8.51132
R20119 VGND.n3260 VGND.t936 8.51132
R20120 VGND.n3259 VGND.t357 8.51132
R20121 VGND.n3258 VGND.t3401 8.51132
R20122 VGND.n3257 VGND.t5488 8.51132
R20123 VGND.n3256 VGND.t5291 8.51132
R20124 VGND.n3255 VGND.t5965 8.51132
R20125 VGND.n3254 VGND.t411 8.51132
R20126 VGND.n3252 VGND.t5190 8.51132
R20127 VGND.n3250 VGND.t4778 8.51132
R20128 VGND.n3249 VGND.t4668 8.51132
R20129 VGND.n3248 VGND.t4145 8.51132
R20130 VGND.n3247 VGND.t6761 8.51132
R20131 VGND.n3246 VGND.t2837 8.51132
R20132 VGND.n3245 VGND.t932 8.51132
R20133 VGND.n3244 VGND.t3466 8.51132
R20134 VGND.n3243 VGND.t5520 8.51132
R20135 VGND.n3241 VGND.t4791 8.51132
R20136 VGND.n3240 VGND.t3693 8.51132
R20137 VGND.n3239 VGND.t1419 8.51132
R20138 VGND.n3238 VGND.t4437 8.51132
R20139 VGND.n3237 VGND.t2854 8.51132
R20140 VGND.n3236 VGND.t5490 8.51132
R20141 VGND.n3235 VGND.t2748 8.51132
R20142 VGND.n2 VGND.t5967 8.51132
R20143 VGND.n3759 VGND.t4410 8.51132
R20144 VGND.n3760 VGND.t5864 8.51132
R20145 VGND.n3761 VGND.t3318 8.51132
R20146 VGND.n3762 VGND.t4628 8.51132
R20147 VGND.n3763 VGND.t4579 8.51132
R20148 VGND.n3764 VGND.t443 8.51132
R20149 VGND.n3765 VGND.t2547 8.51132
R20150 VGND.n3766 VGND.t5341 8.51132
R20151 VGND.n3774 VGND.t5945 8.51132
R20152 VGND.n3773 VGND.t5618 8.51132
R20153 VGND.n3772 VGND.t3373 8.51132
R20154 VGND.n3771 VGND.t338 8.51132
R20155 VGND.n3770 VGND.t5935 8.51132
R20156 VGND.n3769 VGND.t2115 8.51132
R20157 VGND.n3768 VGND.t1328 8.51132
R20158 VGND.n3767 VGND.t2203 8.51132
R20159 VGND.n3785 VGND.t4085 8.51132
R20160 VGND.n3784 VGND.t1301 8.51132
R20161 VGND.n3783 VGND.t2174 8.51132
R20162 VGND.n3782 VGND.t70 8.51132
R20163 VGND.n3781 VGND.t636 8.51132
R20164 VGND.n3780 VGND.t4573 8.51132
R20165 VGND.n3779 VGND.t3488 8.51132
R20166 VGND.n3778 VGND.t1443 8.51132
R20167 VGND.n628 VGND.t3631 8.49619
R20168 VGND.n1926 VGND.t5090 8.49619
R20169 VGND.n856 VGND.t4456 8.49371
R20170 VGND.n852 VGND.t4453 8.49371
R20171 VGND.n1325 VGND.t2517 8.49371
R20172 VGND.n1329 VGND.t2525 8.49371
R20173 VGND.n1330 VGND.t6017 8.49371
R20174 VGND.n1334 VGND.t6015 8.49371
R20175 VGND.n1335 VGND.t5047 8.49371
R20176 VGND.n1331 VGND.t5051 8.49371
R20177 VGND.n1613 VGND.t1349 8.49371
R20178 VGND.n1609 VGND.t1353 8.49371
R20179 VGND.n2077 VGND.t6154 8.48197
R20180 VGND.n754 VGND.t4672 8.48197
R20181 VGND.n1921 VGND.t6576 8.48197
R20182 VGND.n177 VGND.t5211 8.47806
R20183 VGND.n179 VGND.t2456 8.47806
R20184 VGND.n188 VGND.t2199 8.47806
R20185 VGND.n183 VGND.t2044 8.47806
R20186 VGND.n231 VGND.t2463 8.47806
R20187 VGND.n65 VGND.t5129 8.47806
R20188 VGND.n71 VGND.t5651 8.47806
R20189 VGND.n78 VGND.t3969 8.47806
R20190 VGND.n84 VGND.t1305 8.47219
R20191 VGND.n90 VGND.t322 8.47219
R20192 VGND.n94 VGND.t1150 8.47219
R20193 VGND.n104 VGND.t2181 8.47219
R20194 VGND.n1337 VGND.t4886 8.47219
R20195 VGND.n1019 VGND.t6046 8.47023
R20196 VGND.n1017 VGND.t6048 8.47023
R20197 VGND.n1015 VGND.t1427 8.47023
R20198 VGND.n1064 VGND.t1429 8.47023
R20199 VGND.n1062 VGND.t739 8.47023
R20200 VGND.n1060 VGND.t741 8.47023
R20201 VGND.n1056 VGND.t4458 8.47023
R20202 VGND.n1053 VGND.t4460 8.47023
R20203 VGND.n1052 VGND.t512 8.47023
R20204 VGND.n1049 VGND.t510 8.47023
R20205 VGND.n1048 VGND.t5028 8.47023
R20206 VGND.n1046 VGND.t5030 8.47023
R20207 VGND.n1044 VGND.t4347 8.47023
R20208 VGND.n1042 VGND.t4349 8.47023
R20209 VGND.n1041 VGND.t2732 8.47023
R20210 VGND.n1039 VGND.t2734 8.47023
R20211 VGND.n1038 VGND.t1652 8.47023
R20212 VGND.n1036 VGND.t1650 8.47023
R20213 VGND.n1033 VGND.t722 8.47023
R20214 VGND.n1031 VGND.t724 8.47023
R20215 VGND.n1029 VGND.t3836 8.47023
R20216 VGND.n1027 VGND.t3834 8.47023
R20217 VGND.n1025 VGND.t3190 8.47023
R20218 VGND.n574 VGND.t3192 8.47023
R20219 VGND.n2008 VGND.t1632 8.47023
R20220 VGND.n2010 VGND.t1630 8.47023
R20221 VGND.n2015 VGND.t3280 8.47023
R20222 VGND.n2017 VGND.t3282 8.47023
R20223 VGND.n2018 VGND.t5013 8.47023
R20224 VGND.n2021 VGND.t5015 8.47023
R20225 VGND.n2022 VGND.t3276 8.47023
R20226 VGND.n2020 VGND.t3278 8.47023
R20227 VGND.n2016 VGND.t2724 8.47023
R20228 VGND.n2014 VGND.t2722 8.47023
R20229 VGND.n2013 VGND.t2728 8.47023
R20230 VGND.n2011 VGND.t2726 8.47023
R20231 VGND.n2005 VGND.t2378 8.47023
R20232 VGND.n1024 VGND.t2376 8.47023
R20233 VGND.n1026 VGND.t5610 8.47023
R20234 VGND.n1028 VGND.t5608 8.47023
R20235 VGND.n1032 VGND.t2997 8.47023
R20236 VGND.n1034 VGND.t2995 8.47023
R20237 VGND.n1043 VGND.t1682 8.47023
R20238 VGND.n1045 VGND.t1684 8.47023
R20239 VGND.n1051 VGND.t2965 8.47023
R20240 VGND.n1054 VGND.t2963 8.47023
R20241 VGND.n1055 VGND.t316 8.47023
R20242 VGND.n1057 VGND.t314 8.47023
R20243 VGND.n1059 VGND.t3314 8.47023
R20244 VGND.n1061 VGND.t3316 8.47023
R20245 VGND.n932 VGND.t1662 8.47023
R20246 VGND.n930 VGND.t1661 8.47023
R20247 VGND.n813 VGND.t2358 8.47023
R20248 VGND.n812 VGND.t2357 8.47023
R20249 VGND.n810 VGND.t5710 8.47023
R20250 VGND.n809 VGND.t5711 8.47023
R20251 VGND.n920 VGND.t4724 8.47023
R20252 VGND.n922 VGND.t4723 8.47023
R20253 VGND.n934 VGND.t2446 8.47023
R20254 VGND.n917 VGND.t2445 8.47023
R20255 VGND.n915 VGND.t5515 8.47023
R20256 VGND.n914 VGND.t5514 8.47023
R20257 VGND.n913 VGND.t1459 8.47023
R20258 VGND.n911 VGND.t1458 8.47023
R20259 VGND.n900 VGND.t1463 8.47023
R20260 VGND.n902 VGND.t1461 8.47023
R20261 VGND.n904 VGND.t1144 8.47023
R20262 VGND.n906 VGND.t1146 8.47023
R20263 VGND.n908 VGND.t1664 8.47023
R20264 VGND.n1283 VGND.t1666 8.47023
R20265 VGND.n1285 VGND.t5462 8.47023
R20266 VGND.n1287 VGND.t5464 8.47023
R20267 VGND.n1291 VGND.t3643 8.47023
R20268 VGND.n1294 VGND.t3645 8.47023
R20269 VGND.n1319 VGND.t2046 8.47023
R20270 VGND.n1322 VGND.t2048 8.47023
R20271 VGND.n1323 VGND.t3356 8.47023
R20272 VGND.n1321 VGND.t3358 8.47023
R20273 VGND.n1320 VGND.t1859 8.47023
R20274 VGND.n1317 VGND.t1861 8.47023
R20275 VGND.n1295 VGND.t2940 8.47023
R20276 VGND.n1293 VGND.t2942 8.47023
R20277 VGND.n1292 VGND.t4719 8.47023
R20278 VGND.n1290 VGND.t4721 8.47023
R20279 VGND.n1288 VGND.t4224 8.47023
R20280 VGND.n1286 VGND.t4222 8.47023
R20281 VGND.n1284 VGND.t3568 8.47023
R20282 VGND.n1282 VGND.t3566 8.47023
R20283 VGND.n907 VGND.t2781 8.47023
R20284 VGND.n905 VGND.t2779 8.47023
R20285 VGND.n903 VGND.t3131 8.47023
R20286 VGND.n901 VGND.t3129 8.47023
R20287 VGND.n1244 VGND.t2745 8.47023
R20288 VGND.n1244 VGND.t1848 8.47023
R20289 VGND.n1243 VGND.t2746 8.47023
R20290 VGND.n1243 VGND.t1850 8.47023
R20291 VGND.n1242 VGND.t2083 8.47023
R20292 VGND.n1242 VGND.t2167 8.47023
R20293 VGND.n1241 VGND.t2085 8.47023
R20294 VGND.n1241 VGND.t2168 8.47023
R20295 VGND.n1240 VGND.t2170 8.47023
R20296 VGND.n1240 VGND.t5516 8.47023
R20297 VGND.n1277 VGND.t2172 8.47023
R20298 VGND.n1277 VGND.t5517 8.47023
R20299 VGND.n1272 VGND.t900 8.47023
R20300 VGND.n1270 VGND.t898 8.47023
R20301 VGND.n1265 VGND.t2991 8.47023
R20302 VGND.n1263 VGND.t2993 8.47023
R20303 VGND.n1622 VGND.t3739 8.47023
R20304 VGND.n1620 VGND.t3741 8.47023
R20305 VGND.n1617 VGND.t2609 8.47023
R20306 VGND.n1619 VGND.t2611 8.47023
R20307 VGND.n1264 VGND.t2119 8.47023
R20308 VGND.n1266 VGND.t2117 8.47023
R20309 VGND.n1268 VGND.t3749 8.47023
R20310 VGND.n1269 VGND.t3747 8.47023
R20311 VGND.n1274 VGND.t2362 8.47023
R20312 VGND.n1276 VGND.t2360 8.47023
R20313 VGND.n1201 VGND.t5422 8.47023
R20314 VGND.n1199 VGND.t5420 8.47023
R20315 VGND.n1197 VGND.t5426 8.47023
R20316 VGND.n1195 VGND.t5424 8.47023
R20317 VGND.n1193 VGND.t1056 8.47023
R20318 VGND.n1237 VGND.t1058 8.47023
R20319 VGND.n1228 VGND.t5228 8.47023
R20320 VGND.n1228 VGND.t5806 8.47023
R20321 VGND.n1227 VGND.t5232 8.47023
R20322 VGND.n1227 VGND.t5807 8.47023
R20323 VGND.n1226 VGND.t1193 8.47023
R20324 VGND.n1226 VGND.t5804 8.47023
R20325 VGND.n1225 VGND.t1195 8.47023
R20326 VGND.n1225 VGND.t5805 8.47023
R20327 VGND.n1224 VGND.t1029 8.47023
R20328 VGND.n1222 VGND.t1027 8.47023
R20329 VGND.n1635 VGND.t4278 8.47023
R20330 VGND.n1637 VGND.t4276 8.47023
R20331 VGND.n1642 VGND.t1010 8.47023
R20332 VGND.n1644 VGND.t4683 8.47023
R20333 VGND.n1646 VGND.t4685 8.47023
R20334 VGND.n1643 VGND.t1012 8.47023
R20335 VGND.n1641 VGND.t4282 8.47023
R20336 VGND.n1638 VGND.t4280 8.47023
R20337 VGND.n1230 VGND.t4118 8.47023
R20338 VGND.n1232 VGND.t4122 8.47023
R20339 VGND.n1234 VGND.t882 8.47023
R20340 VGND.n1235 VGND.t884 8.47023
R20341 VGND.n1236 VGND.t4338 8.47023
R20342 VGND.n1192 VGND.t4336 8.47023
R20343 VGND.n1194 VGND.t4334 8.47023
R20344 VGND.n1196 VGND.t4332 8.47023
R20345 VGND.n1198 VGND.t826 8.47023
R20346 VGND.n1200 VGND.t828 8.47023
R20347 VGND.n1119 VGND.t6785 8.47023
R20348 VGND.n1116 VGND.t6787 8.47023
R20349 VGND.n1114 VGND.t5909 8.47023
R20350 VGND.n1188 VGND.t5911 8.47023
R20351 VGND.n1187 VGND.t1033 8.47023
R20352 VGND.n1185 VGND.t1035 8.47023
R20353 VGND.n1183 VGND.t3437 8.47023
R20354 VGND.n1181 VGND.t3435 8.47023
R20355 VGND.n1179 VGND.t1775 8.47023
R20356 VGND.n1177 VGND.t1773 8.47023
R20357 VGND.n1175 VGND.t2278 8.47023
R20358 VGND.n1173 VGND.t2280 8.47023
R20359 VGND.n1171 VGND.t2274 8.47023
R20360 VGND.n1169 VGND.t2276 8.47023
R20361 VGND.n1168 VGND.t5985 8.47023
R20362 VGND.n1166 VGND.t5983 8.47023
R20363 VGND.n1164 VGND.t1608 8.47023
R20364 VGND.n1161 VGND.t1606 8.47023
R20365 VGND.n1160 VGND.t4005 8.47023
R20366 VGND.n1158 VGND.t4007 8.47023
R20367 VGND.n1156 VGND.t2020 8.47023
R20368 VGND.n1154 VGND.t2022 8.47023
R20369 VGND.n1153 VGND.t2906 8.47023
R20370 VGND.n1152 VGND.t2908 8.47023
R20371 VGND.n1150 VGND.t1244 8.47023
R20372 VGND.n1147 VGND.t1246 8.47023
R20373 VGND.n1146 VGND.t1242 8.47023
R20374 VGND.n1144 VGND.t1240 8.47023
R20375 VGND.n1141 VGND.t1508 8.47023
R20376 VGND.n1139 VGND.t1510 8.47023
R20377 VGND.n1145 VGND.t542 8.47023
R20378 VGND.n1148 VGND.t540 8.47023
R20379 VGND.n1155 VGND.t1604 8.47023
R20380 VGND.n1157 VGND.t1602 8.47023
R20381 VGND.n1159 VGND.t1502 8.47023
R20382 VGND.n1162 VGND.t1504 8.47023
R20383 VGND.n1170 VGND.t1767 8.47023
R20384 VGND.n1172 VGND.t1769 8.47023
R20385 VGND.n1186 VGND.t4362 8.47023
R20386 VGND.n1189 VGND.t4360 8.47023
R20387 VGND.n1115 VGND.t5683 8.47023
R20388 VGND.n1117 VGND.t5685 8.47023
R20389 VGND.n1118 VGND.t5915 8.47023
R20390 VGND.n1121 VGND.t5913 8.47023
R20391 VGND.n1075 VGND.t2399 8.47023
R20392 VGND.n1072 VGND.t2401 8.47023
R20393 VGND.n1071 VGND.t3597 8.47023
R20394 VGND.n1068 VGND.t3595 8.47023
R20395 VGND.n1111 VGND.t5687 8.47023
R20396 VGND.n1108 VGND.t5689 8.47023
R20397 VGND.n1083 VGND.t3823 8.47023
R20398 VGND.n1081 VGND.t3825 8.47023
R20399 VGND.n2000 VGND.t5410 8.47023
R20400 VGND.n2000 VGND.t538 8.47023
R20401 VGND.n1999 VGND.t5409 8.47023
R20402 VGND.n1999 VGND.t536 8.47023
R20403 VGND.n1998 VGND.t5412 8.47023
R20404 VGND.n1996 VGND.t5414 8.47023
R20405 VGND.n1992 VGND.t2476 8.47023
R20406 VGND.n1994 VGND.t2474 8.47023
R20407 VGND.n1995 VGND.t2478 8.47023
R20408 VGND.n1997 VGND.t2480 8.47023
R20409 VGND.n1079 VGND.t5164 8.47023
R20410 VGND.n1080 VGND.t5166 8.47023
R20411 VGND.n1082 VGND.t4566 8.47023
R20412 VGND.n1084 VGND.t4564 8.47023
R20413 VGND.n1088 VGND.t1654 8.47023
R20414 VGND.n1090 VGND.t1656 8.47023
R20415 VGND.n1093 VGND.t508 8.47023
R20416 VGND.n1095 VGND.t506 8.47023
R20417 VGND.n1097 VGND.t5897 8.47023
R20418 VGND.n1099 VGND.t5899 8.47023
R20419 VGND.n1100 VGND.t3990 8.47023
R20420 VGND.n1102 VGND.t3992 8.47023
R20421 VGND.n1103 VGND.t2957 8.47023
R20422 VGND.n1105 VGND.t2959 8.47023
R20423 VGND.n1107 VGND.t1558 8.47023
R20424 VGND.n1109 VGND.t1556 8.47023
R20425 VGND.n1110 VGND.t2692 8.47023
R20426 VGND.n1069 VGND.t2690 8.47023
R20427 VGND.n1070 VGND.t2688 8.47023
R20428 VGND.n1073 VGND.t2686 8.47023
R20429 VGND.n994 VGND.t4918 8.47023
R20430 VGND.n991 VGND.t4920 8.47023
R20431 VGND.n990 VGND.t5571 8.47023
R20432 VGND.n987 VGND.t5573 8.47023
R20433 VGND.n986 VGND.t4691 8.47023
R20434 VGND.n984 VGND.t4693 8.47023
R20435 VGND.n983 VGND.t1421 8.47023
R20436 VGND.n980 VGND.t1423 8.47023
R20437 VGND.n976 VGND.t4958 8.47023
R20438 VGND.n973 VGND.t4960 8.47023
R20439 VGND.n972 VGND.t5301 8.47023
R20440 VGND.n969 VGND.t5303 8.47023
R20441 VGND.n968 VGND.t2915 8.47023
R20442 VGND.n965 VGND.t2913 8.47023
R20443 VGND.n964 VGND.t4257 8.47023
R20444 VGND.n966 VGND.t4255 8.47023
R20445 VGND.n967 VGND.t5495 8.47023
R20446 VGND.n970 VGND.t5493 8.47023
R20447 VGND.n971 VGND.t2917 8.47023
R20448 VGND.n974 VGND.t2919 8.47023
R20449 VGND.n985 VGND.t2252 8.47023
R20450 VGND.n988 VGND.t2254 8.47023
R20451 VGND.n989 VGND.t2862 8.47023
R20452 VGND.n992 VGND.t2860 8.47023
R20453 VGND.n993 VGND.t5661 8.47023
R20454 VGND.n996 VGND.t5663 8.47023
R20455 VGND.n463 VGND.t1311 8.47023
R20456 VGND.n460 VGND.t1313 8.47023
R20457 VGND.n459 VGND.t5871 8.47023
R20458 VGND.n456 VGND.t5873 8.47023
R20459 VGND.n455 VGND.t5994 8.47023
R20460 VGND.n452 VGND.t5992 8.47023
R20461 VGND.n451 VGND.t5665 8.47023
R20462 VGND.n428 VGND.t5667 8.47023
R20463 VGND.n2437 VGND.t606 8.47023
R20464 VGND.n2437 VGND.t5334 8.47023
R20465 VGND.n2436 VGND.t604 8.47023
R20466 VGND.n2436 VGND.t5335 8.47023
R20467 VGND.n2434 VGND.t2016 8.47023
R20468 VGND.n2432 VGND.t2018 8.47023
R20469 VGND.n2429 VGND.t5722 8.47023
R20470 VGND.n2431 VGND.t5720 8.47023
R20471 VGND.n2433 VGND.t1071 8.47023
R20472 VGND.n2435 VGND.t1069 8.47023
R20473 VGND.n450 VGND.t4385 8.47023
R20474 VGND.n453 VGND.t4383 8.47023
R20475 VGND.n454 VGND.t1326 8.47023
R20476 VGND.n457 VGND.t1324 8.47023
R20477 VGND.n458 VGND.t3016 8.47023
R20478 VGND.n461 VGND.t3018 8.47023
R20479 VGND.n2461 VGND.t2101 8.47023
R20480 VGND.n2458 VGND.t2103 8.47023
R20481 VGND.n2457 VGND.t2097 8.47023
R20482 VGND.n2454 VGND.t2099 8.47023
R20483 VGND.n2453 VGND.t1521 8.47023
R20484 VGND.n2450 VGND.t1523 8.47023
R20485 VGND.n2232 VGND.t5149 8.47023
R20486 VGND.n2234 VGND.t5147 8.47023
R20487 VGND.n2236 VGND.t1075 8.47023
R20488 VGND.n2238 VGND.t1073 8.47023
R20489 VGND.n2240 VGND.t5742 8.47023
R20490 VGND.n2241 VGND.t5744 8.47023
R20491 VGND.n2239 VGND.t2783 8.47023
R20492 VGND.n2237 VGND.t2785 8.47023
R20493 VGND.n2235 VGND.t1453 8.47023
R20494 VGND.n2233 VGND.t1451 8.47023
R20495 VGND.n2231 VGND.t1449 8.47023
R20496 VGND.n2229 VGND.t1447 8.47023
R20497 VGND.n2228 VGND.t3423 8.47023
R20498 VGND.n2225 VGND.t3421 8.47023
R20499 VGND.n426 VGND.t4975 8.47023
R20500 VGND.n2451 VGND.t4973 8.47023
R20501 VGND.n2452 VGND.t1297 8.47023
R20502 VGND.n2455 VGND.t1295 8.47023
R20503 VGND.n2456 VGND.t5758 8.47023
R20504 VGND.n2459 VGND.t5756 8.47023
R20505 VGND.n2532 VGND.t4969 8.47023
R20506 VGND.n2530 VGND.t4971 8.47023
R20507 VGND.n2529 VGND.t943 8.47023
R20508 VGND.n2527 VGND.t945 8.47023
R20509 VGND.n2525 VGND.t4496 8.47023
R20510 VGND.n2522 VGND.t4494 8.47023
R20511 VGND.n2520 VGND.t3910 8.47023
R20512 VGND.n2518 VGND.t3912 8.47023
R20513 VGND.n2517 VGND.t2248 8.47023
R20514 VGND.n2515 VGND.t2250 8.47023
R20515 VGND.n2519 VGND.t5404 8.47023
R20516 VGND.n2521 VGND.t5402 8.47023
R20517 VGND.n2089 VGND.t1674 8.46241
R20518 VGND.n2050 VGND.t1808 8.46241
R20519 VGND.n194 VGND.t4242 8.46241
R20520 VGND.n163 VGND.t6811 8.46241
R20521 VGND.n1415 VGND.t820 8.46241
R20522 VGND.n873 VGND.t2314 8.46241
R20523 VGND.n875 VGND.t2313 8.46241
R20524 VGND.n834 VGND.t5101 8.46241
R20525 VGND.n1312 VGND.t3615 8.46241
R20526 VGND.n1572 VGND.t4295 8.46241
R20527 VGND.n1380 VGND.t1946 8.46241
R20528 VGND.n1378 VGND.t1948 8.46241
R20529 VGND.n3427 VGND.t3378 8.46241
R20530 VGND.n3425 VGND.t3380 8.46241
R20531 VGND.n3417 VGND.t3057 8.46241
R20532 VGND.n1565 VGND.t6037 8.46241
R20533 VGND.n1545 VGND.t5593 8.46241
R20534 VGND.n3394 VGND.t612 8.46241
R20535 VGND.n3383 VGND.t400 8.46241
R20536 VGND.n3402 VGND.t928 8.46241
R20537 VGND.n1553 VGND.t804 8.46241
R20538 VGND.n1480 VGND.t3225 8.46241
R20539 VGND.n1661 VGND.t2156 8.46241
R20540 VGND.n1687 VGND.t3961 8.46241
R20541 VGND.n1688 VGND.t3957 8.46241
R20542 VGND.n1782 VGND.t3838 8.46241
R20543 VGND.n1744 VGND.t3851 8.46241
R20544 VGND.n1756 VGND.t5633 8.46241
R20545 VGND.n1767 VGND.t4052 8.46241
R20546 VGND.n1787 VGND.t3729 8.46241
R20547 VGND.n1789 VGND.t3727 8.46241
R20548 VGND.n1127 VGND.t4759 8.46241
R20549 VGND.n759 VGND.t1920 8.46241
R20550 VGND.n1804 VGND.t2643 8.46241
R20551 VGND.n766 VGND.t5473 8.46241
R20552 VGND.n1950 VGND.t6503 8.46241
R20553 VGND.n1126 VGND.t6508 8.46241
R20554 VGND.n1977 VGND.t1217 8.46241
R20555 VGND.n1911 VGND.t5784 8.46241
R20556 VGND.n1927 VGND.t6521 8.46241
R20557 VGND.n1981 VGND.t3101 8.46241
R20558 VGND.n470 VGND.t4419 8.46241
R20559 VGND.n2400 VGND.t1828 8.46241
R20560 VGND.n482 VGND.t6501 8.46241
R20561 VGND.n2204 VGND.t5501 8.46241
R20562 VGND.n2180 VGND.t584 8.46241
R20563 VGND.n2179 VGND.t588 8.46241
R20564 VGND.n2402 VGND.t2760 8.46241
R20565 VGND.n2404 VGND.t2758 8.46241
R20566 VGND.n516 VGND.t4017 8.46241
R20567 VGND.n2368 VGND.t6003 8.46241
R20568 VGND.n2369 VGND.t5088 8.46241
R20569 VGND.n2370 VGND.t5084 8.46241
R20570 VGND.n1626 VGND.t5534 8.44089
R20571 VGND.n1640 VGND.t330 8.44089
R20572 VGND.n1215 VGND.t2591 8.44089
R20573 VGND.n1218 VGND.t2466 8.44089
R20574 VGND.n587 VGND.t4655 8.43502
R20575 VGND.n1976 VGND.t4649 8.43502
R20576 VGND.n219 VGND.t4866 8.42575
R20577 VGND.n864 VGND.t2447 8.42575
R20578 VGND.n312 VGND.t5793 8.42575
R20579 VGND.n1297 VGND.t4120 8.42575
R20580 VGND.n1481 VGND.t787 8.42575
R20581 VGND.n253 VGND.t394 8.42575
R20582 VGND.n2037 VGND.t4531 8.4135
R20583 VGND.n2052 VGND.t3980 8.4135
R20584 VGND.n2056 VGND.t3982 8.4135
R20585 VGND.n2061 VGND.t6421 8.4135
R20586 VGND.n2078 VGND.t939 8.4135
R20587 VGND.n2062 VGND.t6023 8.4135
R20588 VGND.n2033 VGND.t4309 8.4135
R20589 VGND.n124 VGND.t35 8.4135
R20590 VGND.n171 VGND.t6297 8.4135
R20591 VGND.n225 VGND.t6590 8.4135
R20592 VGND.n1315 VGND.t5057 8.4135
R20593 VGND.n1585 VGND.t5779 8.4135
R20594 VGND.n1576 VGND.t1016 8.4135
R20595 VGND.n311 VGND.t2601 8.4135
R20596 VGND.n1587 VGND.t3678 8.4135
R20597 VGND.n1590 VGND.t4193 8.4135
R20598 VGND.n1344 VGND.t3611 8.4135
R20599 VGND.n1309 VGND.t6344 8.4135
R20600 VGND.n1247 VGND.t3887 8.4135
R20601 VGND.n1600 VGND.t2698 8.4135
R20602 VGND.n1452 VGND.t1252 8.4135
R20603 VGND.n1471 VGND.t1256 8.4135
R20604 VGND.n1504 VGND.t6667 8.4135
R20605 VGND.n3395 VGND.t3483 8.4135
R20606 VGND.n3386 VGND.t3481 8.4135
R20607 VGND.n1512 VGND.t4415 8.4135
R20608 VGND.n1520 VGND.t469 8.4135
R20609 VGND.n1467 VGND.t6435 8.4135
R20610 VGND.n1677 VGND.t5748 8.4135
R20611 VGND.n1691 VGND.t6152 8.4135
R20612 VGND.n1692 VGND.t3122 8.4135
R20613 VGND.n1784 VGND.t467 8.4135
R20614 VGND.n1768 VGND.t6676 8.4135
R20615 VGND.n1701 VGND.t3417 8.4135
R20616 VGND.n1941 VGND.t6574 8.4135
R20617 VGND.n757 VGND.t5850 8.4135
R20618 VGND.n1967 VGND.t1189 8.4135
R20619 VGND.n641 VGND.t5745 8.4135
R20620 VGND.n638 VGND.t4316 8.4135
R20621 VGND.n1978 VGND.t302 8.4135
R20622 VGND.n2386 VGND.t6121 8.4135
R20623 VGND.n2178 VGND.t3253 8.4135
R20624 VGND.n2185 VGND.t5371 8.4135
R20625 VGND.n511 VGND.t6128 8.4135
R20626 VGND.n1462 VGND.t6432 8.41154
R20627 VGND.n1528 VGND.t3329 8.41154
R20628 VGND.n1763 VGND.t6136 8.41154
R20629 VGND.n866 VGND.t2481 8.4101
R20630 VGND.n1299 VGND.t6563 8.4101
R20631 VGND.n1478 VGND.t209 8.4101
R20632 VGND.n551 VGND.t3859 8.4005
R20633 VGND.n551 VGND.t3861 8.4005
R20634 VGND.n562 VGND.t1008 8.4005
R20635 VGND.n562 VGND.t5356 8.4005
R20636 VGND.n227 VGND.t1285 8.4005
R20637 VGND.n227 VGND.t1286 8.4005
R20638 VGND.n181 VGND.t5076 8.4005
R20639 VGND.n181 VGND.t2262 8.4005
R20640 VGND.n160 VGND.t1841 8.4005
R20641 VGND.n160 VGND.t424 8.4005
R20642 VGND.n1402 VGND.t5092 8.4005
R20643 VGND.n1402 VGND.t3001 8.4005
R20644 VGND.n870 VGND.t860 8.4005
R20645 VGND.n870 VGND.t4083 8.4005
R20646 VGND.n1357 VGND.t4931 8.4005
R20647 VGND.n1357 VGND.t1413 8.4005
R20648 VGND.n1373 VGND.t4789 8.4005
R20649 VGND.n1373 VGND.t4498 8.4005
R20650 VGND.n148 VGND.t4849 8.4005
R20651 VGND.n148 VGND.t4366 8.4005
R20652 VGND.n155 VGND.t1533 8.4005
R20653 VGND.n155 VGND.t1689 8.4005
R20654 VGND.n275 VGND.t2506 8.4005
R20655 VGND.n275 VGND.t1788 8.4005
R20656 VGND.n1361 VGND.t2839 8.4005
R20657 VGND.n1361 VGND.t1545 8.4005
R20658 VGND.n1489 VGND.t891 8.4005
R20659 VGND.n1489 VGND.t4862 8.4005
R20660 VGND.n204 VGND.t4087 8.4005
R20661 VGND.n204 VGND.t1596 8.4005
R20662 VGND.n248 VGND.t930 8.4005
R20663 VGND.n248 VGND.t5844 8.4005
R20664 VGND.n201 VGND.t5185 8.4005
R20665 VGND.n201 VGND.t2895 8.4005
R20666 VGND.n1486 VGND.t528 8.4005
R20667 VGND.n1486 VGND.t5278 8.4005
R20668 VGND.n1474 VGND.t4423 8.4005
R20669 VGND.n1474 VGND.t2819 8.4005
R20670 VGND.n792 VGND.t5579 8.4005
R20671 VGND.n792 VGND.t5170 8.4005
R20672 VGND.n775 VGND.t2515 8.4005
R20673 VGND.n775 VGND.t3479 8.4005
R20674 VGND.n1732 VGND.t1334 8.4005
R20675 VGND.n1732 VGND.t5737 8.4005
R20676 VGND.n1728 VGND.t4590 8.4005
R20677 VGND.n1728 VGND.t4934 8.4005
R20678 VGND.n1723 VGND.t2828 8.4005
R20679 VGND.n1723 VGND.t912 8.4005
R20680 VGND.n1717 VGND.t5891 8.4005
R20681 VGND.n1717 VGND.t426 8.4005
R20682 VGND.n730 VGND.t5446 8.4005
R20683 VGND.n730 VGND.t453 8.4005
R20684 VGND.n723 VGND.t2973 8.4005
R20685 VGND.n723 VGND.t2220 8.4005
R20686 VGND.n727 VGND.t530 8.4005
R20687 VGND.n727 VGND.t3754 8.4005
R20688 VGND.n582 VGND.t2800 8.4005
R20689 VGND.n582 VGND.t2798 8.4005
R20690 VGND.n664 VGND.t3576 8.4005
R20691 VGND.n664 VGND.t1956 8.4005
R20692 VGND.n580 VGND.t5894 8.4005
R20693 VGND.n580 VGND.t987 8.4005
R20694 VGND.n946 VGND.t2605 8.4005
R20695 VGND.n946 VGND.t922 8.4005
R20696 VGND.n477 VGND.t1821 8.4005
R20697 VGND.n477 VGND.t457 8.4005
R20698 VGND.n2197 VGND.t1612 8.4005
R20699 VGND.n2197 VGND.t2032 8.4005
R20700 VGND.n481 VGND.t2560 8.4005
R20701 VGND.n481 VGND.t5770 8.4005
R20702 VGND.n471 VGND.t1384 8.4005
R20703 VGND.n471 VGND.t3081 8.4005
R20704 VGND.n509 VGND.t48 8.4005
R20705 VGND.n509 VGND.t4941 8.4005
R20706 VGND.n528 VGND.t4226 8.4005
R20707 VGND.n528 VGND.t1746 8.4005
R20708 VGND.n524 VGND.t1515 8.4005
R20709 VGND.n524 VGND.t1513 8.4005
R20710 VGND.n1513 VGND.t6292 8.38415
R20711 VGND.n178 VGND.t868 8.37615
R20712 VGND.n1472 VGND.t1539 8.37615
R20713 VGND.n2036 VGND.t4307 8.3563
R20714 VGND.n323 VGND.t2597 8.3563
R20715 VGND.n1385 VGND.t6542 8.3563
R20716 VGND.n1458 VGND.t6437 8.3563
R20717 VGND.n1524 VGND.t3331 8.3563
R20718 VGND.n1664 VGND.t113 8.3563
R20719 VGND.n1766 VGND.t6139 8.3563
R20720 VGND.n2406 VGND.t136 8.3563
R20721 VGND.n2058 VGND.t6425 8.35306
R20722 VGND VGND.t1191 8.35306
R20723 VGND.n2086 VGND.t1672 8.0855
R20724 VGND.n564 VGND.t1810 8.0855
R20725 VGND.n180 VGND.t4241 8.0855
R20726 VGND.n161 VGND.t6812 8.0855
R20727 VGND.n1401 VGND.t819 8.0855
R20728 VGND.n871 VGND.t2315 8.0855
R20729 VGND.n1356 VGND.t4297 8.0855
R20730 VGND.n1372 VGND.t1950 8.0855
R20731 VGND.n146 VGND.t3382 8.0855
R20732 VGND.n153 VGND.t3059 8.0855
R20733 VGND.n1358 VGND.t6039 8.0855
R20734 VGND.n1488 VGND.t5591 8.0855
R20735 VGND.n199 VGND.t926 8.0855
R20736 VGND.n1485 VGND.t802 8.0855
R20737 VGND.n1473 VGND.t3227 8.0855
R20738 VGND.n203 VGND.t610 8.0855
R20739 VGND.n789 VGND.t2158 8.0855
R20740 VGND.n774 VGND.t3959 8.0855
R20741 VGND.n1730 VGND.t3853 8.0855
R20742 VGND.n1726 VGND.t5631 8.0855
R20743 VGND.n1722 VGND.t4050 8.0855
R20744 VGND.n768 VGND.t3731 8.0855
R20745 VGND.n731 VGND.t1922 8.0855
R20746 VGND.n724 VGND.t2645 8.0855
R20747 VGND.n728 VGND.t5475 8.0855
R20748 VGND.n584 VGND.t1219 8.0855
R20749 VGND.n663 VGND.t5786 8.0855
R20750 VGND.n581 VGND.t3103 8.0855
R20751 VGND.n949 VGND.t4417 8.0855
R20752 VGND.n475 VGND.t1830 8.0855
R20753 VGND.n2194 VGND.t5503 8.0855
R20754 VGND.n2176 VGND.t586 8.0855
R20755 VGND.n473 VGND.t2762 8.0855
R20756 VGND.n508 VGND.t4019 8.0855
R20757 VGND.n527 VGND.t6001 8.0855
R20758 VGND.n526 VGND.t5086 8.0855
R20759 VGND.n3755 VGND.n3 7.4975
R20760 VGND.n803 VGND.t5053 7.37611
R20761 VGND.n805 VGND.t6346 7.37611
R20762 VGND.n281 VGND.t6589 7.37611
R20763 VGND.n778 VGND.t5384 7.37611
R20764 VGND.n622 VGND.t4998 7.37611
R20765 VGND.n209 VGND.t4869 6.64191
R20766 VGND.n277 VGND.t5791 6.64191
R20767 VGND.n249 VGND.t396 6.64191
R20768 VGND.n807 VGND.t20 6.63343
R20769 VGND.n806 VGND.t5 6.63343
R20770 VGND.n212 VGND.t6225 6.63343
R20771 VGND.n553 VGND.t6150 6.56999
R20772 VGND.n549 VGND.t2450 6.56999
R20773 VGND.n286 VGND.t4732 6.56999
R20774 VGND.n285 VGND.t1181 6.56999
R20775 VGND.n844 VGND.t178 6.56999
R20776 VGND.n733 VGND.t6548 6.56999
R20777 VGND.n1814 VGND.t166 6.56999
R20778 VGND.n1125 VGND.t717 6.56999
R20779 VGND.n662 VGND.t6111 6.56999
R20780 VGND.n2195 VGND.t2570 6.56999
R20781 VGND.n2087 VGND.n2086 6.54898
R20782 VGND.n2051 VGND.n564 6.54898
R20783 VGND.n192 VGND.n180 6.54898
R20784 VGND.n165 VGND.n161 6.54898
R20785 VGND.n1413 VGND.n1401 6.54898
R20786 VGND.n876 VGND.n871 6.54898
R20787 VGND.n1570 VGND.n1356 6.54898
R20788 VGND.n1376 VGND.n1372 6.54898
R20789 VGND.n3424 VGND.n146 6.54898
R20790 VGND.n3415 VGND.n153 6.54898
R20791 VGND.n1564 VGND.n1358 6.54898
R20792 VGND.n1543 VGND.n1488 6.54898
R20793 VGND.n3400 VGND.n199 6.54898
R20794 VGND.n1552 VGND.n1485 6.54898
R20795 VGND.n1479 VGND.n1473 6.54898
R20796 VGND VGND.n203 6.54898
R20797 VGND.n1660 VGND.n789 6.54898
R20798 VGND.n1686 VGND.n774 6.54898
R20799 VGND.n1742 VGND.n1730 6.54898
R20800 VGND.n1754 VGND.n1726 6.54898
R20801 VGND.n1765 VGND.n1722 6.54898
R20802 VGND.n1785 VGND.n768 6.54898
R20803 VGND.n760 VGND.n731 6.54898
R20804 VGND.n1805 VGND.n724 6.54898
R20805 VGND VGND.n728 6.54898
R20806 VGND.n1979 VGND.n584 6.54898
R20807 VGND.n1909 VGND.n663 6.54898
R20808 VGND.n1983 VGND.n581 6.54898
R20809 VGND.n951 VGND.n949 6.54898
R20810 VGND.n2398 VGND.n475 6.54898
R20811 VGND.n2203 VGND.n2194 6.54898
R20812 VGND.n2177 VGND.n2176 6.54898
R20813 VGND.n2405 VGND.n473 6.54898
R20814 VGND.n514 VGND.n508 6.54898
R20815 VGND.n2367 VGND.n527 6.54898
R20816 VGND.n2371 VGND.n526 6.54898
R20817 VGND.n822 VGND.n801 6.54311
R20818 VGND.n1530 VGND.n1493 6.54311
R20819 VGND.n1773 VGND.n1719 6.54311
R20820 VGND.n1914 VGND.n661 6.54311
R20821 VGND.n2184 VGND.n2173 6.54311
R20822 VGND.n2372 VGND.n525 6.54311
R20823 VGND.n566 VGND.t3984 6.5255
R20824 VGND.n848 VGND.t3613 6.5255
R20825 VGND.n738 VGND.t6636 6.5255
R20826 VGND.n658 VGND.t5598 6.5255
R20827 VGND.n826 VGND.t6747 6.50373
R20828 VGND.n898 VGND.t6692 6.50373
R20829 VGND.n1345 VGND.n1338 6.47463
R20830 VGND.n2160 VGND.n2094 6.46859
R20831 VGND.n2059 VGND.n561 6.46859
R20832 VGND.n237 VGND.n228 6.46859
R20833 VGND.n185 VGND.n182 6.46859
R20834 VGND.n173 VGND.n159 6.46859
R20835 VGND.n1405 VGND.n1403 6.46859
R20836 VGND.n884 VGND.n868 6.46859
R20837 VGND.n1399 VGND.n1359 6.46859
R20838 VGND.n3430 VGND.n142 6.46859
R20839 VGND.n3419 VGND.n150 6.46859
R20840 VGND.n157 VGND.n156 6.46859
R20841 VGND.n327 VGND.n274 6.46859
R20842 VGND.n1392 VGND.n1363 6.46859
R20843 VGND.n1535 VGND.n1491 6.46859
R20844 VGND.n3385 VGND.n207 6.46859
R20845 VGND.n266 VGND.n247 6.46859
R20846 VGND.n3392 VGND.n202 6.46859
R20847 VGND.n1544 VGND.n1487 6.46859
R20848 VGND.n1557 VGND.n1444 6.46859
R20849 VGND.n1651 VGND.n795 6.46859
R20850 VGND.n1680 VGND.n777 6.46859
R20851 VGND.n1759 VGND.n1724 6.46859
R20852 VGND.n1734 VGND.n1733 6.46859
R20853 VGND.n1748 VGND.n1729 6.46859
R20854 VGND.n1778 VGND.n1718 6.46859
R20855 VGND.n1795 VGND.n729 6.46859
R20856 VGND.n1821 VGND.n1813 6.46859
R20857 VGND.n1802 VGND.n725 6.46859
R20858 VGND.n1986 VGND.n579 6.46859
R20859 VGND.n1901 VGND.n666 6.46859
R20860 VGND.n1990 VGND.n578 6.46859
R20861 VGND.n957 VGND.n945 6.46859
R20862 VGND.n2390 VGND.n479 6.46859
R20863 VGND.n2218 VGND.n2171 6.46859
R20864 VGND.n2389 VGND.n480 6.46859
R20865 VGND.n952 VGND.n948 6.46859
R20866 VGND.n2378 VGND.n487 6.46859
R20867 VGND.n2358 VGND.n530 6.46859
R20868 VGND.n2379 VGND.n486 6.46859
R20869 VGND.n2046 VGND.n566 6.46462
R20870 VGND.n1440 VGND.n1421 6.46462
R20871 VGND.n860 VGND.n848 6.46462
R20872 VGND.n1674 VGND.n780 6.46462
R20873 VGND.n1673 VGND.n781 6.46462
R20874 VGND.n1672 VGND.n782 6.46462
R20875 VGND.n1962 VGND.n595 6.46462
R20876 VGND.n1960 VGND.n597 6.46462
R20877 VGND.n1958 VGND.n598 6.46462
R20878 VGND.n743 VGND.n738 6.46462
R20879 VGND.n639 VGND.n621 6.46462
R20880 VGND.n641 VGND.n620 6.46462
R20881 VGND.n642 VGND.n619 6.46462
R20882 VGND.n1924 VGND.n658 6.46462
R20883 VGND.n1505 VGND.n1501 6.45932
R20884 VGND.n924 VGND.n919 6.45138
R20885 VGND.n853 VGND.n850 6.45138
R20886 VGND.n3446 VGND.n113 6.45138
R20887 VGND.n1433 VGND.n1425 6.45138
R20888 VGND.n1435 VGND.n1423 6.45138
R20889 VGND.n1436 VGND.n1422 6.45138
R20890 VGND.n931 VGND.n918 6.45138
R20891 VGND.n1393 VGND.n1362 6.45138
R20892 VGND.n1459 VGND.n1447 6.45138
R20893 VGND.n1668 VGND.n784 6.45138
R20894 VGND.n1666 VGND.n786 6.45138
R20895 VGND.n1663 VGND.n787 6.45138
R20896 VGND.n1662 VGND.n788 6.45138
R20897 VGND.n1659 VGND.n790 6.45138
R20898 VGND.n1658 VGND.n791 6.45138
R20899 VGND.n1656 VGND.n793 6.45138
R20900 VGND.n1954 VGND.n601 6.45138
R20901 VGND.n1952 VGND.n602 6.45138
R20902 VGND.n1951 VGND.n603 6.45138
R20903 VGND.n1949 VGND.n604 6.45138
R20904 VGND.n1947 VGND.n606 6.45138
R20905 VGND.n1946 VGND.n607 6.45138
R20906 VGND.n1944 VGND.n609 6.45138
R20907 VGND.n652 VGND.n645 6.45138
R20908 VGND.n651 VGND.n646 6.45138
R20909 VGND.n650 VGND.n647 6.45138
R20910 VGND.n649 VGND.n648 6.45138
R20911 VGND.n614 VGND.n613 6.45138
R20912 VGND.n1935 VGND.n616 6.45138
R20913 VGND.n1934 VGND.n617 6.45138
R20914 VGND.n811 VGND.n807 6.45115
R20915 VGND.n814 VGND.n806 6.45115
R20916 VGND.n217 VGND.n212 6.45115
R20917 VGND.n1508 VGND.n1500 6.45006
R20918 VGND.n1621 VGND.n842 6.44333
R20919 VGND.n1624 VGND.n841 6.44333
R20920 VGND.n1642 VGND.n797 6.44333
R20921 VGND.n1210 VGND.n1207 6.44333
R20922 VGND.n1213 VGND.n1205 6.44333
R20923 VGND.n1220 VGND.n1204 6.44333
R20924 VGND.n1223 VGND.n1203 6.44333
R20925 VGND VGND.n796 6.44333
R20926 VGND.n1580 VGND.n1352 6.44137
R20927 VGND.n1584 VGND.n1350 6.44137
R20928 VGND.n1466 VGND.n1446 6.44137
R20929 VGND.n753 VGND.n734 6.44137
R20930 VGND.n749 VGND.n735 6.44137
R20931 VGND.n1929 VGND.n657 6.44137
R20932 VGND.n2054 VGND.n563 6.4355
R20933 VGND.n1582 VGND.n1351 6.4355
R20934 VGND.n3413 VGND.n154 6.4355
R20935 VGND.n1302 VGND.n896 6.4355
R20936 VGND.n1211 VGND.n1206 6.4355
R20937 VGND.n748 VGND.n736 6.4355
R20938 VGND.n1817 VGND.n1815 6.4355
R20939 VGND.n1957 VGND.n599 6.4355
R20940 VGND.n1975 VGND.n585 6.4355
R20941 VGND.n820 VGND.n803 6.43354
R20942 VGND.n817 VGND.n805 6.43354
R20943 VGND.n313 VGND.n281 6.43354
R20944 VGND.n1678 VGND.n778 6.43354
R20945 VGND.n634 VGND.n622 6.43354
R20946 VGND.n882 VGND.n869 6.41829
R20947 VGND.n1430 VGND.n1427 6.41829
R20948 VGND.n854 VGND.n849 6.41789
R20949 VGND.n1327 VGND.n890 6.41789
R20950 VGND.n1332 VGND.n889 6.41789
R20951 VGND.n1333 VGND.n888 6.41789
R20952 VGND.n1611 VGND.n843 6.41789
R20953 VGND.n2079 VGND.n553 6.41593
R20954 VGND.n550 VGND.n549 6.41593
R20955 VGND.n223 VGND.n210 6.41593
R20956 VGND VGND.n209 6.41593
R20957 VGND.n297 VGND.n286 6.41593
R20958 VGND.n319 VGND.n277 6.41593
R20959 VGND.n317 VGND.n279 6.41593
R20960 VGND.n298 VGND.n285 6.41593
R20961 VGND.n259 VGND.n249 6.41593
R20962 VGND.n257 VGND.n251 6.41593
R20963 VGND.n845 VGND.n844 6.41593
R20964 VGND.n756 VGND.n733 6.41593
R20965 VGND.n1818 VGND.n1814 6.41593
R20966 VGND.n1128 VGND.n1125 6.41593
R20967 VGND.n1910 VGND.n662 6.41593
R20968 VGND.n2202 VGND.n2195 6.41593
R20969 VGND.n2164 VGND.n552 6.40771
R20970 VGND.n126 VGND.n123 6.40771
R20971 VGND.n1341 VGND.n1339 6.40771
R20972 VGND.n299 VGND.n284 6.40771
R20973 VGND.n1575 VGND.n1353 6.40771
R20974 VGND.n1503 VGND.n1502 6.40771
R20975 VGND.n3389 VGND.n205 6.40771
R20976 VGND.n1752 VGND.n1727 6.40771
R20977 VGND.n1772 VGND.n1720 6.40771
R20978 VGND.n1709 VGND.n769 6.40771
R20979 VGND.n1704 VGND.n770 6.40771
R20980 VGND.n1930 VGND.n656 6.40771
R20981 VGND.n1915 VGND.n660 6.40771
R20982 VGND.n630 VGND.n624 6.40771
R20983 VGND.n2182 VGND.n2174 6.40771
R20984 VGND.n2200 VGND.n2196 6.40771
R20985 VGND.n2219 VGND.n2170 6.40771
R20986 VGND.n2395 VGND.n476 6.40771
R20987 VGND.n2375 VGND.n523 6.40771
R20988 VGND.n2038 VGND.n569 6.39182
R20989 VGND.n321 VGND.n276 6.39182
R20990 VGND.n1382 VGND.n1369 6.39182
R20991 VGND.n1667 VGND.n785 6.39182
R20992 VGND.n1955 VGND.n600 6.39182
R20993 VGND.n1974 VGND.n586 6.39182
R20994 VGND.n2403 VGND.n474 6.39182
R20995 VGND.n830 VGND.n826 6.38785
R20996 VGND.n1296 VGND.n898 6.38785
R20997 VGND.n2063 VGND.n559 6.38659
R20998 VGND.n916 VGND.n909 6.38659
R20999 VGND.n821 VGND.n802 6.38659
R21000 VGND.n823 VGND.n800 6.38659
R21001 VGND.n861 VGND.n847 6.38659
R21002 VGND.n741 VGND.n740 6.38659
R21003 VGND.n1961 VGND.n596 6.38659
R21004 VGND.n1305 VGND.n893 6.38521
R21005 VGND.n1307 VGND.n892 6.38521
R21006 VGND.n1455 VGND.n1449 6.38521
R21007 VGND.n1454 VGND.n1450 6.38521
R21008 VGND.n1968 VGND.n591 6.38521
R21009 VGND.n1966 VGND.n592 6.38521
R21010 VGND VGND.n1424 6.37859
R21011 VGND.n221 VGND.n211 6.37859
R21012 VGND.n176 VGND.n158 6.37859
R21013 VGND VGND.n897 6.37859
R21014 VGND.n314 VGND.n280 6.37859
R21015 VGND.n1387 VGND.n1366 6.37859
R21016 VGND.n1389 VGND.n1364 6.37859
R21017 VGND VGND.n1492 6.37859
R21018 VGND.n256 VGND.n252 6.37859
R21019 VGND.n1469 VGND.n1445 6.37859
R21020 VGND VGND.n722 6.37859
R21021 VGND VGND.n2172 6.37859
R21022 VGND.n742 VGND.n739 6.36006
R21023 VGND.n1963 VGND.n594 6.36006
R21024 VGND.n633 VGND.n623 6.36006
R21025 VGND.n2034 VGND.n571 6.35874
R21026 VGND.n2043 VGND.n568 6.35874
R21027 VGND.n2065 VGND.n557 6.35874
R21028 VGND.n2067 VGND.n556 6.35874
R21029 VGND.n2064 VGND.n558 6.35874
R21030 VGND.n912 VGND.n910 6.35874
R21031 VGND.n818 VGND.n804 6.35874
R21032 VGND.n835 VGND.n825 6.35874
R21033 VGND.n865 VGND.n846 6.35874
R21034 VGND.n1430 VGND.n1426 6.35874
R21035 VGND.n1429 VGND.n1428 6.35874
R21036 VGND.n3449 VGND.n112 6.35874
R21037 VGND.n3440 VGND.n114 6.35874
R21038 VGND.n3439 VGND.n115 6.35874
R21039 VGND.n132 VGND.n119 6.35874
R21040 VGND.n130 VGND.n121 6.35874
R21041 VGND.n127 VGND.n122 6.35874
R21042 VGND.n131 VGND.n120 6.35874
R21043 VGND.n133 VGND.n118 6.35874
R21044 VGND.n135 VGND.n117 6.35874
R21045 VGND.n3438 VGND.n116 6.35874
R21046 VGND.n1388 VGND.n1365 6.35874
R21047 VGND.n1386 VGND.n1367 6.35874
R21048 VGND.n1384 VGND.n1368 6.35874
R21049 VGND.n3421 VGND.n149 6.35874
R21050 VGND.n3423 VGND.n147 6.35874
R21051 VGND.n1628 VGND.n839 6.35874
R21052 VGND.n1453 VGND.n1451 6.35874
R21053 VGND.n1522 VGND.n1495 6.35874
R21054 VGND.n1521 VGND.n1496 6.35874
R21055 VGND.n1518 VGND.n1497 6.35874
R21056 VGND.n1511 VGND.n1498 6.35874
R21057 VGND.n1248 VGND.n1246 6.35874
R21058 VGND.n1676 VGND.n779 6.35874
R21059 VGND.n1693 VGND.n772 6.35874
R21060 VGND.n1690 VGND.n773 6.35874
R21061 VGND.n590 VGND.n589 6.35874
R21062 VGND.n1942 VGND.n610 6.35874
R21063 VGND.n1945 VGND.n608 6.35874
R21064 VGND.n1933 VGND.n618 6.35874
R21065 VGND.n1936 VGND.n615 6.35874
R21066 VGND.n953 VGND.n947 6.35874
R21067 VGND.n296 VGND.n287 6.3555
R21068 VGND.n293 VGND.n288 6.3555
R21069 VGND.n3426 VGND.n145 6.3555
R21070 VGND.n3429 VGND.n143 6.3555
R21071 VGND.n569 VGND.t306 6.32611
R21072 VGND.n276 VGND.t6583 6.32611
R21073 VGND.n1369 VGND.t6429 6.32611
R21074 VGND.n785 VGND.t13 6.32611
R21075 VGND.n599 VGND.t1254 6.32611
R21076 VGND.n585 VGND.t134 6.32611
R21077 VGND.n474 VGND.t4653 6.32611
R21078 VGND.n869 VGND.t2011 5.79141
R21079 VGND.n1427 VGND.t3073 5.79141
R21080 VGND.n559 VGND.t5981 5.66271
R21081 VGND.n740 VGND.t3591 5.66271
R21082 VGND.n1500 VGND.t3429 5.43579
R21083 VGND.n596 VGND.t5386 5.38302
R21084 VGND VGND.n2922 5.32526
R21085 VGND.n2060 VGND.n560 5.32359
R21086 VGND.n2048 VGND.n565 5.32359
R21087 VGND.n2035 VGND.n570 5.32359
R21088 VGND.n2019 VGND.n572 5.32359
R21089 VGND.n1030 VGND.n1023 5.32359
R21090 VGND.n1050 VGND.n1022 5.32359
R21091 VGND.n3348 VGND.n357 5.32359
R21092 VGND.n2105 VGND.n2096 5.32359
R21093 VGND VGND.t2112 5.32359
R21094 VGND.n2141 VGND.t2741 5.32359
R21095 VGND.n2158 VGND.n2095 5.32359
R21096 VGND.n2092 VGND.n2091 5.32359
R21097 VGND.n2071 VGND.n554 5.32359
R21098 VGND.n3452 VGND.n3451 5.32359
R21099 VGND.n3451 VGND.n111 5.32359
R21100 VGND.n3451 VGND.n61 5.32359
R21101 VGND.n3451 VGND 5.32359
R21102 VGND.n3451 VGND.n60 5.32359
R21103 VGND.n3451 VGND.n59 5.32359
R21104 VGND.n3451 VGND.n58 5.32359
R21105 VGND.n3451 VGND.n57 5.32359
R21106 VGND.n3451 VGND.n56 5.32359
R21107 VGND.n3451 VGND 5.32359
R21108 VGND.n3691 VGND.n42 5.32359
R21109 VGND.n1377 VGND.n1371 5.32359
R21110 VGND.n1573 VGND.n1355 5.32359
R21111 VGND.n1348 VGND.n1347 5.32359
R21112 VGND.n3416 VGND.n152 5.32359
R21113 VGND.n340 VGND.n246 5.32359
R21114 VGND.n306 VGND.n282 5.32359
R21115 VGND.n1304 VGND.n894 5.32359
R21116 VGND.n3388 VGND.n206 5.32359
R21117 VGND.n1510 VGND.n1499 5.32359
R21118 VGND.n1539 VGND.n1490 5.32359
R21119 VGND.n1483 VGND.n1482 5.32359
R21120 VGND.n1607 VGND.t4319 5.32359
R21121 VGND.n1255 VGND.t4376 5.32359
R21122 VGND.n1741 VGND.n1731 5.32359
R21123 VGND.n1769 VGND.n1721 5.32359
R21124 VGND.n1684 VGND.n776 5.32359
R21125 VGND.n1654 VGND.n794 5.32359
R21126 VGND.n1217 VGND.t3760 5.32359
R21127 VGND.t3013 VGND 5.32359
R21128 VGND.n1852 VGND.t2265 5.32359
R21129 VGND.n1823 VGND.n1822 5.32359
R21130 VGND.n758 VGND.n732 5.32359
R21131 VGND.n1948 VGND.n605 5.32359
R21132 VGND.n1130 VGND.n1124 5.32359
R21133 VGND.n1163 VGND.n1123 5.32359
R21134 VGND.n654 VGND.n653 5.32359
R21135 VGND.n1980 VGND.n583 5.32359
R21136 VGND.n695 VGND.t4944 5.32359
R21137 VGND.n1889 VGND.t4174 5.32359
R21138 VGND.n1922 VGND.n659 5.32359
R21139 VGND.n1087 VGND.n1077 5.32359
R21140 VGND.n2393 VGND.n478 5.32359
R21141 VGND.n958 VGND.n944 5.32359
R21142 VGND.n998 VGND.n942 5.32359
R21143 VGND.n2206 VGND 5.32359
R21144 VGND.t418 VGND.n2862 5.32359
R21145 VGND.n2571 VGND.t5917 5.32359
R21146 VGND.n2795 VGND.t4378 5.32359
R21147 VGND.t5346 VGND.n2766 5.32359
R21148 VGND.n2643 VGND.n2634 5.32359
R21149 VGND.n2662 VGND.n2632 5.32359
R21150 VGND.n2698 VGND.t2656 5.32359
R21151 VGND.n2715 VGND.n2631 5.32359
R21152 VGND.n2629 VGND.n2628 5.32359
R21153 VGND VGND.t5556 5.32359
R21154 VGND.n2362 VGND.n529 5.32359
R21155 VGND.n521 VGND.n520 5.32359
R21156 VGND.n2427 VGND.t1917 5.32359
R21157 VGND.n466 VGND.n465 5.32359
R21158 VGND.t852 VGND.n2331 5.32359
R21159 VGND.n2284 VGND.t2204 5.32359
R21160 VGND.n2247 VGND.t6808 5.32359
R21161 VGND.n2464 VGND.t5193 5.32359
R21162 VGND.n2911 VGND.n404 5.32359
R21163 VGND.n2502 VGND.n2497 5.32359
R21164 VGND.n2533 VGND.n2494 5.32359
R21165 VGND.t5221 VGND 5.32359
R21166 VGND.n3737 VGND.n6 5.32359
R21167 VGND.n3324 VGND.n3312 5.32359
R21168 VGND.n3291 VGND.n361 5.32359
R21169 VGND.n3196 VGND.n3182 5.32359
R21170 VGND.n3162 VGND.n368 5.32359
R21171 VGND.n3091 VGND.n3076 5.32359
R21172 VGND.n3057 VGND.n376 5.32359
R21173 VGND.n2986 VGND.n2970 5.32359
R21174 VGND.n2044 VGND.n567 5.32226
R21175 VGND.n2012 VGND.n573 5.32226
R21176 VGND.n1058 VGND.n1021 5.32226
R21177 VGND.n3347 VGND.n358 5.32226
R21178 VGND.n2124 VGND.t3600 5.32226
R21179 VGND.n2161 VGND.n2093 5.32226
R21180 VGND.n2069 VGND.n555 5.32226
R21181 VGND.t3414 VGND.n3465 5.32226
R21182 VGND.t2008 VGND.n3667 5.32226
R21183 VGND.t2646 VGND.n3638 5.32226
R21184 VGND.t2535 VGND.n3653 5.32226
R21185 VGND.t2267 VGND.n3479 5.32226
R21186 VGND.t2606 VGND.n3571 5.32226
R21187 VGND.t4826 VGND.n3603 5.32226
R21188 VGND.t2225 VGND.n3619 5.32226
R21189 VGND.t1659 VGND.n3587 5.32226
R21190 VGND.t6782 VGND.n3555 5.32226
R21191 VGND.t4363 VGND.n3543 5.32226
R21192 VGND.t4213 VGND.n20 5.32226
R21193 VGND.t4178 VGND.n35 5.32226
R21194 VGND.t3581 VGND.n3498 5.32226
R21195 VGND.t73 VGND.n3513 5.32226
R21196 VGND.t3779 VGND.n3528 5.32226
R21197 VGND.n3452 VGND.n55 5.32226
R21198 VGND.n3462 VGND.n55 5.32226
R21199 VGND.n110 VGND.n55 5.32226
R21200 VGND.n81 VGND.n55 5.32226
R21201 VGND.n63 VGND.n55 5.32226
R21202 VGND.n240 VGND.n55 5.32226
R21203 VGND.n213 VGND.n55 5.32226
R21204 VGND.n195 VGND.n55 5.32226
R21205 VGND.n166 VGND.n55 5.32226
R21206 VGND.n136 VGND.n55 5.32226
R21207 VGND.n3445 VGND.n55 5.32226
R21208 VGND.n1437 VGND.n55 5.32226
R21209 VGND.n1409 VGND.n55 5.32226
R21210 VGND.n881 VGND.n55 5.32226
R21211 VGND.n858 VGND.n55 5.32226
R21212 VGND.n833 VGND.n55 5.32226
R21213 VGND.n816 VGND.n55 5.32226
R21214 VGND.n929 VGND.n55 5.32226
R21215 VGND.n56 VGND.n55 5.32226
R21216 VGND.n356 VGND.n355 5.32226
R21217 VGND.n3698 VGND.n3697 5.32226
R21218 VGND.n53 VGND.n43 5.32226
R21219 VGND.n1381 VGND.n1370 5.32226
R21220 VGND.n1398 VGND.n1360 5.32226
R21221 VGND.n1574 VGND.n1354 5.32226
R21222 VGND.n1591 VGND.n1349 5.32226
R21223 VGND.n1336 VGND.n887 5.32226
R21224 VGND.n1318 VGND.n891 5.32226
R21225 VGND.n1303 VGND.n895 5.32226
R21226 VGND.n1289 VGND.n899 5.32226
R21227 VGND.n3428 VGND.n144 5.32226
R21228 VGND.n3418 VGND.n151 5.32226
R21229 VGND.n290 VGND.n289 5.32226
R21230 VGND.n333 VGND.n273 5.32226
R21231 VGND.n318 VGND.n278 5.32226
R21232 VGND.n303 VGND.n283 5.32226
R21233 VGND.n258 VGND.n250 5.32226
R21234 VGND.n3399 VGND.n200 5.32226
R21235 VGND.n1526 VGND.n1494 5.32226
R21236 VGND.n1554 VGND.n1484 5.32226
R21237 VGND.n1456 VGND.n1448 5.32226
R21238 VGND.n1625 VGND.n840 5.32226
R21239 VGND.n1273 VGND.n1245 5.32226
R21240 VGND.n3369 VGND.t2652 5.32226
R21241 VGND.n1755 VGND.n1725 5.32226
R21242 VGND.n1783 VGND.n1716 5.32226
R21243 VGND.n1694 VGND.n771 5.32226
R21244 VGND.n1671 VGND.n783 5.32226
R21245 VGND.n1639 VGND.n798 5.32226
R21246 VGND.n1231 VGND.n1202 5.32226
R21247 VGND.n1833 VGND.t3389 5.32226
R21248 VGND.n1870 VGND.t2954 5.32226
R21249 VGND.n1799 VGND.n726 5.32226
R21250 VGND.n745 VGND.n737 5.32226
R21251 VGND.n1964 VGND.n593 5.32226
R21252 VGND.n1143 VGND.t1151 5.32226
R21253 VGND VGND.n1122 5.32226
R21254 VGND.n629 VGND.n625 5.32226
R21255 VGND.n1993 VGND.n577 5.32226
R21256 VGND.n1104 VGND.n1076 5.32226
R21257 VGND.n676 VGND.t2257 5.32226
R21258 VGND.n713 VGND.t1923 5.32226
R21259 VGND.n1905 VGND.n665 5.32226
R21260 VGND.n1931 VGND.n655 5.32226
R21261 VGND VGND.t3888 5.32226
R21262 VGND.n2181 VGND.n2175 5.32226
R21263 VGND.n2407 VGND.n472 5.32226
R21264 VGND.n978 VGND.n943 5.32226
R21265 VGND.n1008 VGND.t5822 5.32226
R21266 VGND.n2589 VGND.t2824 5.32226
R21267 VGND.n2838 VGND.t3473 5.32226
R21268 VGND.n2872 VGND.t1491 5.32226
R21269 VGND VGND.t5938 5.32226
R21270 VGND VGND.t3370 5.32226
R21271 VGND VGND.t3491 5.32226
R21272 VGND.t3701 VGND 5.32226
R21273 VGND.n2742 VGND.t2323 5.32226
R21274 VGND.n2813 VGND.t1818 5.32226
R21275 VGND.n2776 VGND.t547 5.32226
R21276 VGND.n2718 VGND.n2630 5.32226
R21277 VGND.n2681 VGND.t3368 5.32226
R21278 VGND.n2644 VGND.n2633 5.32226
R21279 VGND.n541 VGND.t3243 5.32226
R21280 VGND.n2376 VGND.n522 5.32226
R21281 VGND.n491 VGND.t4170 5.32226
R21282 VGND.n2442 VGND.n467 5.32226
R21283 VGND.n440 VGND.t3241 5.32226
R21284 VGND.n2342 VGND.t4039 5.32226
R21285 VGND.n2303 VGND.t414 5.32226
R21286 VGND.n2266 VGND.t1396 5.32226
R21287 VGND.n2227 VGND.n2223 5.32226
R21288 VGND.n2482 VGND.t397 5.32226
R21289 VGND.n2552 VGND.n2492 5.32226
R21290 VGND.n2535 VGND.n2493 5.32226
R21291 VGND.n2514 VGND.n2495 5.32226
R21292 VGND.n2504 VGND.n2496 5.32226
R21293 VGND.n2891 VGND.n406 5.32226
R21294 VGND.n2908 VGND.n405 5.32226
R21295 VGND.n2951 VGND.n2950 5.32226
R21296 VGND.n2941 VGND.n2920 5.32226
R21297 VGND.n2931 VGND.n2921 5.32226
R21298 VGND.n18 VGND.n8 5.32226
R21299 VGND.n3735 VGND.n7 5.32226
R21300 VGND.n3753 VGND.n5 5.32226
R21301 VGND.n3322 VGND.n3313 5.32226
R21302 VGND.n3333 VGND.n3311 5.32226
R21303 VGND.n3310 VGND.n3309 5.32226
R21304 VGND.n3277 VGND.n362 5.32226
R21305 VGND.n3192 VGND.n3183 5.32226
R21306 VGND.n3204 VGND.n3181 5.32226
R21307 VGND.n3180 VGND.n3179 5.32226
R21308 VGND.n3150 VGND.n369 5.32226
R21309 VGND.n3085 VGND.n3077 5.32226
R21310 VGND.n3098 VGND.n3075 5.32226
R21311 VGND.n3074 VGND.n3073 5.32226
R21312 VGND.n3047 VGND.n377 5.32226
R21313 VGND.n2978 VGND.n2971 5.32226
R21314 VGND.n2992 VGND.n2969 5.32226
R21315 VGND.n3786 VGND.n3777 5.32226
R21316 VGND.n3776 VGND.n3775 5.32226
R21317 VGND.n3758 VGND.n1 5.32226
R21318 VGND.n3242 VGND.n3234 5.32226
R21319 VGND.n3251 VGND.n3233 5.32226
R21320 VGND.n3261 VGND.n3232 5.32226
R21321 VGND.n3270 VGND.n3231 5.32226
R21322 VGND.n3230 VGND.n3229 5.32226
R21323 VGND.n3214 VGND.n365 5.32226
R21324 VGND.n3132 VGND.n3126 5.32226
R21325 VGND.n3141 VGND.n3125 5.32226
R21326 VGND.n3124 VGND.n3123 5.32226
R21327 VGND.n3109 VGND.n372 5.32226
R21328 VGND.n3027 VGND.n3021 5.32226
R21329 VGND.n3036 VGND.n3020 5.32226
R21330 VGND.n3019 VGND.n3018 5.32226
R21331 VGND.n3005 VGND.n380 5.32226
R21332 VGND.n3274 VGND.n363 5.2925
R21333 VGND.n3337 VGND.n3336 5.2925
R21334 VGND.t146 VGND 5.15045
R21335 VGND.n892 VGND.t947 5.06876
R21336 VGND.n1450 VGND.t989 5.06876
R21337 VGND.n592 VGND.t1703 5.06876
R21338 VGND.n3409 VGND.n196 4.9415
R21339 VGND.n1280 VGND.n935 4.9415
R21340 VGND.n837 VGND.n836 4.9415
R21341 VGND.n1596 VGND.n885 4.9415
R21342 VGND.n1562 VGND.n1442 4.9415
R21343 VGND.n3433 VGND.n3432 4.9415
R21344 VGND.n244 VGND.n243 4.9415
R21345 VGND.n3685 VGND.n3463 4.9415
R21346 VGND.n80 VGND.n3 4.9415
R21347 VGND.t5778 VGND.t3800 4.61698
R21348 VGND.t6434 VGND.t642 4.61698
R21349 VGND.t3469 VGND.t3216 4.61698
R21350 VGND.t3418 VGND.t3214 4.61698
R21351 VGND.t2058 VGND.t6551 4.61698
R21352 VGND.n557 VGND.t5256 4.5505
R21353 VGND.n557 VGND.t4894 4.5505
R21354 VGND.n556 VGND.t2381 4.5505
R21355 VGND.n556 VGND.t6638 4.5505
R21356 VGND.n910 VGND.t6512 4.5505
R21357 VGND.n910 VGND.t3175 4.5505
R21358 VGND.n804 VGND.t46 4.5505
R21359 VGND.n804 VGND.t1361 4.5505
R21360 VGND.n825 VGND.t3084 4.5505
R21361 VGND.n825 VGND.t6735 4.5505
R21362 VGND.n846 VGND.t5272 4.5505
R21363 VGND.n846 VGND.t176 4.5505
R21364 VGND.n869 VGND.t81 4.5505
R21365 VGND.n1424 VGND.t4519 4.5505
R21366 VGND.n1427 VGND.t5707 4.5505
R21367 VGND.n897 VGND.t6566 4.5505
R21368 VGND.n1352 VGND.t3803 4.5505
R21369 VGND.n1352 VGND.t4069 4.5505
R21370 VGND.n1350 VGND.t3801 4.5505
R21371 VGND.n1350 VGND.t1014 4.5505
R21372 VGND.n1446 VGND.t3675 4.5505
R21373 VGND.n1446 VGND.t4539 4.5505
R21374 VGND.n1492 VGND.t2242 4.5505
R21375 VGND.n722 VGND.t170 4.5505
R21376 VGND.n734 VGND.t6552 4.5505
R21377 VGND.n734 VGND.t951 4.5505
R21378 VGND.n735 VGND.t3769 4.5505
R21379 VGND.n735 VGND.t5511 4.5505
R21380 VGND.n610 VGND.t4838 4.5505
R21381 VGND.n610 VGND.t4840 4.5505
R21382 VGND.n608 VGND.t2416 4.5505
R21383 VGND.n608 VGND.t1699 4.5505
R21384 VGND.n600 VGND.t122 4.5505
R21385 VGND.n600 VGND.t6718 4.5505
R21386 VGND.n586 VGND.t6334 4.5505
R21387 VGND.n586 VGND.t180 4.5505
R21388 VGND.n657 VGND.t3772 4.5505
R21389 VGND.n657 VGND.t6643 4.5505
R21390 VGND.n2172 VGND.t6159 4.5505
R21391 VGND.n3410 VGND.n3409 4.5005
R21392 VGND.n3408 VGND.n3407 4.5005
R21393 VGND.n1762 VGND.n197 4.5005
R21394 VGND.n1876 VGND.n1875 4.5005
R21395 VGND.n1878 VGND.n1877 4.5005
R21396 VGND.n1113 VGND.n1112 4.5005
R21397 VGND.n1014 VGND.n1013 4.5005
R21398 VGND.n2600 VGND.n2599 4.5005
R21399 VGND.n2622 VGND.n2621 4.5005
R21400 VGND.n2611 VGND.n2610 4.5005
R21401 VGND.n393 VGND.n384 4.5005
R21402 VGND.n2962 VGND.n2961 4.5005
R21403 VGND.n1191 VGND.n1190 4.5005
R21404 VGND.n1239 VGND.n1238 4.5005
R21405 VGND.n1279 VGND.n1278 4.5005
R21406 VGND.n1281 VGND.n1280 4.5005
R21407 VGND.n2732 VGND.n2731 4.5005
R21408 VGND.n2825 VGND.n2824 4.5005
R21409 VGND.n2827 VGND.n2826 4.5005
R21410 VGND.n982 VGND.n427 4.5005
R21411 VGND.n2002 VGND.n2001 4.5005
R21412 VGND.n1151 VGND.n575 4.5005
R21413 VGND.n1632 VGND.n1631 4.5005
R21414 VGND.n1630 VGND.n1629 4.5005
R21415 VGND.n1313 VGND.n837 4.5005
R21416 VGND.n2692 VGND.n378 4.5005
R21417 VGND.n2730 VGND.n2729 4.5005
R21418 VGND.n2655 VGND.n374 4.5005
R21419 VGND.n2787 VGND.n408 4.5005
R21420 VGND.n2884 VGND.n2883 4.5005
R21421 VGND.n2411 VGND.n2410 4.5005
R21422 VGND.n1972 VGND.n1971 4.5005
R21423 VGND.n1970 VGND.n1969 4.5005
R21424 VGND.n1665 VGND.n588 4.5005
R21425 VGND.n1598 VGND.n1597 4.5005
R21426 VGND.n1596 VGND.n1595 4.5005
R21427 VGND.n2413 VGND.n2412 4.5005
R21428 VGND.n2447 VGND.n2446 4.5005
R21429 VGND.n435 VGND.n419 4.5005
R21430 VGND.n2382 VGND.n2381 4.5005
R21431 VGND.n2384 VGND.n2383 4.5005
R21432 VGND.n1938 VGND.n1937 4.5005
R21433 VGND.n1940 VGND.n1939 4.5005
R21434 VGND.n1689 VGND.n612 4.5005
R21435 VGND.n1561 VGND.n1560 4.5005
R21436 VGND.n1563 VGND.n1562 4.5005
R21437 VGND.n2297 VGND.n484 4.5005
R21438 VGND.n2261 VGND.n407 4.5005
R21439 VGND.n2449 VGND.n2448 4.5005
R21440 VGND.n2488 VGND.n2487 4.5005
R21441 VGND.n2350 VGND.n2349 4.5005
R21442 VGND.n2352 VGND.n2351 4.5005
R21443 VGND.n2221 VGND.n2220 4.5005
R21444 VGND.n1912 VGND.n548 4.5005
R21445 VGND.n1794 VGND.n1793 4.5005
R21446 VGND.n1792 VGND.n1791 4.5005
R21447 VGND.n1532 VGND.n141 4.5005
R21448 VGND.n3432 VGND.n3431 4.5005
R21449 VGND.n2935 VGND.n367 4.5005
R21450 VGND.n2916 VGND.n370 4.5005
R21451 VGND.n2886 VGND.n2885 4.5005
R21452 VGND.n2524 VGND.n411 4.5005
R21453 VGND.n2558 VGND.n2557 4.5005
R21454 VGND.n2132 VGND.n363 4.5005
R21455 VGND.n2168 VGND.n2167 4.5005
R21456 VGND.n2066 VGND.n483 4.5005
R21457 VGND.n2040 VGND.n469 4.5005
R21458 VGND.n2004 VGND.n2003 4.5005
R21459 VGND.n1067 VGND.n1066 4.5005
R21460 VGND.n3338 VGND.n3337 4.5005
R21461 VGND.n685 VGND.n359 4.5005
R21462 VGND.n1842 VGND.n245 4.5005
R21463 VGND.n3378 VGND.n3377 4.5005
R21464 VGND.n3380 VGND.n3379 4.5005
R21465 VGND.n315 VGND.n244 4.5005
R21466 VGND.n3336 VGND.n3335 4.5005
R21467 VGND.n3275 VGND.n3274 4.5005
R21468 VGND.n3209 VGND.n3208 4.5005
R21469 VGND.n3147 VGND.n3146 4.5005
R21470 VGND.n3104 VGND.n3103 4.5005
R21471 VGND.n3043 VGND.n3042 4.5005
R21472 VGND.n2999 VGND.n2998 4.5005
R21473 VGND.n3718 VGND.n3717 4.5005
R21474 VGND.n3715 VGND.n3714 4.5005
R21475 VGND.n34 VGND.n19 4.5005
R21476 VGND.n3509 VGND.n3508 4.5005
R21477 VGND.n3524 VGND.n3523 4.5005
R21478 VGND.n3539 VGND.n3538 4.5005
R21479 VGND.n3554 VGND.n3553 4.5005
R21480 VGND.n3570 VGND.n3569 4.5005
R21481 VGND.n3586 VGND.n3585 4.5005
R21482 VGND.n3602 VGND.n3601 4.5005
R21483 VGND.n3618 VGND.n3617 4.5005
R21484 VGND.n3634 VGND.n3633 4.5005
R21485 VGND.n3649 VGND.n3648 4.5005
R21486 VGND.n3664 VGND.n3663 4.5005
R21487 VGND.n3666 VGND.n3665 4.5005
R21488 VGND.n3478 VGND.n3464 4.5005
R21489 VGND.n3684 VGND.n3683 4.5005
R21490 VGND.n3686 VGND.n3685 4.5005
R21491 VGND.n3716 VGND.n0 4.5005
R21492 VGND.n3253 VGND.n360 4.5005
R21493 VGND.n3273 VGND.n3272 4.5005
R21494 VGND.n3211 VGND.n3210 4.5005
R21495 VGND.n3145 VGND.n3144 4.5005
R21496 VGND.n3106 VGND.n3105 4.5005
R21497 VGND.n3041 VGND.n3040 4.5005
R21498 VGND.n3001 VGND.n3000 4.5005
R21499 VGND.n3757 VGND.n3756 4.5005
R21500 VGND.n3755 VGND.n3754 4.5005
R21501 VGND.n346 VGND.n3 4.5005
R21502 VGND.n909 VGND.t3176 4.48817
R21503 VGND.n802 VGND.t349 4.48817
R21504 VGND.n800 VGND.t5329 4.48817
R21505 VGND.n847 VGND.t5728 4.48817
R21506 VGND.n739 VGND.t3468 4.30241
R21507 VGND.n623 VGND.t1403 4.30241
R21508 VGND VGND.t45 4.14907
R21509 VGND.n2086 VGND.t3893 4.0955
R21510 VGND.n564 VGND.t2930 4.0955
R21511 VGND.n180 VGND.t5061 4.0955
R21512 VGND.n161 VGND.t2177 4.0955
R21513 VGND.n1401 VGND.t2053 4.0955
R21514 VGND.n871 VGND.t4896 4.0955
R21515 VGND.n893 VGND.t2133 4.0955
R21516 VGND.n893 VGND.t874 4.0955
R21517 VGND.n892 VGND.t6009 4.0955
R21518 VGND.n1356 VGND.t5293 4.0955
R21519 VGND.n1372 VGND.t665 4.0955
R21520 VGND.n146 VGND.t3376 4.0955
R21521 VGND.n153 VGND.t4898 4.0955
R21522 VGND.n1358 VGND.t1573 4.0955
R21523 VGND.n1488 VGND.t985 4.0955
R21524 VGND.n199 VGND.t3510 4.0955
R21525 VGND.n1485 VGND.t5280 4.0955
R21526 VGND.n1473 VGND.t2821 4.0955
R21527 VGND.n1449 VGND.t6427 4.0955
R21528 VGND.n1449 VGND.t3689 4.0955
R21529 VGND.n1450 VGND.t4529 4.0955
R21530 VGND.n203 VGND.t2393 4.0955
R21531 VGND.n789 VGND.t2154 4.0955
R21532 VGND.n774 VGND.t3955 4.0955
R21533 VGND.n1730 VGND.t5616 4.0955
R21534 VGND.n1726 VGND.t3924 4.0955
R21535 VGND.n1722 VGND.t455 4.0955
R21536 VGND.n768 VGND.t5693 4.0955
R21537 VGND.n591 VGND.t3158 4.0955
R21538 VGND.n591 VGND.t6664 4.0955
R21539 VGND.n592 VGND.t124 4.0955
R21540 VGND.n731 VGND.t1590 4.0955
R21541 VGND.n724 VGND.t3003 4.0955
R21542 VGND.n728 VGND.t683 4.0955
R21543 VGND.n584 VGND.t2179 4.0955
R21544 VGND.n663 VGND.t2137 4.0955
R21545 VGND.n581 VGND.t859 4.0955
R21546 VGND.n949 VGND.t2603 4.0955
R21547 VGND.n475 VGND.t2338 4.0955
R21548 VGND.n2194 VGND.t1265 4.0955
R21549 VGND.n2176 VGND.t328 4.0955
R21550 VGND.n473 VGND.t5245 4.0955
R21551 VGND.n508 VGND.t3047 4.0955
R21552 VGND.n527 VGND.t1705 4.0955
R21553 VGND.n526 VGND.t1378 4.0955
R21554 VGND.n2094 VGND.t41 4.04494
R21555 VGND.n2094 VGND.t6364 4.04494
R21556 VGND.n561 VGND.t192 4.04494
R21557 VGND.n561 VGND.t6362 4.04494
R21558 VGND.n228 VGND.t140 4.04494
R21559 VGND.n228 VGND.t6195 4.04494
R21560 VGND.n182 VGND.t156 4.04494
R21561 VGND.n182 VGND.t6196 4.04494
R21562 VGND.n159 VGND.t6095 4.04494
R21563 VGND.n159 VGND.t6199 4.04494
R21564 VGND.n1421 VGND.t6410 4.04494
R21565 VGND.n1421 VGND.t6412 4.04494
R21566 VGND.n1403 VGND.t6459 4.04494
R21567 VGND.n1403 VGND.t6742 4.04494
R21568 VGND.n868 VGND.t6455 4.04494
R21569 VGND.n868 VGND.t6633 4.04494
R21570 VGND.n1359 VGND.t6729 4.04494
R21571 VGND.n1359 VGND.t6205 4.04494
R21572 VGND.n142 VGND.t6741 4.04494
R21573 VGND.n142 VGND.t6211 4.04494
R21574 VGND.n150 VGND.t88 4.04494
R21575 VGND.n150 VGND.t6215 4.04494
R21576 VGND.n156 VGND.t6557 4.04494
R21577 VGND.n156 VGND.t6219 4.04494
R21578 VGND.n274 VGND.t6595 4.04494
R21579 VGND.n274 VGND.t6213 4.04494
R21580 VGND.n1363 VGND.t6779 4.04494
R21581 VGND.n1363 VGND.t6221 4.04494
R21582 VGND.n1491 VGND.t6328 4.04494
R21583 VGND.n1491 VGND.t6354 4.04494
R21584 VGND.n207 VGND.t101 4.04494
R21585 VGND.n207 VGND.t6207 4.04494
R21586 VGND.n247 VGND.t6114 4.04494
R21587 VGND.n247 VGND.t6217 4.04494
R21588 VGND.n202 VGND.t6070 4.04494
R21589 VGND.n202 VGND.t6201 4.04494
R21590 VGND.n1487 VGND.t226 4.04494
R21591 VGND.n1487 VGND.t6356 4.04494
R21592 VGND.n1444 VGND.t145 4.04494
R21593 VGND.n1444 VGND.t6374 4.04494
R21594 VGND.n795 VGND.t6461 4.04494
R21595 VGND.n795 VGND.t6097 4.04494
R21596 VGND.n777 VGND.t6447 4.04494
R21597 VGND.n777 VGND.t174 4.04494
R21598 VGND.n1724 VGND.t6476 4.04494
R21599 VGND.n1724 VGND.t6209 4.04494
R21600 VGND.n1733 VGND.t6684 4.04494
R21601 VGND.n1733 VGND.t6194 4.04494
R21602 VGND.n1729 VGND.t6707 4.04494
R21603 VGND.n1729 VGND.t6203 4.04494
R21604 VGND.n1718 VGND.t33 4.04494
R21605 VGND.n1718 VGND.t6198 4.04494
R21606 VGND.n780 VGND.t251 4.04494
R21607 VGND.n780 VGND.t267 4.04494
R21608 VGND.n781 VGND.t257 4.04494
R21609 VGND.n781 VGND.t255 4.04494
R21610 VGND.n782 VGND.t265 4.04494
R21611 VGND.n782 VGND.t253 4.04494
R21612 VGND.n595 VGND.t6529 4.04494
R21613 VGND.n595 VGND.t6533 4.04494
R21614 VGND.n597 VGND.t6531 4.04494
R21615 VGND.n597 VGND.t6527 4.04494
R21616 VGND.n598 VGND.t6525 4.04494
R21617 VGND.n598 VGND.t6523 4.04494
R21618 VGND.n729 VGND.t6133 4.04494
R21619 VGND.n729 VGND.t6360 4.04494
R21620 VGND.n1813 VGND.t6116 4.04494
R21621 VGND.n1813 VGND.t6223 4.04494
R21622 VGND.n725 VGND.t152 4.04494
R21623 VGND.n725 VGND.t6380 4.04494
R21624 VGND.n579 VGND.t6457 4.04494
R21625 VGND.n579 VGND.t22 4.04494
R21626 VGND.n621 VGND.t261 4.04494
R21627 VGND.n621 VGND.t259 4.04494
R21628 VGND.n620 VGND.t263 4.04494
R21629 VGND.n620 VGND.t249 4.04494
R21630 VGND.n619 VGND.t245 4.04494
R21631 VGND.n619 VGND.t247 4.04494
R21632 VGND.n666 VGND.t93 4.04494
R21633 VGND.n666 VGND.t6366 4.04494
R21634 VGND.n578 VGND.t6451 4.04494
R21635 VGND.n578 VGND.t6310 4.04494
R21636 VGND.n945 VGND.t6453 4.04494
R21637 VGND.n945 VGND.t6147 4.04494
R21638 VGND.n479 VGND.t6712 4.04494
R21639 VGND.n479 VGND.t6358 4.04494
R21640 VGND.n2171 VGND.t86 4.04494
R21641 VGND.n2171 VGND.t6372 4.04494
R21642 VGND.n480 VGND.t6376 4.04494
R21643 VGND.n480 VGND.t6190 4.04494
R21644 VGND.n948 VGND.t6449 4.04494
R21645 VGND.n948 VGND.t127 4.04494
R21646 VGND.n487 VGND.t6734 4.04494
R21647 VGND.n487 VGND.t6370 4.04494
R21648 VGND.n530 VGND.t6632 4.04494
R21649 VGND.n530 VGND.t6378 4.04494
R21650 VGND.n486 VGND.t6368 4.04494
R21651 VGND.n486 VGND.t161 4.04494
R21652 VGND.n1425 VGND.t6406 3.8098
R21653 VGND.n1425 VGND.t6404 3.8098
R21654 VGND.n1423 VGND.t6401 3.8098
R21655 VGND.n1423 VGND.t6407 3.8098
R21656 VGND.n1422 VGND.t6408 3.8098
R21657 VGND.n1422 VGND.t6402 3.8098
R21658 VGND.n1424 VGND.t5968 3.77367
R21659 VGND.n897 VGND.t3266 3.77367
R21660 VGND.n1492 VGND.t1986 3.77367
R21661 VGND.n722 VGND.t5507 3.77367
R21662 VGND.n2172 VGND.t1934 3.77367
R21663 VGND.n919 VGND.t5881 3.6005
R21664 VGND.n919 VGND.t5883 3.6005
R21665 VGND.n850 VGND.t4515 3.6005
R21666 VGND.n850 VGND.t4516 3.6005
R21667 VGND.n113 VGND.t4814 3.6005
R21668 VGND.n113 VGND.t4815 3.6005
R21669 VGND.n918 VGND.t1062 3.6005
R21670 VGND.n918 VGND.t1060 3.6005
R21671 VGND.n1362 VGND.t4027 3.6005
R21672 VGND.n1362 VGND.t4031 3.6005
R21673 VGND.n1447 VGND.t2864 3.6005
R21674 VGND.n1447 VGND.t2870 3.6005
R21675 VGND.n3146 VGND.n370 3.5285
R21676 VGND.n3209 VGND.n367 3.5285
R21677 VGND.n563 VGND.t3042 3.52308
R21678 VGND.n563 VGND.t203 3.52308
R21679 VGND.n552 VGND.t2454 3.52308
R21680 VGND.n552 VGND.t207 3.52308
R21681 VGND.n123 VGND.t5564 3.52308
R21682 VGND.n123 VGND.t6471 3.52308
R21683 VGND.n1339 VGND.t6745 3.52308
R21684 VGND.n1339 VGND.t6444 3.52308
R21685 VGND.n1351 VGND.t2545 3.52308
R21686 VGND.n1351 VGND.t4152 3.52308
R21687 VGND.n284 VGND.t6395 3.52308
R21688 VGND.n284 VGND.t1101 3.52308
R21689 VGND.n154 VGND.t5524 3.52308
R21690 VGND.n154 VGND.t6469 3.52308
R21691 VGND.n1353 VGND.t5132 3.52308
R21692 VGND.n1353 VGND.t1425 3.52308
R21693 VGND.n896 VGND.t2383 3.52308
R21694 VGND.n896 VGND.t4906 3.52308
R21695 VGND.n1502 VGND.t6230 3.52308
R21696 VGND.n1502 VGND.t3427 3.52308
R21697 VGND.n205 VGND.t3071 3.52308
R21698 VGND.n205 VGND.t6397 3.52308
R21699 VGND.n1206 VGND.t1115 3.52308
R21700 VGND.n1206 VGND.t770 3.52308
R21701 VGND.n1727 VGND.t3105 3.52308
R21702 VGND.n1727 VGND.t6388 3.52308
R21703 VGND.n1720 VGND.t4689 3.52308
R21704 VGND.n1720 VGND.t6390 3.52308
R21705 VGND.n769 VGND.t6107 3.52308
R21706 VGND.n769 VGND.t201 3.52308
R21707 VGND.n770 VGND.t570 3.52308
R21708 VGND.n770 VGND.t205 3.52308
R21709 VGND.n736 VGND.t5400 3.52308
R21710 VGND.n736 VGND.t5644 3.52308
R21711 VGND.n1815 VGND.t2858 3.52308
R21712 VGND.n1815 VGND.t6384 3.52308
R21713 VGND.n656 VGND.t2261 3.52308
R21714 VGND.n656 VGND.t3248 3.52308
R21715 VGND.n660 VGND.t220 3.52308
R21716 VGND.n660 VGND.t4326 3.52308
R21717 VGND.n624 VGND.t4993 3.52308
R21718 VGND.n624 VGND.t916 3.52308
R21719 VGND.n2174 VGND.t224 3.52308
R21720 VGND.n2174 VGND.t5466 3.52308
R21721 VGND.n2196 VGND.t6124 3.52308
R21722 VGND.n2196 VGND.t211 3.52308
R21723 VGND.n2170 VGND.t1127 3.52308
R21724 VGND.n2170 VGND.t222 3.52308
R21725 VGND.n476 VGND.t6026 3.52308
R21726 VGND.n476 VGND.t198 3.52308
R21727 VGND.n523 VGND.t217 3.52308
R21728 VGND.n523 VGND.t3584 3.52308
R21729 VGND.n1364 VGND.t3447 3.45782
R21730 VGND.n784 VGND.t6277 3.37782
R21731 VGND.n784 VGND.t6272 3.37782
R21732 VGND.n786 VGND.t6278 3.37782
R21733 VGND.n786 VGND.t6273 3.37782
R21734 VGND.n787 VGND.t6286 3.37782
R21735 VGND.n787 VGND.t6284 3.37782
R21736 VGND.n788 VGND.t6288 3.37782
R21737 VGND.n788 VGND.t6290 3.37782
R21738 VGND.n790 VGND.t6262 3.37782
R21739 VGND.n790 VGND.t6264 3.37782
R21740 VGND.n791 VGND.t6270 3.37782
R21741 VGND.n791 VGND.t6266 3.37782
R21742 VGND.n793 VGND.t6282 3.37782
R21743 VGND.n793 VGND.t6280 3.37782
R21744 VGND.n601 VGND.t291 3.37782
R21745 VGND.n601 VGND.t295 3.37782
R21746 VGND.n602 VGND.t283 3.37782
R21747 VGND.n602 VGND.t279 3.37782
R21748 VGND.n603 VGND.t281 3.37782
R21749 VGND.n603 VGND.t277 3.37782
R21750 VGND.n604 VGND.t273 3.37782
R21751 VGND.n604 VGND.t271 3.37782
R21752 VGND.n606 VGND.t243 3.37782
R21753 VGND.n606 VGND.t269 3.37782
R21754 VGND.n607 VGND.t287 3.37782
R21755 VGND.n607 VGND.t293 3.37782
R21756 VGND.n609 VGND.t289 3.37782
R21757 VGND.n609 VGND.t285 3.37782
R21758 VGND.n645 VGND.t6621 3.37782
R21759 VGND.n645 VGND.t6617 3.37782
R21760 VGND.n646 VGND.t6601 3.37782
R21761 VGND.n646 VGND.t6607 3.37782
R21762 VGND.n647 VGND.t6603 3.37782
R21763 VGND.n647 VGND.t6605 3.37782
R21764 VGND.n648 VGND.t6627 3.37782
R21765 VGND.n648 VGND.t6625 3.37782
R21766 VGND.n613 VGND.t6597 3.37782
R21767 VGND.n613 VGND.t6623 3.37782
R21768 VGND.n616 VGND.t6615 3.37782
R21769 VGND.n616 VGND.t6611 3.37782
R21770 VGND.n617 VGND.t6609 3.37782
R21771 VGND.n617 VGND.t6613 3.37782
R21772 VGND.n1501 VGND.t3431 3.21226
R21773 VGND.n1501 VGND.t3425 3.21226
R21774 VGND.n594 VGND.t3150 3.18108
R21775 VGND.n594 VGND.t3152 3.18108
R21776 VGND.n210 VGND.t4868 2.93792
R21777 VGND.n279 VGND.t5795 2.93792
R21778 VGND.n251 VGND.t388 2.93792
R21779 VGND.n1426 VGND.t6249 2.89962
R21780 VGND.n1426 VGND.t6246 2.89962
R21781 VGND.n1428 VGND.t3514 2.89962
R21782 VGND.n1428 VGND.t3515 2.89962
R21783 VGND.n112 VGND.t6243 2.89962
R21784 VGND.n112 VGND.t6239 2.89962
R21785 VGND.n114 VGND.t6481 2.89962
R21786 VGND.n114 VGND.t6479 2.89962
R21787 VGND.n115 VGND.t6066 2.89962
R21788 VGND.n115 VGND.t6065 2.89962
R21789 VGND.n119 VGND.t6485 2.89962
R21790 VGND.n119 VGND.t6483 2.89962
R21791 VGND.n121 VGND.t1140 2.89962
R21792 VGND.n121 VGND.t1141 2.89962
R21793 VGND.n122 VGND.t6482 2.89962
R21794 VGND.n122 VGND.t6480 2.89962
R21795 VGND.n120 VGND.t6484 2.89962
R21796 VGND.n120 VGND.t6490 2.89962
R21797 VGND.n118 VGND.t149 2.89962
R21798 VGND.n118 VGND.t148 2.89962
R21799 VGND.n117 VGND.t6496 2.89962
R21800 VGND.n117 VGND.t6495 2.89962
R21801 VGND.n116 VGND.t6494 2.89962
R21802 VGND.n116 VGND.t6491 2.89962
R21803 VGND.n1365 VGND.t6238 2.89962
R21804 VGND.n1365 VGND.t6248 2.89962
R21805 VGND.n1367 VGND.t5701 2.89962
R21806 VGND.n1367 VGND.t5703 2.89962
R21807 VGND.n1368 VGND.t6245 2.89962
R21808 VGND.n1368 VGND.t6241 2.89962
R21809 VGND.n1495 VGND.t6478 2.89962
R21810 VGND.n1495 VGND.t6493 2.89962
R21811 VGND.n1496 VGND.t1932 2.89962
R21812 VGND.n1496 VGND.t1928 2.89962
R21813 VGND.n1497 VGND.t6487 2.89962
R21814 VGND.n1497 VGND.t6489 2.89962
R21815 VGND.n739 VGND.t2332 2.89962
R21816 VGND.n623 VGND.t6419 2.89962
R21817 VGND.n158 VGND.t6465 2.72794
R21818 VGND.n158 VGND.t867 2.72794
R21819 VGND.n1445 VGND.t188 2.72794
R21820 VGND.n1445 VGND.t1537 2.72794
R21821 VGND.n3673 VGND 2.66571
R21822 VGND.n3668 VGND 2.66571
R21823 VGND VGND.n3482 2.66571
R21824 VGND VGND.n3481 2.66571
R21825 VGND.n3480 VGND 2.66571
R21826 VGND.n3575 VGND 2.66571
R21827 VGND.n3607 VGND 2.66571
R21828 VGND.n3623 VGND 2.66571
R21829 VGND.n3591 VGND 2.66571
R21830 VGND.n3559 VGND 2.66571
R21831 VGND VGND.n40 2.66571
R21832 VGND.n3704 VGND 2.66571
R21833 VGND.n36 VGND 2.66571
R21834 VGND VGND.n37 2.66571
R21835 VGND VGND.n21 2.66571
R21836 VGND VGND.n38 2.66571
R21837 VGND VGND.n403 2.66571
R21838 VGND VGND.n401 2.66571
R21839 VGND VGND.n402 2.66571
R21840 VGND.n3357 VGND 2.66471
R21841 VGND.n270 VGND 2.66471
R21842 VGND VGND.n3359 2.66471
R21843 VGND VGND.n271 2.66471
R21844 VGND VGND.n272 2.66471
R21845 VGND VGND.n2207 2.66471
R21846 VGND VGND.n388 2.66471
R21847 VGND VGND.n389 2.66471
R21848 VGND.n400 VGND 2.66471
R21849 VGND VGND.n2954 2.66471
R21850 VGND VGND.n531 2.66471
R21851 VGND VGND.n2332 2.66471
R21852 VGND.n566 VGND.t6781 2.52151
R21853 VGND.n848 VGND.t5382 2.52151
R21854 VGND.n738 VGND.t5428 2.52151
R21855 VGND.n658 VGND.t5606 2.52151
R21856 VGND.n596 VGND.t872 2.34987
R21857 VGND.n1500 VGND.t6294 2.27826
R21858 VGND.n3042 VGND.n378 2.2055
R21859 VGND.n3104 VGND.n374 2.2055
R21860 VGND.n801 VGND.t3 2.11405
R21861 VGND.n1493 VGND.t3027 2.11405
R21862 VGND.n1719 VGND.t1039 2.11405
R21863 VGND.n661 VGND.t2272 2.11405
R21864 VGND.n2173 VGND.t5782 2.11405
R21865 VGND.n525 VGND.t878 2.11405
R21866 VGND.n553 VGND.t4982 2.01032
R21867 VGND.n549 VGND.t3789 2.01032
R21868 VGND.n210 VGND.t1853 2.01032
R21869 VGND.n211 VGND.t4867 2.01032
R21870 VGND.n211 VGND.t4865 2.01032
R21871 VGND.n209 VGND.t1854 2.01032
R21872 VGND.n286 VGND.t4910 2.01032
R21873 VGND.n277 VGND.t3522 2.01032
R21874 VGND.n279 VGND.t3520 2.01032
R21875 VGND.n280 VGND.t5789 2.01032
R21876 VGND.n280 VGND.t5797 2.01032
R21877 VGND.n285 VGND.t2121 2.01032
R21878 VGND.n249 VGND.t1271 2.01032
R21879 VGND.n251 VGND.t1269 2.01032
R21880 VGND.n252 VGND.t390 2.01032
R21881 VGND.n252 VGND.t392 2.01032
R21882 VGND.n844 VGND.t3973 2.01032
R21883 VGND.n733 VGND.t1966 2.01032
R21884 VGND.n1814 VGND.t3699 2.01032
R21885 VGND.n1125 VGND.t5218 2.01032
R21886 VGND.n662 VGND.t3065 2.01032
R21887 VGND.n2195 VGND.t1907 2.01032
R21888 VGND.n571 VGND.t3813 1.99806
R21889 VGND.n571 VGND.t3786 1.99806
R21890 VGND.n568 VGND.t6332 1.99806
R21891 VGND.n568 VGND.t5216 1.99806
R21892 VGND.n558 VGND.t4541 1.99806
R21893 VGND.n558 VGND.t4521 1.99806
R21894 VGND.n569 VGND.t461 1.99806
R21895 VGND.n807 VGND.t2404 1.99806
R21896 VGND.n806 VGND.t5456 1.99806
R21897 VGND.n212 VGND.t1291 1.99806
R21898 VGND.n849 VGND.t4455 1.99806
R21899 VGND.n849 VGND.t4454 1.99806
R21900 VGND.n803 VGND.t4967 1.99806
R21901 VGND.n805 VGND.t5824 1.99806
R21902 VGND.n890 VGND.t2519 1.99806
R21903 VGND.n890 VGND.t2523 1.99806
R21904 VGND.n889 VGND.t6013 1.99806
R21905 VGND.n889 VGND.t6011 1.99806
R21906 VGND.n1338 VGND.t5674 1.99806
R21907 VGND.n1338 VGND.t2521 1.99806
R21908 VGND.n281 VGND.t5809 1.99806
R21909 VGND.n276 VGND.t4232 1.99806
R21910 VGND.n287 VGND.t2433 1.99806
R21911 VGND.n287 VGND.t2438 1.99806
R21912 VGND.n288 VGND.t2431 1.99806
R21913 VGND.n288 VGND.t2435 1.99806
R21914 VGND.n149 VGND.t779 1.99806
R21915 VGND.n149 VGND.t775 1.99806
R21916 VGND.n147 VGND.t777 1.99806
R21917 VGND.n147 VGND.t781 1.99806
R21918 VGND.n145 VGND.t6656 1.99806
R21919 VGND.n145 VGND.t6658 1.99806
R21920 VGND.n143 VGND.t6660 1.99806
R21921 VGND.n143 VGND.t6654 1.99806
R21922 VGND.n1369 VGND.t3895 1.99806
R21923 VGND.n1366 VGND.t2984 1.99806
R21924 VGND.n1366 VGND.t2982 1.99806
R21925 VGND.n1364 VGND.t2980 1.99806
R21926 VGND.n888 VGND.t5049 1.99806
R21927 VGND.n888 VGND.t5045 1.99806
R21928 VGND.n839 VGND.t5289 1.99806
R21929 VGND.n839 VGND.t2385 1.99806
R21930 VGND.n843 VGND.t1347 1.99806
R21931 VGND.n843 VGND.t1351 1.99806
R21932 VGND.n1451 VGND.t1863 1.99806
R21933 VGND.n1451 VGND.t6330 1.99806
R21934 VGND.n1498 VGND.t6299 1.99806
R21935 VGND.n1498 VGND.t6296 1.99806
R21936 VGND.n842 VGND.t3737 1.99806
R21937 VGND.n842 VGND.t6694 1.99806
R21938 VGND.n841 VGND.t5532 1.99806
R21939 VGND.n841 VGND.t4687 1.99806
R21940 VGND.n1246 VGND.t5828 1.99806
R21941 VGND.n1246 VGND.t5055 1.99806
R21942 VGND.n797 VGND.t332 1.99806
R21943 VGND.n797 VGND.t1511 1.99806
R21944 VGND.n785 VGND.t2354 1.99806
R21945 VGND.n779 VGND.t760 1.99806
R21946 VGND.n779 VGND.t758 1.99806
R21947 VGND.n772 VGND.t2418 1.99806
R21948 VGND.n772 VGND.t2414 1.99806
R21949 VGND.n773 VGND.t2412 1.99806
R21950 VGND.n773 VGND.t2420 1.99806
R21951 VGND.n778 VGND.t2665 1.99806
R21952 VGND.n1207 VGND.t4003 1.99806
R21953 VGND.n1207 VGND.t6704 1.99806
R21954 VGND.n1205 VGND.t2593 1.99806
R21955 VGND.n1205 VGND.t1506 1.99806
R21956 VGND.n1204 VGND.t5230 1.99806
R21957 VGND.n1204 VGND.t2468 1.99806
R21958 VGND.n1203 VGND.t6702 1.99806
R21959 VGND.n1203 VGND.t1771 1.99806
R21960 VGND.n796 VGND.t4284 1.99806
R21961 VGND.n796 VGND.t6690 1.99806
R21962 VGND.n589 VGND.t6335 1.99806
R21963 VGND.n589 VGND.t5725 1.99806
R21964 VGND.n599 VGND.t832 1.99806
R21965 VGND.n585 VGND.t430 1.99806
R21966 VGND.n618 VGND.t239 1.99806
R21967 VGND.n618 VGND.t241 1.99806
R21968 VGND.n615 VGND.t235 1.99806
R21969 VGND.n615 VGND.t237 1.99806
R21970 VGND.n622 VGND.t1113 1.99806
R21971 VGND.n474 VGND.t3456 1.99806
R21972 VGND.n947 VGND.t6337 1.99806
R21973 VGND.n947 VGND.t2511 1.99806
R21974 VGND.n826 VGND.t5672 1.61041
R21975 VGND.n898 VGND.t1465 1.61041
R21976 VGND.t4150 VGND.t80 0.954194
R21977 VGND.t2 VGND.t1077 0.858825
R21978 VGND.t1059 VGND.t6400 0.763456
R21979 VGND.t45 VGND.t6793 0.715771
R21980 VGND.n1375 VGND.n1374 0.6965
R21981 VGND.n1686 VGND.n1685 0.6965
R21982 VGND VGND.n1375 0.6485
R21983 VGND.t3209 VGND.t4 0.572717
R21984 VGND.t6 VGND.t4514 0.572717
R21985 VGND.n1984 VGND.n1983 0.5525
R21986 VGND.n2067 VGND 0.548
R21987 VGND.n1796 VGND 0.4925
R21988 VGND VGND.n2055 0.4805
R21989 VGND.n955 VGND 0.4745
R21990 VGND.n1675 VGND.n1674 0.45275
R21991 VGND.n1772 VGND 0.4505
R21992 VGND.n2164 VGND 0.4505
R21993 VGND.n3409 VGND.n3408 0.4415
R21994 VGND.n3408 VGND.n197 0.4415
R21995 VGND.n1876 VGND.n197 0.4415
R21996 VGND.n1877 VGND.n1876 0.4415
R21997 VGND.n1877 VGND.n363 0.4415
R21998 VGND.n3274 VGND.n3273 0.4415
R21999 VGND.n1280 VGND.n1279 0.4415
R22000 VGND.n1279 VGND.n1239 0.4415
R22001 VGND.n1239 VGND.n1191 0.4415
R22002 VGND.n1191 VGND.n1113 0.4415
R22003 VGND.n1113 VGND.n1067 0.4415
R22004 VGND.n1067 VGND.n1014 0.4415
R22005 VGND.n1014 VGND.n419 0.4415
R22006 VGND.n2488 VGND.n419 0.4415
R22007 VGND.n2558 VGND.n2488 0.4415
R22008 VGND.n2600 VGND.n2558 0.4415
R22009 VGND.n2731 VGND.n2600 0.4415
R22010 VGND.n2731 VGND.n2730 0.4415
R22011 VGND.n2730 VGND.n2622 0.4415
R22012 VGND.n2622 VGND.n2611 0.4415
R22013 VGND.n2611 VGND.n384 0.4415
R22014 VGND.n2962 VGND.n384 0.4415
R22015 VGND.n2999 VGND.n2962 0.4415
R22016 VGND.n3000 VGND.n2999 0.4415
R22017 VGND.n1630 VGND.n837 0.4415
R22018 VGND.n1631 VGND.n1630 0.4415
R22019 VGND.n1631 VGND.n575 0.4415
R22020 VGND.n2002 VGND.n575 0.4415
R22021 VGND.n2003 VGND.n2002 0.4415
R22022 VGND.n2003 VGND.n427 0.4415
R22023 VGND.n2447 VGND.n427 0.4415
R22024 VGND.n2448 VGND.n2447 0.4415
R22025 VGND.n2448 VGND.n411 0.4415
R22026 VGND.n2826 VGND.n411 0.4415
R22027 VGND.n2826 VGND.n2825 0.4415
R22028 VGND.n2825 VGND.n378 0.4415
R22029 VGND.n3042 VGND.n3041 0.4415
R22030 VGND.n1597 VGND.n1596 0.4415
R22031 VGND.n1597 VGND.n588 0.4415
R22032 VGND.n1970 VGND.n588 0.4415
R22033 VGND.n1971 VGND.n1970 0.4415
R22034 VGND.n1971 VGND.n469 0.4415
R22035 VGND.n2411 VGND.n469 0.4415
R22036 VGND.n2412 VGND.n2411 0.4415
R22037 VGND.n2412 VGND.n407 0.4415
R22038 VGND.n2885 VGND.n407 0.4415
R22039 VGND.n2885 VGND.n2884 0.4415
R22040 VGND.n2884 VGND.n408 0.4415
R22041 VGND.n408 VGND.n374 0.4415
R22042 VGND.n3105 VGND.n3104 0.4415
R22043 VGND.n1562 VGND.n1561 0.4415
R22044 VGND.n1561 VGND.n612 0.4415
R22045 VGND.n1939 VGND.n612 0.4415
R22046 VGND.n1939 VGND.n1938 0.4415
R22047 VGND.n1938 VGND.n483 0.4415
R22048 VGND.n2383 VGND.n483 0.4415
R22049 VGND.n2383 VGND.n2382 0.4415
R22050 VGND.n2382 VGND.n484 0.4415
R22051 VGND.n484 VGND.n370 0.4415
R22052 VGND.n3146 VGND.n3145 0.4415
R22053 VGND.n3432 VGND.n141 0.4415
R22054 VGND.n1792 VGND.n141 0.4415
R22055 VGND.n1793 VGND.n1792 0.4415
R22056 VGND.n1793 VGND.n548 0.4415
R22057 VGND.n2168 VGND.n548 0.4415
R22058 VGND.n2221 VGND.n2168 0.4415
R22059 VGND.n2351 VGND.n2221 0.4415
R22060 VGND.n2351 VGND.n2350 0.4415
R22061 VGND.n2350 VGND.n367 0.4415
R22062 VGND.n3210 VGND.n3209 0.4415
R22063 VGND.n3379 VGND.n244 0.4415
R22064 VGND.n3379 VGND.n3378 0.4415
R22065 VGND.n3378 VGND.n245 0.4415
R22066 VGND.n359 VGND.n245 0.4415
R22067 VGND.n3337 VGND.n359 0.4415
R22068 VGND.n3336 VGND.n360 0.4415
R22069 VGND.n3685 VGND.n3684 0.4415
R22070 VGND.n3684 VGND.n3464 0.4415
R22071 VGND.n3665 VGND.n3464 0.4415
R22072 VGND.n3665 VGND.n3664 0.4415
R22073 VGND.n3664 VGND.n3649 0.4415
R22074 VGND.n3649 VGND.n3634 0.4415
R22075 VGND.n3634 VGND.n3618 0.4415
R22076 VGND.n3618 VGND.n3602 0.4415
R22077 VGND.n3602 VGND.n3586 0.4415
R22078 VGND.n3586 VGND.n3570 0.4415
R22079 VGND.n3570 VGND.n3554 0.4415
R22080 VGND.n3554 VGND.n3539 0.4415
R22081 VGND.n3539 VGND.n3524 0.4415
R22082 VGND.n3524 VGND.n3509 0.4415
R22083 VGND.n3509 VGND.n19 0.4415
R22084 VGND.n3715 VGND.n19 0.4415
R22085 VGND.n3717 VGND.n3715 0.4415
R22086 VGND.n3717 VGND.n3716 0.4415
R22087 VGND.n3756 VGND.n3755 0.4415
R22088 VGND.n953 VGND 0.4325
R22089 VGND.n2064 VGND 0.4325
R22090 VGND.n55 VGND.t102 0.429663
R22091 VGND VGND.n3411 0.4205
R22092 VGND VGND.n821 0.40325
R22093 VGND VGND.n1302 0.38675
R22094 VGND.n3451 VGND.t325 0.381978
R22095 VGND.n3421 VGND 0.3755
R22096 VGND.n3389 VGND 0.3725
R22097 VGND VGND.n835 0.36725
R22098 VGND.n355 VGND.n354 0.3665
R22099 VGND.n3697 VGND.n3696 0.3665
R22100 VGND VGND.n1926 0.3665
R22101 VGND.n2376 VGND.n2375 0.3665
R22102 VGND.n2950 VGND.n2949 0.3665
R22103 VGND.n2941 VGND.n2940 0.3665
R22104 VGND.n2931 VGND.n2930 0.3665
R22105 VGND.n3006 VGND.n3005 0.3665
R22106 VGND.n3018 VGND.n3017 0.3665
R22107 VGND.n3036 VGND.n3035 0.3665
R22108 VGND.n3027 VGND.n3026 0.3665
R22109 VGND.n3110 VGND.n3109 0.3665
R22110 VGND.n3123 VGND.n3122 0.3665
R22111 VGND.n3141 VGND.n3140 0.3665
R22112 VGND.n3132 VGND.n3131 0.3665
R22113 VGND.n3215 VGND.n3214 0.3665
R22114 VGND.n3229 VGND.n3228 0.3665
R22115 VGND.n3270 VGND.n3269 0.3665
R22116 VGND.n3261 VGND.n3260 0.3665
R22117 VGND.n3251 VGND.n3250 0.3665
R22118 VGND.n3242 VGND.n3241 0.3665
R22119 VGND.n3759 VGND.n3758 0.3665
R22120 VGND.n3775 VGND.n3774 0.3665
R22121 VGND.n3786 VGND.n3785 0.3665
R22122 VGND.n1396 VGND.n1395 0.3635
R22123 VGND.n3423 VGND.n3422 0.3635
R22124 VGND VGND.n297 0.3635
R22125 VGND.n321 VGND.n320 0.3635
R22126 VGND.n1461 VGND.n1460 0.3635
R22127 VGND.n1974 VGND.n1973 0.3635
R22128 VGND.n2199 VGND 0.3605
R22129 VGND VGND.n1764 0.3575
R22130 VGND.n881 VGND.n880 0.3545
R22131 VGND.n1685 VGND.n1684 0.3545
R22132 VGND.n2065 VGND.n2064 0.353
R22133 VGND VGND.n3384 0.3515
R22134 VGND.n2387 VGND 0.3515
R22135 VGND VGND.n485 0.3515
R22136 VGND.n1248 VGND 0.3485
R22137 VGND.n1599 VGND 0.3485
R22138 VGND.n1765 VGND 0.3395
R22139 VGND.n1981 VGND 0.338
R22140 VGND.n3681 VGND.n3680 0.3365
R22141 VGND.n3680 VGND.n3679 0.3365
R22142 VGND.n3679 VGND.n3678 0.3365
R22143 VGND.n3677 VGND.n3676 0.3365
R22144 VGND.n3676 VGND.n3675 0.3365
R22145 VGND.n3675 VGND.n3674 0.3365
R22146 VGND.n3493 VGND.n3492 0.3365
R22147 VGND.n3492 VGND.n3491 0.3365
R22148 VGND.n3491 VGND.n3490 0.3365
R22149 VGND.n3489 VGND.n3488 0.3365
R22150 VGND.n3488 VGND.n3487 0.3365
R22151 VGND.n3487 VGND.n3486 0.3365
R22152 VGND.n3646 VGND.n3645 0.3365
R22153 VGND.n3645 VGND.n3644 0.3365
R22154 VGND.n3644 VGND.n3643 0.3365
R22155 VGND.n3642 VGND.n3641 0.3365
R22156 VGND.n3641 VGND.n3640 0.3365
R22157 VGND.n3640 VGND.n3639 0.3365
R22158 VGND.n3661 VGND.n3660 0.3365
R22159 VGND.n3660 VGND.n3659 0.3365
R22160 VGND.n3659 VGND.n3658 0.3365
R22161 VGND.n3657 VGND.n3656 0.3365
R22162 VGND.n3656 VGND.n3655 0.3365
R22163 VGND.n3655 VGND.n3654 0.3365
R22164 VGND.n3476 VGND.n3475 0.3365
R22165 VGND.n3475 VGND.n3474 0.3365
R22166 VGND.n3474 VGND.n3473 0.3365
R22167 VGND.n3472 VGND.n3471 0.3365
R22168 VGND.n3471 VGND.n3470 0.3365
R22169 VGND.n3470 VGND.n3469 0.3365
R22170 VGND.n3583 VGND.n3582 0.3365
R22171 VGND.n3582 VGND.n3581 0.3365
R22172 VGND.n3581 VGND.n3580 0.3365
R22173 VGND.n3579 VGND.n3578 0.3365
R22174 VGND.n3578 VGND.n3577 0.3365
R22175 VGND.n3577 VGND.n3576 0.3365
R22176 VGND.n3615 VGND.n3614 0.3365
R22177 VGND.n3614 VGND.n3613 0.3365
R22178 VGND.n3613 VGND.n3612 0.3365
R22179 VGND.n3611 VGND.n3610 0.3365
R22180 VGND.n3610 VGND.n3609 0.3365
R22181 VGND.n3609 VGND.n3608 0.3365
R22182 VGND.n3631 VGND.n3630 0.3365
R22183 VGND.n3630 VGND.n3629 0.3365
R22184 VGND.n3629 VGND.n3628 0.3365
R22185 VGND.n3627 VGND.n3626 0.3365
R22186 VGND.n3626 VGND.n3625 0.3365
R22187 VGND.n3625 VGND.n3624 0.3365
R22188 VGND.n3599 VGND.n3598 0.3365
R22189 VGND.n3598 VGND.n3597 0.3365
R22190 VGND.n3597 VGND.n3596 0.3365
R22191 VGND.n3595 VGND.n3594 0.3365
R22192 VGND.n3594 VGND.n3593 0.3365
R22193 VGND.n3593 VGND.n3592 0.3365
R22194 VGND.n3567 VGND.n3566 0.3365
R22195 VGND.n3566 VGND.n3565 0.3365
R22196 VGND.n3565 VGND.n3564 0.3365
R22197 VGND.n3563 VGND.n3562 0.3365
R22198 VGND.n3562 VGND.n3561 0.3365
R22199 VGND.n3561 VGND.n3560 0.3365
R22200 VGND.n3551 VGND.n3550 0.3365
R22201 VGND.n3550 VGND.n3549 0.3365
R22202 VGND.n3549 VGND.n3548 0.3365
R22203 VGND.n3547 VGND.n3546 0.3365
R22204 VGND.n3546 VGND.n3545 0.3365
R22205 VGND.n3545 VGND.n3544 0.3365
R22206 VGND.n3712 VGND.n3711 0.3365
R22207 VGND.n3711 VGND.n3710 0.3365
R22208 VGND.n3710 VGND.n3709 0.3365
R22209 VGND.n3708 VGND.n3707 0.3365
R22210 VGND.n3707 VGND.n3706 0.3365
R22211 VGND.n3706 VGND.n3705 0.3365
R22212 VGND.n32 VGND.n31 0.3365
R22213 VGND.n31 VGND.n30 0.3365
R22214 VGND.n30 VGND.n29 0.3365
R22215 VGND.n28 VGND.n27 0.3365
R22216 VGND.n27 VGND.n26 0.3365
R22217 VGND.n26 VGND.n25 0.3365
R22218 VGND.n3506 VGND.n3505 0.3365
R22219 VGND.n3505 VGND.n3504 0.3365
R22220 VGND.n3504 VGND.n3503 0.3365
R22221 VGND.n3502 VGND.n3501 0.3365
R22222 VGND.n3501 VGND.n3500 0.3365
R22223 VGND.n3500 VGND.n3499 0.3365
R22224 VGND.n3521 VGND.n3520 0.3365
R22225 VGND.n3520 VGND.n3519 0.3365
R22226 VGND.n3519 VGND.n3518 0.3365
R22227 VGND.n3517 VGND.n3516 0.3365
R22228 VGND.n3516 VGND.n3515 0.3365
R22229 VGND.n3515 VGND.n3514 0.3365
R22230 VGND.n3536 VGND.n3535 0.3365
R22231 VGND.n3535 VGND.n3534 0.3365
R22232 VGND.n3534 VGND.n3533 0.3365
R22233 VGND.n3532 VGND.n3531 0.3365
R22234 VGND.n3531 VGND.n3530 0.3365
R22235 VGND.n3530 VGND.n3529 0.3365
R22236 VGND.n879 VGND.n878 0.3365
R22237 VGND.n878 VGND.n877 0.3365
R22238 VGND.n1412 VGND.n1411 0.3365
R22239 VGND.n1433 VGND.n1432 0.3365
R22240 VGND.n3460 VGND.n3459 0.3365
R22241 VGND.n3459 VGND.n3458 0.3365
R22242 VGND.n3458 VGND.n3457 0.3365
R22243 VGND.n3456 VGND.n3455 0.3365
R22244 VGND.n3455 VGND.n3454 0.3365
R22245 VGND.n3454 VGND.n3453 0.3365
R22246 VGND.n343 VGND.n342 0.3365
R22247 VGND.n344 VGND.n343 0.3365
R22248 VGND.n345 VGND.n344 0.3365
R22249 VGND.n354 VGND.n353 0.3365
R22250 VGND.n353 VGND.n352 0.3365
R22251 VGND.n352 VGND.n351 0.3365
R22252 VGND.n350 VGND.n349 0.3365
R22253 VGND.n349 VGND.n348 0.3365
R22254 VGND.n348 VGND.n347 0.3365
R22255 VGND.n3696 VGND.n3695 0.3365
R22256 VGND.n3695 VGND.n3694 0.3365
R22257 VGND.n3694 VGND.n3693 0.3365
R22258 VGND.n52 VGND.n51 0.3365
R22259 VGND.n51 VGND.n50 0.3365
R22260 VGND.n50 VGND.n49 0.3365
R22261 VGND.n49 VGND.n48 0.3365
R22262 VGND.n47 VGND.n46 0.3365
R22263 VGND.n46 VGND.n45 0.3365
R22264 VGND.n45 VGND.n44 0.3365
R22265 VGND.n1475 VGND.n1443 0.3365
R22266 VGND.n261 VGND.n260 0.3365
R22267 VGND.n264 VGND.n263 0.3365
R22268 VGND.n268 VGND.n267 0.3365
R22269 VGND.n1656 VGND.n1655 0.3365
R22270 VGND.n1659 VGND.n1658 0.3365
R22271 VGND.n1663 VGND.n1662 0.3365
R22272 VGND.n1673 VGND.n1672 0.3365
R22273 VGND.n1713 VGND.n1712 0.3365
R22274 VGND.n1738 VGND.n1737 0.3365
R22275 VGND.n3367 VGND.n3366 0.3365
R22276 VGND.n3366 VGND.n3365 0.3365
R22277 VGND.n3365 VGND.n3364 0.3365
R22278 VGND.n3363 VGND.n3362 0.3365
R22279 VGND.n3362 VGND.n3361 0.3365
R22280 VGND.n3361 VGND.n3360 0.3365
R22281 VGND.n1135 VGND.n1134 0.3365
R22282 VGND.n1134 VGND.n1133 0.3365
R22283 VGND.n1952 VGND.n1951 0.3365
R22284 VGND.n1944 VGND.n1943 0.3365
R22285 VGND.n762 VGND.n761 0.3365
R22286 VGND.n765 VGND.n764 0.3365
R22287 VGND.n1807 VGND.n1806 0.3365
R22288 VGND.n1831 VGND.n1830 0.3365
R22289 VGND.n1830 VGND.n1829 0.3365
R22290 VGND.n1829 VGND.n1828 0.3365
R22291 VGND.n1827 VGND.n1826 0.3365
R22292 VGND.n1826 VGND.n1825 0.3365
R22293 VGND.n1825 VGND.n1824 0.3365
R22294 VGND.n652 VGND.n651 0.3365
R22295 VGND.n651 VGND.n650 0.3365
R22296 VGND.n650 VGND.n649 0.3365
R22297 VGND.n1935 VGND.n1934 0.3365
R22298 VGND.n674 VGND.n673 0.3365
R22299 VGND.n673 VGND.n672 0.3365
R22300 VGND.n672 VGND.n671 0.3365
R22301 VGND.n670 VGND.n669 0.3365
R22302 VGND.n669 VGND.n668 0.3365
R22303 VGND.n668 VGND.n667 0.3365
R22304 VGND.n1005 VGND.n1004 0.3365
R22305 VGND.n1004 VGND.n1003 0.3365
R22306 VGND.n1002 VGND.n1001 0.3365
R22307 VGND.n1000 VGND.n999 0.3365
R22308 VGND.n2192 VGND.n2191 0.3365
R22309 VGND.n2215 VGND.n2214 0.3365
R22310 VGND.n2214 VGND.n2213 0.3365
R22311 VGND.n2213 VGND.n2212 0.3365
R22312 VGND.n2211 VGND.n2210 0.3365
R22313 VGND.n2210 VGND.n2209 0.3365
R22314 VGND.n2209 VGND.n2208 0.3365
R22315 VGND.n2870 VGND.n2869 0.3365
R22316 VGND.n2869 VGND.n2868 0.3365
R22317 VGND.n2868 VGND.n2867 0.3365
R22318 VGND.n2866 VGND.n2865 0.3365
R22319 VGND.n2865 VGND.n2864 0.3365
R22320 VGND.n2864 VGND.n2863 0.3365
R22321 VGND.n2614 VGND.n2613 0.3365
R22322 VGND.n2620 VGND.n2619 0.3365
R22323 VGND.n2618 VGND.n2617 0.3365
R22324 VGND.n2617 VGND.n2616 0.3365
R22325 VGND.n2616 VGND.n2615 0.3365
R22326 VGND.n2603 VGND.n2602 0.3365
R22327 VGND.n2609 VGND.n2608 0.3365
R22328 VGND.n2607 VGND.n2606 0.3365
R22329 VGND.n2606 VGND.n2605 0.3365
R22330 VGND.n2605 VGND.n2604 0.3365
R22331 VGND.n392 VGND.n391 0.3365
R22332 VGND.n395 VGND.n394 0.3365
R22333 VGND.n397 VGND.n396 0.3365
R22334 VGND.n398 VGND.n397 0.3365
R22335 VGND.n399 VGND.n398 0.3365
R22336 VGND.n386 VGND.n385 0.3365
R22337 VGND.n2960 VGND.n2959 0.3365
R22338 VGND.n2958 VGND.n2957 0.3365
R22339 VGND.n2957 VGND.n2956 0.3365
R22340 VGND.n2956 VGND.n2955 0.3365
R22341 VGND.n2774 VGND.n2773 0.3365
R22342 VGND.n2773 VGND.n2772 0.3365
R22343 VGND.n2772 VGND.n2771 0.3365
R22344 VGND.n2770 VGND.n2769 0.3365
R22345 VGND.n2769 VGND.n2768 0.3365
R22346 VGND.n2768 VGND.n2767 0.3365
R22347 VGND.n2642 VGND.n2641 0.3365
R22348 VGND.n2641 VGND.n2640 0.3365
R22349 VGND.n2640 VGND.n2639 0.3365
R22350 VGND.n2638 VGND.n2637 0.3365
R22351 VGND.n2637 VGND.n2636 0.3365
R22352 VGND.n2636 VGND.n2635 0.3365
R22353 VGND.n443 VGND.n442 0.3365
R22354 VGND.n444 VGND.n443 0.3365
R22355 VGND.n445 VGND.n444 0.3365
R22356 VGND.n448 VGND.n447 0.3365
R22357 VGND.n449 VGND.n448 0.3365
R22358 VGND.n513 VGND.n512 0.3365
R22359 VGND.n2370 VGND.n2369 0.3365
R22360 VGND.n539 VGND.n538 0.3365
R22361 VGND.n538 VGND.n537 0.3365
R22362 VGND.n537 VGND.n536 0.3365
R22363 VGND.n535 VGND.n534 0.3365
R22364 VGND.n534 VGND.n533 0.3365
R22365 VGND.n533 VGND.n532 0.3365
R22366 VGND.n2340 VGND.n2339 0.3365
R22367 VGND.n2339 VGND.n2338 0.3365
R22368 VGND.n2338 VGND.n2337 0.3365
R22369 VGND.n2336 VGND.n2335 0.3365
R22370 VGND.n2335 VGND.n2334 0.3365
R22371 VGND.n2334 VGND.n2333 0.3365
R22372 VGND.n2491 VGND.n2490 0.3365
R22373 VGND.n2556 VGND.n2555 0.3365
R22374 VGND.n2554 VGND.n2553 0.3365
R22375 VGND.n2512 VGND.n2511 0.3365
R22376 VGND.n2511 VGND.n2510 0.3365
R22377 VGND.n2510 VGND.n2509 0.3365
R22378 VGND.n2507 VGND.n2506 0.3365
R22379 VGND.n2506 VGND.n2505 0.3365
R22380 VGND.n2500 VGND.n2499 0.3365
R22381 VGND.n2499 VGND.n2498 0.3365
R22382 VGND.n2888 VGND.n2887 0.3365
R22383 VGND.n2889 VGND.n2888 0.3365
R22384 VGND.n2890 VGND.n2889 0.3365
R22385 VGND.n2910 VGND.n2909 0.3365
R22386 VGND.n2913 VGND.n2912 0.3365
R22387 VGND.n2914 VGND.n2913 0.3365
R22388 VGND.n2918 VGND.n2917 0.3365
R22389 VGND.n2919 VGND.n2918 0.3365
R22390 VGND.n2949 VGND.n2948 0.3365
R22391 VGND.n2948 VGND.n2947 0.3365
R22392 VGND.n2947 VGND.n2946 0.3365
R22393 VGND.n2945 VGND.n2944 0.3365
R22394 VGND.n2944 VGND.n2943 0.3365
R22395 VGND.n2943 VGND.n2942 0.3365
R22396 VGND.n2940 VGND.n2939 0.3365
R22397 VGND.n2939 VGND.n2938 0.3365
R22398 VGND.n2938 VGND.n2937 0.3365
R22399 VGND.n2934 VGND.n2933 0.3365
R22400 VGND.n2933 VGND.n2932 0.3365
R22401 VGND.n2930 VGND.n2929 0.3365
R22402 VGND.n2929 VGND.n2928 0.3365
R22403 VGND.n2928 VGND.n2927 0.3365
R22404 VGND.n2926 VGND.n2925 0.3365
R22405 VGND.n2925 VGND.n2924 0.3365
R22406 VGND.n2924 VGND.n2923 0.3365
R22407 VGND.n3350 VGND.n3349 0.3365
R22408 VGND.n3351 VGND.n3350 0.3365
R22409 VGND.n3352 VGND.n3351 0.3365
R22410 VGND.n3354 VGND.n3353 0.3365
R22411 VGND.n3355 VGND.n3354 0.3365
R22412 VGND.n3356 VGND.n3355 0.3365
R22413 VGND.n2990 VGND.n2989 0.3365
R22414 VGND.n2989 VGND.n2988 0.3365
R22415 VGND.n2988 VGND.n2987 0.3365
R22416 VGND.n2977 VGND.n2976 0.3365
R22417 VGND.n2976 VGND.n2975 0.3365
R22418 VGND.n2975 VGND.n2974 0.3365
R22419 VGND.n2974 VGND.n2973 0.3365
R22420 VGND.n3045 VGND.n3044 0.3365
R22421 VGND.n3046 VGND.n3045 0.3365
R22422 VGND.n3060 VGND.n3059 0.3365
R22423 VGND.n3061 VGND.n3060 0.3365
R22424 VGND.n3097 VGND.n3096 0.3365
R22425 VGND.n3096 VGND.n3095 0.3365
R22426 VGND.n3095 VGND.n3094 0.3365
R22427 VGND.n3094 VGND.n3093 0.3365
R22428 VGND.n3084 VGND.n3083 0.3365
R22429 VGND.n3083 VGND.n3082 0.3365
R22430 VGND.n3082 VGND.n3081 0.3365
R22431 VGND.n3081 VGND.n3080 0.3365
R22432 VGND.n3079 VGND.n3078 0.3365
R22433 VGND.n3149 VGND.n3148 0.3365
R22434 VGND.n3165 VGND.n3164 0.3365
R22435 VGND.n3203 VGND.n3202 0.3365
R22436 VGND.n3202 VGND.n3201 0.3365
R22437 VGND.n3201 VGND.n3200 0.3365
R22438 VGND.n3200 VGND.n3199 0.3365
R22439 VGND.n3198 VGND.n3197 0.3365
R22440 VGND.n3191 VGND.n3190 0.3365
R22441 VGND.n3190 VGND.n3189 0.3365
R22442 VGND.n3189 VGND.n3188 0.3365
R22443 VGND.n3188 VGND.n3187 0.3365
R22444 VGND.n3186 VGND.n3185 0.3365
R22445 VGND.n3185 VGND.n3184 0.3365
R22446 VGND.n3332 VGND.n3331 0.3365
R22447 VGND.n3331 VGND.n3330 0.3365
R22448 VGND.n3330 VGND.n3329 0.3365
R22449 VGND.n3329 VGND.n3328 0.3365
R22450 VGND.n3327 VGND.n3326 0.3365
R22451 VGND.n3326 VGND.n3325 0.3365
R22452 VGND.n3321 VGND.n3320 0.3365
R22453 VGND.n3320 VGND.n3319 0.3365
R22454 VGND.n3319 VGND.n3318 0.3365
R22455 VGND.n3318 VGND.n3317 0.3365
R22456 VGND.n3316 VGND.n3315 0.3365
R22457 VGND.n3315 VGND.n3314 0.3365
R22458 VGND.n3314 VGND.n4 0.3365
R22459 VGND.n16 VGND.n15 0.3365
R22460 VGND.n15 VGND.n14 0.3365
R22461 VGND.n14 VGND.n13 0.3365
R22462 VGND.n12 VGND.n11 0.3365
R22463 VGND.n11 VGND.n10 0.3365
R22464 VGND.n10 VGND.n9 0.3365
R22465 VGND.n383 VGND.n382 0.3365
R22466 VGND.n3004 VGND.n3003 0.3365
R22467 VGND.n3007 VGND.n3006 0.3365
R22468 VGND.n3008 VGND.n3007 0.3365
R22469 VGND.n3009 VGND.n3008 0.3365
R22470 VGND.n3011 VGND.n3010 0.3365
R22471 VGND.n3012 VGND.n3011 0.3365
R22472 VGND.n3013 VGND.n3012 0.3365
R22473 VGND.n3017 VGND.n3016 0.3365
R22474 VGND.n3016 VGND.n3015 0.3365
R22475 VGND.n3015 VGND.n3014 0.3365
R22476 VGND.n3039 VGND.n3038 0.3365
R22477 VGND.n3038 VGND.n3037 0.3365
R22478 VGND.n3035 VGND.n3034 0.3365
R22479 VGND.n3034 VGND.n3033 0.3365
R22480 VGND.n3033 VGND.n3032 0.3365
R22481 VGND.n3031 VGND.n3030 0.3365
R22482 VGND.n3030 VGND.n3029 0.3365
R22483 VGND.n3029 VGND.n3028 0.3365
R22484 VGND.n3026 VGND.n3025 0.3365
R22485 VGND.n3025 VGND.n3024 0.3365
R22486 VGND.n3024 VGND.n3023 0.3365
R22487 VGND.n3022 VGND.n373 0.3365
R22488 VGND.n3108 VGND.n3107 0.3365
R22489 VGND.n3111 VGND.n3110 0.3365
R22490 VGND.n3112 VGND.n3111 0.3365
R22491 VGND.n3113 VGND.n3112 0.3365
R22492 VGND.n3115 VGND.n3114 0.3365
R22493 VGND.n3116 VGND.n3115 0.3365
R22494 VGND.n3117 VGND.n3116 0.3365
R22495 VGND.n3122 VGND.n3121 0.3365
R22496 VGND.n3121 VGND.n3120 0.3365
R22497 VGND.n3120 VGND.n3119 0.3365
R22498 VGND.n3118 VGND.n371 0.3365
R22499 VGND.n3143 VGND.n3142 0.3365
R22500 VGND.n3140 VGND.n3139 0.3365
R22501 VGND.n3139 VGND.n3138 0.3365
R22502 VGND.n3138 VGND.n3137 0.3365
R22503 VGND.n3136 VGND.n3135 0.3365
R22504 VGND.n3135 VGND.n3134 0.3365
R22505 VGND.n3134 VGND.n3133 0.3365
R22506 VGND.n3131 VGND.n3130 0.3365
R22507 VGND.n3130 VGND.n3129 0.3365
R22508 VGND.n3129 VGND.n3128 0.3365
R22509 VGND.n3127 VGND.n366 0.3365
R22510 VGND.n3213 VGND.n3212 0.3365
R22511 VGND.n3216 VGND.n3215 0.3365
R22512 VGND.n3217 VGND.n3216 0.3365
R22513 VGND.n3218 VGND.n3217 0.3365
R22514 VGND.n3220 VGND.n3219 0.3365
R22515 VGND.n3221 VGND.n3220 0.3365
R22516 VGND.n3222 VGND.n3221 0.3365
R22517 VGND.n3228 VGND.n3227 0.3365
R22518 VGND.n3227 VGND.n3226 0.3365
R22519 VGND.n3226 VGND.n3225 0.3365
R22520 VGND.n3224 VGND.n3223 0.3365
R22521 VGND.n3223 VGND.n364 0.3365
R22522 VGND.n3269 VGND.n3268 0.3365
R22523 VGND.n3268 VGND.n3267 0.3365
R22524 VGND.n3267 VGND.n3266 0.3365
R22525 VGND.n3265 VGND.n3264 0.3365
R22526 VGND.n3264 VGND.n3263 0.3365
R22527 VGND.n3263 VGND.n3262 0.3365
R22528 VGND.n3260 VGND.n3259 0.3365
R22529 VGND.n3259 VGND.n3258 0.3365
R22530 VGND.n3258 VGND.n3257 0.3365
R22531 VGND.n3256 VGND.n3255 0.3365
R22532 VGND.n3255 VGND.n3254 0.3365
R22533 VGND.n3250 VGND.n3249 0.3365
R22534 VGND.n3249 VGND.n3248 0.3365
R22535 VGND.n3248 VGND.n3247 0.3365
R22536 VGND.n3246 VGND.n3245 0.3365
R22537 VGND.n3245 VGND.n3244 0.3365
R22538 VGND.n3244 VGND.n3243 0.3365
R22539 VGND.n3241 VGND.n3240 0.3365
R22540 VGND.n3240 VGND.n3239 0.3365
R22541 VGND.n3239 VGND.n3238 0.3365
R22542 VGND.n3237 VGND.n3236 0.3365
R22543 VGND.n3236 VGND.n3235 0.3365
R22544 VGND.n3235 VGND.n2 0.3365
R22545 VGND.n3760 VGND.n3759 0.3365
R22546 VGND.n3761 VGND.n3760 0.3365
R22547 VGND.n3762 VGND.n3761 0.3365
R22548 VGND.n3764 VGND.n3763 0.3365
R22549 VGND.n3765 VGND.n3764 0.3365
R22550 VGND.n3766 VGND.n3765 0.3365
R22551 VGND.n3774 VGND.n3773 0.3365
R22552 VGND.n3773 VGND.n3772 0.3365
R22553 VGND.n3772 VGND.n3771 0.3365
R22554 VGND.n3770 VGND.n3769 0.3365
R22555 VGND.n3769 VGND.n3768 0.3365
R22556 VGND.n3768 VGND.n3767 0.3365
R22557 VGND.n3785 VGND.n3784 0.3365
R22558 VGND.n3784 VGND.n3783 0.3365
R22559 VGND.n3783 VGND.n3782 0.3365
R22560 VGND.n3781 VGND.n3780 0.3365
R22561 VGND.n3780 VGND.n3779 0.3365
R22562 VGND.n3779 VGND.n3778 0.3365
R22563 VGND.t5880 VGND.t6 0.334293
R22564 VGND VGND.n3413 0.33425
R22565 VGND VGND.n1817 0.33425
R22566 VGND.n2054 VGND 0.33425
R22567 VGND VGND.n1435 0.3335
R22568 VGND.n3424 VGND.n3423 0.3335
R22569 VGND VGND.n3417 0.3335
R22570 VGND.n1533 VGND.n1532 0.3335
R22571 VGND.n653 VGND.n652 0.3335
R22572 VGND VGND.n2400 0.3335
R22573 VGND.n2202 VGND.n2201 0.3335
R22574 VGND.n3211 VGND.n366 0.3335
R22575 VGND.n1302 VGND.n1301 0.33125
R22576 VGND.n1530 VGND.n1529 0.3305
R22577 VGND.n2403 VGND.n2402 0.3305
R22578 VGND.n2373 VGND.n2372 0.3305
R22579 VGND.n741 VGND.n611 0.32975
R22580 VGND.n1945 VGND.n1944 0.326
R22581 VGND.n192 VGND.n191 0.3245
R22582 VGND VGND.n236 0.3245
R22583 VGND.n1581 VGND 0.3245
R22584 VGND.n1552 VGND.n1551 0.3245
R22585 VGND.n1522 VGND 0.3245
R22586 VGND VGND.n3681 0.32225
R22587 VGND VGND.n3493 0.32225
R22588 VGND VGND.n3646 0.32225
R22589 VGND VGND.n3661 0.32225
R22590 VGND VGND.n3476 0.32225
R22591 VGND VGND.n3583 0.32225
R22592 VGND VGND.n3615 0.32225
R22593 VGND VGND.n3631 0.32225
R22594 VGND VGND.n3599 0.32225
R22595 VGND VGND.n3567 0.32225
R22596 VGND VGND.n3551 0.32225
R22597 VGND VGND.n3712 0.32225
R22598 VGND VGND.n32 0.32225
R22599 VGND VGND.n3506 0.32225
R22600 VGND VGND.n3521 0.32225
R22601 VGND VGND.n3536 0.32225
R22602 VGND.n304 VGND 0.32225
R22603 VGND VGND.n1477 0.32225
R22604 VGND VGND.n1538 0.32225
R22605 VGND.n260 VGND 0.32225
R22606 VGND VGND.n1006 0.32225
R22607 VGND VGND.n2215 0.32225
R22608 VGND.n2613 VGND 0.32225
R22609 VGND.n2602 VGND 0.32225
R22610 VGND.n391 VGND 0.32225
R22611 VGND VGND.n386 0.32225
R22612 VGND VGND.n2642 0.32225
R22613 VGND VGND.n2462 0.32225
R22614 VGND.n2042 VGND 0.32225
R22615 VGND.n3349 VGND 0.32225
R22616 VGND.n381 VGND 0.32225
R22617 VGND.n1658 VGND.n1657 0.3215
R22618 VGND.n632 VGND.n631 0.3215
R22619 VGND.n2385 VGND 0.3185
R22620 VGND.n3040 VGND.n379 0.314
R22621 VGND.n1440 VGND.n1439 0.3125
R22622 VGND.n1811 VGND.n1810 0.3125
R22623 VGND.n1566 VGND.n1565 0.3095
R22624 VGND.n3395 VGND.n3394 0.3095
R22625 VGND.n766 VGND.n765 0.3095
R22626 VGND.n2557 VGND.n2556 0.3095
R22627 VGND VGND.n1429 0.3065
R22628 VGND VGND.n1583 0.3065
R22629 VGND.n1251 VGND 0.3065
R22630 VGND.n1126 VGND 0.3065
R22631 VGND VGND.n1975 0.3065
R22632 VGND.n1927 VGND 0.3065
R22633 VGND.n882 VGND 0.305
R22634 VGND.n1875 VGND.n1874 0.305
R22635 VGND.n1963 VGND.n1962 0.3035
R22636 VGND.n1305 VGND 0.3005
R22637 VGND.n263 VGND.n262 0.3005
R22638 VGND VGND.n187 0.29825
R22639 VGND VGND.n1297 0.29825
R22640 VGND.n313 VGND.n312 0.29825
R22641 VGND.n1800 VGND 0.29825
R22642 VGND.n1666 VGND.n1665 0.2975
R22643 VGND VGND.n1693 0.2975
R22644 VGND.n1435 VGND.n1434 0.2945
R22645 VGND.n876 VGND.n875 0.2915
R22646 VGND.n1565 VGND.n1564 0.2915
R22647 VGND.n3425 VGND.n3424 0.2915
R22648 VGND.n1661 VGND.n1660 0.2915
R22649 VGND.n1687 VGND.n1686 0.2915
R22650 VGND.n760 VGND.n759 0.2915
R22651 VGND.n2917 VGND.n2916 0.29
R22652 VGND.n1408 VGND.n1407 0.2885
R22653 VGND.n1808 VGND.n1807 0.2885
R22654 VGND VGND.n1940 0.287
R22655 VGND.n742 VGND.n741 0.28625
R22656 VGND.n1954 VGND.n1953 0.2855
R22657 VGND VGND.n190 0.2825
R22658 VGND.n1384 VGND 0.2825
R22659 VGND.n305 VGND 0.2825
R22660 VGND.n334 VGND.n333 0.2825
R22661 VGND VGND.n1550 0.2825
R22662 VGND.n269 VGND 0.2825
R22663 VGND.n1672 VGND.n1671 0.2825
R22664 VGND VGND.n1713 0.2825
R22665 VGND VGND.n1711 0.2825
R22666 VGND.n1753 VGND 0.2825
R22667 VGND VGND.n1135 0.2825
R22668 VGND.n1810 VGND 0.2825
R22669 VGND VGND.n1871 0.2825
R22670 VGND VGND.n1987 0.2825
R22671 VGND VGND.n1913 0.2825
R22672 VGND VGND.n1005 0.2825
R22673 VGND.n2396 VGND 0.2825
R22674 VGND.n2201 VGND 0.2825
R22675 VGND.n2628 VGND.n2627 0.2825
R22676 VGND.n2715 VGND.n2714 0.2825
R22677 VGND VGND.n2439 0.2825
R22678 VGND VGND.n2438 0.2825
R22679 VGND VGND.n2489 0.2825
R22680 VGND VGND.n2554 0.2825
R22681 VGND VGND.n2512 0.2825
R22682 VGND.n2076 VGND 0.2825
R22683 VGND.n2081 VGND 0.2825
R22684 VGND.n2158 VGND.n2157 0.2825
R22685 VGND.n382 VGND 0.2825
R22686 VGND.n3003 VGND 0.2825
R22687 VGND VGND.n3677 0.28175
R22688 VGND VGND.n3489 0.28175
R22689 VGND VGND.n3642 0.28175
R22690 VGND VGND.n3657 0.28175
R22691 VGND VGND.n3472 0.28175
R22692 VGND VGND.n3579 0.28175
R22693 VGND VGND.n3611 0.28175
R22694 VGND VGND.n3627 0.28175
R22695 VGND VGND.n3595 0.28175
R22696 VGND VGND.n3563 0.28175
R22697 VGND VGND.n3547 0.28175
R22698 VGND VGND.n3708 0.28175
R22699 VGND VGND.n28 0.28175
R22700 VGND VGND.n3502 0.28175
R22701 VGND VGND.n3517 0.28175
R22702 VGND VGND.n3532 0.28175
R22703 VGND VGND.n3456 0.28175
R22704 VGND.n342 VGND 0.28175
R22705 VGND VGND.n350 0.28175
R22706 VGND VGND.n3692 0.28175
R22707 VGND VGND.n47 0.28175
R22708 VGND VGND.n3363 0.28175
R22709 VGND VGND.n1136 0.28175
R22710 VGND VGND.n1827 0.28175
R22711 VGND VGND.n670 0.28175
R22712 VGND VGND.n1002 0.28175
R22713 VGND VGND.n1000 0.28175
R22714 VGND VGND.n2211 0.28175
R22715 VGND VGND.n2866 0.28175
R22716 VGND VGND.n2618 0.28175
R22717 VGND VGND.n2607 0.28175
R22718 VGND.n396 VGND 0.28175
R22719 VGND VGND.n2958 0.28175
R22720 VGND VGND.n2770 0.28175
R22721 VGND VGND.n2638 0.28175
R22722 VGND.n446 VGND 0.28175
R22723 VGND.n447 VGND 0.28175
R22724 VGND VGND.n535 0.28175
R22725 VGND VGND.n2336 0.28175
R22726 VGND VGND.n2508 0.28175
R22727 VGND VGND.n2507 0.28175
R22728 VGND.n2915 VGND 0.28175
R22729 VGND VGND.n2945 0.28175
R22730 VGND VGND.n2936 0.28175
R22731 VGND VGND.n2926 0.28175
R22732 VGND.n3353 VGND 0.28175
R22733 VGND VGND.n2990 0.28175
R22734 VGND VGND.n2972 0.28175
R22735 VGND VGND.n3092 0.28175
R22736 VGND VGND.n3079 0.28175
R22737 VGND VGND.n3198 0.28175
R22738 VGND VGND.n3186 0.28175
R22739 VGND VGND.n3327 0.28175
R22740 VGND VGND.n3316 0.28175
R22741 VGND VGND.n12 0.28175
R22742 VGND.n3010 VGND 0.28175
R22743 VGND VGND.n379 0.28175
R22744 VGND VGND.n3031 0.28175
R22745 VGND VGND.n3022 0.28175
R22746 VGND.n3114 VGND 0.28175
R22747 VGND VGND.n3118 0.28175
R22748 VGND VGND.n3136 0.28175
R22749 VGND VGND.n3127 0.28175
R22750 VGND.n3219 VGND 0.28175
R22751 VGND VGND.n3224 0.28175
R22752 VGND VGND.n3265 0.28175
R22753 VGND VGND.n3256 0.28175
R22754 VGND VGND.n3246 0.28175
R22755 VGND VGND.n3237 0.28175
R22756 VGND.n3763 VGND 0.28175
R22757 VGND VGND.n3770 0.28175
R22758 VGND VGND.n3781 0.28175
R22759 VGND VGND.n3460 0.281
R22760 VGND VGND.n3367 0.281
R22761 VGND VGND.n1831 0.281
R22762 VGND VGND.n674 0.281
R22763 VGND VGND.n2870 0.281
R22764 VGND VGND.n2774 0.281
R22765 VGND VGND.n2661 0.281
R22766 VGND VGND.n539 0.281
R22767 VGND VGND.n2340 0.281
R22768 VGND VGND.n2104 0.281
R22769 VGND VGND.n16 0.281
R22770 VGND.n856 VGND.n855 0.2795
R22771 VGND.n341 VGND.n340 0.2795
R22772 VGND.n1791 VGND 0.2795
R22773 VGND.n1744 VGND.n1743 0.2795
R22774 VGND.n2187 VGND.n2186 0.2795
R22775 VGND.n1453 VGND.n1452 0.27725
R22776 VGND.n884 VGND.n883 0.2765
R22777 VGND.n238 VGND.n237 0.2765
R22778 VGND VGND.n108 0.2765
R22779 VGND.n1400 VGND.n1399 0.2765
R22780 VGND.n3420 VGND.n3419 0.2765
R22781 VGND VGND.n296 0.2765
R22782 VGND.n3393 VGND.n3392 0.2765
R22783 VGND.n266 VGND.n265 0.2765
R22784 VGND.n1652 VGND.n1651 0.2765
R22785 VGND.n1760 VGND.n1759 0.2765
R22786 VGND VGND.n962 0.2765
R22787 VGND VGND.n819 0.27425
R22788 VGND VGND.n632 0.27425
R22789 VGND.n1410 VGND.n1409 0.2705
R22790 VGND.n1786 VGND.n1785 0.2675
R22791 VGND.n2381 VGND.n2380 0.266
R22792 VGND.n1413 VGND.n1412 0.2645
R22793 VGND.n223 VGND.n222 0.2645
R22794 VGND VGND.n224 0.2645
R22795 VGND.n3391 VGND.n3390 0.2645
R22796 VGND VGND.n1699 0.2645
R22797 VGND.n1969 VGND.n590 0.2645
R22798 VGND.n1987 VGND 0.2645
R22799 VGND VGND.n1976 0.2645
R22800 VGND.n1909 VGND.n1908 0.2645
R22801 VGND.n2374 VGND.n2373 0.2645
R22802 VGND VGND.n2043 0.2645
R22803 VGND.n2088 VGND.n2087 0.2645
R22804 VGND VGND.n1430 0.26225
R22805 VGND.n2068 VGND 0.26075
R22806 VGND.n1481 VGND.n1480 0.25925
R22807 VGND.n1958 VGND.n1957 0.2585
R22808 VGND.n3043 VGND 0.2585
R22809 VGND.n2377 VGND 0.257
R22810 VGND.n821 VGND.n820 0.2555
R22811 VGND VGND.n2089 0.2555
R22812 VGND VGND.n1211 0.25475
R22813 VGND.n74 VGND.n73 0.2525
R22814 VGND.n76 VGND.n75 0.2525
R22815 VGND.n331 VGND.n330 0.2525
R22816 VGND.n336 VGND.n335 0.2525
R22817 VGND.n338 VGND.n337 0.2525
R22818 VGND.n1258 VGND.n1257 0.2525
R22819 VGND VGND.n1543 0.2525
R22820 VGND.n3399 VGND 0.2525
R22821 VGND.n1220 VGND.n1219 0.2525
R22822 VGND.n1650 VGND.n1649 0.2525
R22823 VGND.n1779 VGND.n1778 0.2525
R22824 VGND.n1749 VGND.n1748 0.2525
R22825 VGND.n1746 VGND.n1745 0.2525
R22826 VGND.n1741 VGND 0.2525
R22827 VGND.n3374 VGND.n3373 0.2525
R22828 VGND.n1867 VGND.n1866 0.2525
R22829 VGND.n1865 VGND.n1864 0.2525
R22830 VGND.n1863 VGND.n1862 0.2525
R22831 VGND.n1859 VGND.n1858 0.2525
R22832 VGND.n1857 VGND.n1856 0.2525
R22833 VGND.n1855 VGND.n1854 0.2525
R22834 VGND.n1849 VGND.n1848 0.2525
R22835 VGND.n1847 VGND.n1846 0.2525
R22836 VGND.n1845 VGND.n1844 0.2525
R22837 VGND.n1840 VGND.n1839 0.2525
R22838 VGND.n1838 VGND.n1837 0.2525
R22839 VGND.n1836 VGND.n1835 0.2525
R22840 VGND.n1905 VGND 0.2525
R22841 VGND.n1898 VGND.n1897 0.2525
R22842 VGND.n1896 VGND.n1895 0.2525
R22843 VGND.n1892 VGND.n1891 0.2525
R22844 VGND.n1886 VGND.n1885 0.2525
R22845 VGND.n1884 VGND.n1883 0.2525
R22846 VGND.n1882 VGND.n1881 0.2525
R22847 VGND.n1880 VGND.n1879 0.2525
R22848 VGND.n720 VGND.n719 0.2525
R22849 VGND.n718 VGND.n717 0.2525
R22850 VGND.n716 VGND.n715 0.2525
R22851 VGND.n710 VGND.n709 0.2525
R22852 VGND.n708 VGND.n707 0.2525
R22853 VGND.n706 VGND.n705 0.2525
R22854 VGND.n704 VGND.n703 0.2525
R22855 VGND.n702 VGND.n701 0.2525
R22856 VGND.n700 VGND.n699 0.2525
R22857 VGND.n698 VGND.n697 0.2525
R22858 VGND.n692 VGND.n691 0.2525
R22859 VGND.n690 VGND.n689 0.2525
R22860 VGND.n688 VGND.n687 0.2525
R22861 VGND.n683 VGND.n682 0.2525
R22862 VGND.n681 VGND.n680 0.2525
R22863 VGND.n679 VGND.n678 0.2525
R22864 VGND.n940 VGND.n939 0.2525
R22865 VGND.n938 VGND.n937 0.2525
R22866 VGND.n1011 VGND.n1010 0.2525
R22867 VGND.n2393 VGND 0.2525
R22868 VGND.n2564 VGND.n2563 0.2525
R22869 VGND.n2562 VGND.n2561 0.2525
R22870 VGND.n2560 VGND.n2559 0.2525
R22871 VGND.n2596 VGND.n2595 0.2525
R22872 VGND.n2594 VGND.n2593 0.2525
R22873 VGND.n2592 VGND.n2591 0.2525
R22874 VGND.n2586 VGND.n2585 0.2525
R22875 VGND.n2584 VGND.n2583 0.2525
R22876 VGND.n2582 VGND.n2581 0.2525
R22877 VGND.n2580 VGND.n2579 0.2525
R22878 VGND.n2578 VGND.n2577 0.2525
R22879 VGND.n2576 VGND.n2575 0.2525
R22880 VGND.n2574 VGND.n2573 0.2525
R22881 VGND.n2568 VGND.n2567 0.2525
R22882 VGND.n2566 VGND.n2565 0.2525
R22883 VGND.n2830 VGND.n2829 0.2525
R22884 VGND.n2832 VGND.n2831 0.2525
R22885 VGND.n2834 VGND.n2833 0.2525
R22886 VGND.n2836 VGND.n2835 0.2525
R22887 VGND.n2842 VGND.n2841 0.2525
R22888 VGND.n2844 VGND.n2843 0.2525
R22889 VGND.n2846 VGND.n2845 0.2525
R22890 VGND.n2848 VGND.n2847 0.2525
R22891 VGND.n2850 VGND.n2849 0.2525
R22892 VGND.n2852 VGND.n2851 0.2525
R22893 VGND.n2854 VGND.n2853 0.2525
R22894 VGND.n2859 VGND.n2858 0.2525
R22895 VGND.n2857 VGND.n2856 0.2525
R22896 VGND.n2881 VGND.n2880 0.2525
R22897 VGND.n2879 VGND.n2878 0.2525
R22898 VGND.n2877 VGND.n2876 0.2525
R22899 VGND.n2875 VGND.n2874 0.2525
R22900 VGND.n414 VGND.n413 0.2525
R22901 VGND.n416 VGND.n415 0.2525
R22902 VGND.n418 VGND.n417 0.2525
R22903 VGND.n2736 VGND.n2735 0.2525
R22904 VGND.n2738 VGND.n2737 0.2525
R22905 VGND.n2740 VGND.n2739 0.2525
R22906 VGND.n2746 VGND.n2745 0.2525
R22907 VGND.n2748 VGND.n2747 0.2525
R22908 VGND.n2750 VGND.n2749 0.2525
R22909 VGND.n2752 VGND.n2751 0.2525
R22910 VGND.n2754 VGND.n2753 0.2525
R22911 VGND.n2756 VGND.n2755 0.2525
R22912 VGND.n2758 VGND.n2757 0.2525
R22913 VGND.n2763 VGND.n2762 0.2525
R22914 VGND.n2761 VGND.n2760 0.2525
R22915 VGND.n2822 VGND.n2821 0.2525
R22916 VGND.n2820 VGND.n2819 0.2525
R22917 VGND.n2818 VGND.n2817 0.2525
R22918 VGND.n2816 VGND.n2815 0.2525
R22919 VGND.n2810 VGND.n2809 0.2525
R22920 VGND.n2808 VGND.n2807 0.2525
R22921 VGND.n2806 VGND.n2805 0.2525
R22922 VGND.n2804 VGND.n2803 0.2525
R22923 VGND.n2802 VGND.n2801 0.2525
R22924 VGND.n2800 VGND.n2799 0.2525
R22925 VGND.n2798 VGND.n2797 0.2525
R22926 VGND.n2792 VGND.n2791 0.2525
R22927 VGND.n2790 VGND.n2789 0.2525
R22928 VGND.n2785 VGND.n2784 0.2525
R22929 VGND.n2783 VGND.n2782 0.2525
R22930 VGND.n2781 VGND.n2780 0.2525
R22931 VGND.n2779 VGND.n2778 0.2525
R22932 VGND.n2626 VGND.n2625 0.2525
R22933 VGND.n2727 VGND.n2726 0.2525
R22934 VGND.n2723 VGND.n2722 0.2525
R22935 VGND.n2721 VGND.n2720 0.2525
R22936 VGND.n2718 VGND 0.2525
R22937 VGND.n2713 VGND.n2712 0.2525
R22938 VGND.n2711 VGND.n2710 0.2525
R22939 VGND.n2709 VGND.n2708 0.2525
R22940 VGND.n2705 VGND.n2704 0.2525
R22941 VGND.n2703 VGND.n2702 0.2525
R22942 VGND.n2701 VGND.n2700 0.2525
R22943 VGND.n2697 VGND.n2696 0.2525
R22944 VGND.n2695 VGND.n2694 0.2525
R22945 VGND.n2690 VGND.n2689 0.2525
R22946 VGND.n2688 VGND.n2687 0.2525
R22947 VGND.n2686 VGND.n2685 0.2525
R22948 VGND.n2684 VGND.n2683 0.2525
R22949 VGND.n2679 VGND.n2678 0.2525
R22950 VGND.n2677 VGND.n2676 0.2525
R22951 VGND.n2675 VGND.n2674 0.2525
R22952 VGND.n2673 VGND.n2672 0.2525
R22953 VGND.n2671 VGND.n2670 0.2525
R22954 VGND.n2669 VGND.n2668 0.2525
R22955 VGND.n2667 VGND.n2666 0.2525
R22956 VGND.n2665 VGND.n2664 0.2525
R22957 VGND.n2660 VGND.n2659 0.2525
R22958 VGND.n2658 VGND.n2657 0.2525
R22959 VGND.n2651 VGND.n2650 0.2525
R22960 VGND.n2649 VGND.n2648 0.2525
R22961 VGND.n2647 VGND.n2646 0.2525
R22962 VGND.n431 VGND.n430 0.2525
R22963 VGND.n433 VGND.n432 0.2525
R22964 VGND.n438 VGND.n437 0.2525
R22965 VGND.n2424 VGND.n2423 0.2525
R22966 VGND.n2422 VGND.n2421 0.2525
R22967 VGND.n2420 VGND.n2419 0.2525
R22968 VGND.n2416 VGND.n2415 0.2525
R22969 VGND.n489 VGND.n488 0.2525
R22970 VGND.n2362 VGND 0.2525
R22971 VGND.n2355 VGND.n2354 0.2525
R22972 VGND.n544 VGND.n543 0.2525
R22973 VGND.n424 VGND.n423 0.2525
R22974 VGND.n422 VGND.n421 0.2525
R22975 VGND.n2485 VGND.n2484 0.2525
R22976 VGND.n2481 VGND.n2480 0.2525
R22977 VGND.n2479 VGND.n2478 0.2525
R22978 VGND.n2477 VGND.n2476 0.2525
R22979 VGND.n2475 VGND.n2474 0.2525
R22980 VGND.n2471 VGND.n2470 0.2525
R22981 VGND.n2469 VGND.n2468 0.2525
R22982 VGND.n2467 VGND.n2466 0.2525
R22983 VGND.n2251 VGND.n2250 0.2525
R22984 VGND.n2253 VGND.n2252 0.2525
R22985 VGND.n2255 VGND.n2254 0.2525
R22986 VGND.n2259 VGND.n2258 0.2525
R22987 VGND.n2264 VGND.n2263 0.2525
R22988 VGND.n2270 VGND.n2269 0.2525
R22989 VGND.n2272 VGND.n2271 0.2525
R22990 VGND.n2274 VGND.n2273 0.2525
R22991 VGND.n2276 VGND.n2275 0.2525
R22992 VGND.n2278 VGND.n2277 0.2525
R22993 VGND.n2280 VGND.n2279 0.2525
R22994 VGND.n2282 VGND.n2281 0.2525
R22995 VGND.n2288 VGND.n2287 0.2525
R22996 VGND.n2290 VGND.n2289 0.2525
R22997 VGND.n2292 VGND.n2291 0.2525
R22998 VGND.n2294 VGND.n2293 0.2525
R22999 VGND.n2296 VGND.n2295 0.2525
R23000 VGND.n2299 VGND.n2298 0.2525
R23001 VGND.n2301 VGND.n2300 0.2525
R23002 VGND.n2307 VGND.n2306 0.2525
R23003 VGND.n2309 VGND.n2308 0.2525
R23004 VGND.n2311 VGND.n2310 0.2525
R23005 VGND.n2313 VGND.n2312 0.2525
R23006 VGND.n2315 VGND.n2314 0.2525
R23007 VGND.n2317 VGND.n2316 0.2525
R23008 VGND.n2319 VGND.n2318 0.2525
R23009 VGND.n2328 VGND.n2327 0.2525
R23010 VGND.n2326 VGND.n2325 0.2525
R23011 VGND.n2324 VGND.n2323 0.2525
R23012 VGND.n2322 VGND.n2321 0.2525
R23013 VGND.n2347 VGND.n2346 0.2525
R23014 VGND.n2345 VGND.n2344 0.2525
R23015 VGND.n2074 VGND.n2073 0.2525
R23016 VGND.n2156 VGND.n2155 0.2525
R23017 VGND.n2154 VGND.n2153 0.2525
R23018 VGND.n2152 VGND.n2151 0.2525
R23019 VGND.n2148 VGND.n2147 0.2525
R23020 VGND.n2146 VGND.n2145 0.2525
R23021 VGND.n2144 VGND.n2143 0.2525
R23022 VGND.n2140 VGND.n2139 0.2525
R23023 VGND.n2138 VGND.n2137 0.2525
R23024 VGND.n2136 VGND.n2135 0.2525
R23025 VGND.n2134 VGND.n2133 0.2525
R23026 VGND.n2131 VGND.n2130 0.2525
R23027 VGND.n2129 VGND.n2128 0.2525
R23028 VGND.n2127 VGND.n2126 0.2525
R23029 VGND.n2122 VGND.n2121 0.2525
R23030 VGND.n2120 VGND.n2119 0.2525
R23031 VGND.n2118 VGND.n2117 0.2525
R23032 VGND.n2116 VGND.n2115 0.2525
R23033 VGND.n2114 VGND.n2113 0.2525
R23034 VGND.n2112 VGND.n2111 0.2525
R23035 VGND.n2110 VGND.n2109 0.2525
R23036 VGND.n2108 VGND.n2107 0.2525
R23037 VGND.n2103 VGND.n2102 0.2525
R23038 VGND.n2101 VGND.n2100 0.2525
R23039 VGND.n2099 VGND.n2098 0.2525
R23040 VGND.n3341 VGND.n3340 0.2525
R23041 VGND.n3343 VGND.n3342 0.2525
R23042 VGND.n3345 VGND.n3344 0.2525
R23043 VGND.n2079 VGND.n2078 0.25025
R23044 VGND.n3422 VGND.n3421 0.2495
R23045 VGND.n1546 VGND.n1545 0.2495
R23046 VGND.n2204 VGND 0.2495
R23047 VGND VGND.n2370 0.2495
R23048 VGND.n2353 VGND.n2352 0.2495
R23049 VGND.n2349 VGND.n2222 0.2495
R23050 VGND VGND.n873 0.24875
R23051 VGND.n1620 VGND.n1619 0.248
R23052 VGND.n219 VGND.n218 0.2465
R23053 VGND.n1817 VGND.n1816 0.24275
R23054 VGND.n173 VGND 0.2405
R23055 VGND.n1570 VGND.n1569 0.2405
R23056 VGND VGND.n1601 0.2405
R23057 VGND.n1455 VGND 0.2405
R23058 VGND.n1968 VGND 0.2405
R23059 VGND.n2413 VGND.n468 0.2405
R23060 VGND.n2262 VGND.n2261 0.2405
R23061 VGND.n3107 VGND.n3106 0.2405
R23062 VGND.n824 VGND.n823 0.23975
R23063 VGND.n860 VGND 0.23975
R23064 VGND.t1138 VGND.t4150 0.238924
R23065 VGND.t6793 VGND.t1138 0.238924
R23066 VGND.n86 VGND 0.23825
R23067 VGND VGND.n1533 0.23825
R23068 VGND.n2182 VGND 0.23825
R23069 VGND.n2189 VGND 0.23825
R23070 VGND VGND.n518 0.23825
R23071 VGND.n323 VGND.n322 0.2375
R23072 VGND.n1873 VGND.n1872 0.2375
R23073 VGND.n1222 VGND 0.236
R23074 VGND.n763 VGND 0.2345
R23075 VGND.n1843 VGND.n1842 0.2345
R23076 VGND.n1975 VGND 0.2345
R23077 VGND.n686 VGND.n685 0.2345
R23078 VGND.n3254 VGND.n3253 0.2345
R23079 VGND.n1751 VGND 0.23075
R23080 VGND.n2827 VGND.n410 0.23
R23081 VGND.n2824 VGND.n412 0.23
R23082 VGND.n2693 VGND.n2692 0.23
R23083 VGND.n1406 VGND.n1405 0.2285
R23084 VGND.n327 VGND.n326 0.2285
R23085 VGND.n1538 VGND.n1537 0.2285
R23086 VGND.n3396 VGND 0.2285
R23087 VGND.n1737 VGND.n1736 0.2285
R23088 VGND.n1990 VGND.n1989 0.2285
R23089 VGND.n1904 VGND.n1903 0.2285
R23090 VGND.n2379 VGND.n2378 0.2285
R23091 VGND.n2361 VGND.n2360 0.2285
R23092 VGND.n3427 VGND.n3426 0.2255
R23093 VGND.n517 VGND.n516 0.2255
R23094 VGND.n3411 VGND.n3410 0.224
R23095 VGND VGND.n834 0.2225
R23096 VGND.n127 VGND 0.2225
R23097 VGND VGND.n216 0.2225
R23098 VGND VGND.n82 0.2225
R23099 VGND.n1548 VGND 0.2225
R23100 VGND.n3382 VGND 0.2225
R23101 VGND VGND.n1676 0.2225
R23102 VGND VGND.n1950 0.2225
R23103 VGND VGND.n755 0.2225
R23104 VGND.n1916 VGND 0.2225
R23105 VGND.n2441 VGND 0.2225
R23106 VGND.n2501 VGND 0.2225
R23107 VGND.n2167 VGND.n550 0.2225
R23108 VGND VGND.n3058 0.2225
R23109 VGND VGND.n3163 0.2225
R23110 VGND VGND.n3292 0.2225
R23111 VGND.n1762 VGND.n1761 0.221
R23112 VGND.n1871 VGND 0.221
R23113 VGND.n3276 VGND.n3275 0.221
R23114 VGND.n3272 VGND.n3271 0.221
R23115 VGND.n311 VGND 0.22025
R23116 VGND VGND.n1512 0.22025
R23117 VGND.n757 VGND 0.22025
R23118 VGND VGND.n2037 0.22025
R23119 VGND.n1415 VGND.n1414 0.2195
R23120 VGND.n3692 VGND.n3691 0.2195
R23121 VGND.n2530 VGND.n2529 0.2195
R23122 VGND.n1017 VGND.n1015 0.2195
R23123 VGND VGND.n2179 0.21575
R23124 VGND.n3144 VGND.n371 0.215
R23125 VGND VGND.n745 0.2105
R23126 VGND.n2405 VGND 0.2105
R23127 VGND VGND.n2398 0.2105
R23128 VGND.n2886 VGND 0.20975
R23129 VGND VGND.n2066 0.209
R23130 VGND VGND.n748 0.20825
R23131 VGND.n1480 VGND 0.2075
R23132 VGND.n1763 VGND 0.2075
R23133 VGND VGND.n2050 0.2075
R23134 VGND.n861 VGND.n860 0.206
R23135 VGND.n1210 VGND 0.2045
R23136 VGND.n1740 VGND.n1739 0.2045
R23137 VGND.n1933 VGND.n1932 0.2045
R23138 VGND.n951 VGND.n950 0.2045
R23139 VGND.n2198 VGND.n2169 0.2045
R23140 VGND VGND.n2367 0.2045
R23141 VGND.n1393 VGND.n1392 0.2015
R23142 VGND VGND.n1385 0.2015
R23143 VGND.n2407 VGND.n2406 0.2015
R23144 VGND.n2036 VGND.n2035 0.2015
R23145 VGND.n1263 VGND 0.2
R23146 VGND.n1093 VGND 0.2
R23147 VGND.n1079 VGND 0.2
R23148 VGND VGND.n426 0.2
R23149 VGND VGND.n3671 0.1985
R23150 VGND.n3484 VGND 0.1985
R23151 VGND.n3636 VGND 0.1985
R23152 VGND.n3651 VGND 0.1985
R23153 VGND.n3467 VGND 0.1985
R23154 VGND VGND.n3573 0.1985
R23155 VGND VGND.n3605 0.1985
R23156 VGND VGND.n3621 0.1985
R23157 VGND VGND.n3589 0.1985
R23158 VGND VGND.n3557 0.1985
R23159 VGND.n3541 VGND 0.1985
R23160 VGND VGND.n3702 0.1985
R23161 VGND.n23 VGND 0.1985
R23162 VGND.n3496 VGND 0.1985
R23163 VGND.n3511 VGND 0.1985
R23164 VGND.n3526 VGND 0.1985
R23165 VGND.n915 VGND 0.1985
R23166 VGND.n932 VGND 0.1985
R23167 VGND VGND.n812 0.1985
R23168 VGND.n863 VGND 0.1985
R23169 VGND.n1404 VGND.n59 0.1985
R23170 VGND VGND.n3441 0.1985
R23171 VGND.n3440 VGND 0.1985
R23172 VGND.n3434 VGND 0.1985
R23173 VGND VGND.n132 0.1985
R23174 VGND.n131 VGND 0.1985
R23175 VGND VGND.n167 0.1985
R23176 VGND.n175 VGND 0.1985
R23177 VGND VGND.n185 0.1985
R23178 VGND VGND.n226 0.1985
R23179 VGND.n79 VGND 0.1985
R23180 VGND.n88 VGND 0.1985
R23181 VGND VGND.n106 0.1985
R23182 VGND.n1295 VGND 0.1985
R23183 VGND VGND.n1331 0.1985
R23184 VGND.n1334 VGND 0.1985
R23185 VGND.n1343 VGND 0.1985
R23186 VGND.n1341 VGND 0.1985
R23187 VGND VGND.n291 0.1985
R23188 VGND VGND.n294 0.1985
R23189 VGND VGND.n324 0.1985
R23190 VGND VGND.n1243 0.1985
R23191 VGND.n1242 VGND 0.1985
R23192 VGND.n1272 VGND 0.1985
R23193 VGND VGND.n1259 0.1985
R23194 VGND.n1622 VGND 0.1985
R23195 VGND VGND.n1615 0.1985
R23196 VGND VGND.n1453 0.1985
R23197 VGND.n1542 VGND 0.1985
R23198 VGND VGND.n1517 0.1985
R23199 VGND.n1510 VGND.n1509 0.1985
R23200 VGND VGND.n1227 0.1985
R23201 VGND.n1226 VGND 0.1985
R23202 VGND.n1637 VGND 0.1985
R23203 VGND VGND.n1642 0.1985
R23204 VGND VGND.n1679 0.1985
R23205 VGND VGND.n1695 0.1985
R23206 VGND.n1783 VGND.n1782 0.1985
R23207 VGND.n1758 VGND 0.1985
R23208 VGND VGND.n3371 0.1985
R23209 VGND VGND.n1185 0.1985
R23210 VGND VGND.n1177 0.1985
R23211 VGND VGND.n1166 0.1985
R23212 VGND VGND.n1139 0.1985
R23213 VGND VGND.n590 0.1985
R23214 VGND.n1802 VGND 0.1985
R23215 VGND.n1095 VGND 0.1985
R23216 VGND VGND.n1999 0.1985
R23217 VGND.n1931 VGND.n1930 0.1985
R23218 VGND.n1908 VGND 0.1985
R23219 VGND VGND.n1893 0.1985
R23220 VGND VGND.n960 0.1985
R23221 VGND VGND.n2205 0.1985
R23222 VGND.n465 VGND.n464 0.1985
R23223 VGND VGND.n2436 0.1985
R23224 VGND.n2365 VGND 0.1985
R23225 VGND VGND.n545 0.1985
R23226 VGND VGND.n2229 0.1985
R23227 VGND.n2245 VGND 0.1985
R23228 VGND.n2552 VGND.n2551 0.1985
R23229 VGND.n2532 VGND 0.1985
R23230 VGND VGND.n2527 0.1985
R23231 VGND.n2504 VGND.n2503 0.1985
R23232 VGND.n2892 VGND.n2891 0.1985
R23233 VGND.n1019 VGND 0.1985
R23234 VGND VGND.n1064 0.1985
R23235 VGND.n1041 VGND 0.1985
R23236 VGND.n2043 VGND 0.1985
R23237 VGND.n2986 VGND.n2985 0.1985
R23238 VGND.n3048 VGND.n3047 0.1985
R23239 VGND.n3073 VGND.n3072 0.1985
R23240 VGND.n3091 VGND.n3090 0.1985
R23241 VGND.n3151 VGND.n3150 0.1985
R23242 VGND.n3179 VGND.n3178 0.1985
R23243 VGND.n3196 VGND.n3195 0.1985
R23244 VGND.n3278 VGND.n3277 0.1985
R23245 VGND.n3309 VGND.n3308 0.1985
R23246 VGND.n3324 VGND.n3323 0.1985
R23247 VGND.n3753 VGND.n3752 0.1985
R23248 VGND VGND.n1860 0.19775
R23249 VGND.n1924 VGND 0.19775
R23250 VGND VGND.n2597 0.19775
R23251 VGND.n2734 VGND 0.19775
R23252 VGND VGND.n2724 0.19775
R23253 VGND VGND.n2706 0.19775
R23254 VGND VGND.n2652 0.19775
R23255 VGND VGND.n2417 0.19775
R23256 VGND VGND.n2472 0.19775
R23257 VGND.n2257 VGND 0.19775
R23258 VGND VGND.n2149 0.19775
R23259 VGND.n1390 VGND.n1389 0.197
R23260 VGND.n921 VGND.n920 0.1955
R23261 VGND.n3449 VGND.n3448 0.1955
R23262 VGND.n1572 VGND.n1571 0.1955
R23263 VGND.n1278 VGND 0.1955
R23264 VGND.n3402 VGND.n3401 0.1955
R23265 VGND.n1669 VGND.n1668 0.1955
R23266 VGND.n1698 VGND 0.1955
R23267 VGND.n1789 VGND.n1788 0.1955
R23268 VGND.n2621 VGND.n2614 0.1955
R23269 VGND.n2610 VGND.n2603 0.1955
R23270 VGND.n393 VGND.n392 0.1955
R23271 VGND.n2961 VGND.n385 0.1955
R23272 VGND.n2729 VGND.n2623 0.1955
R23273 VGND.n2912 VGND.n2911 0.1955
R23274 VGND.n2049 VGND.n2048 0.1955
R23275 VGND.n3001 VGND.n383 0.1955
R23276 VGND.n3413 VGND.n3412 0.19475
R23277 VGND.n911 VGND 0.194
R23278 VGND.n2450 VGND 0.194
R23279 VGND VGND.n2005 0.194
R23280 VGND.n221 VGND 0.1925
R23281 VGND VGND.n3689 0.1925
R23282 VGND VGND.n1253 0.1925
R23283 VGND.n1610 VGND.n1609 0.1925
R23284 VGND VGND.n1605 0.1925
R23285 VGND VGND.n1555 0.1925
R23286 VGND VGND.n3404 0.1925
R23287 VGND.n1224 VGND.n1223 0.1925
R23288 VGND.n1214 VGND.n1213 0.1925
R23289 VGND.n1634 VGND 0.1925
R23290 VGND.n1682 VGND.n1681 0.1925
R23291 VGND VGND.n587 0.1925
R23292 VGND.n644 VGND.n643 0.1925
R23293 VGND VGND.n2444 0.1925
R23294 VGND.n493 VGND 0.1925
R23295 VGND.n2515 VGND 0.1925
R23296 VGND VGND.n2968 0.1925
R23297 VGND.n755 VGND.n754 0.19175
R23298 VGND.t1077 VGND.t146 0.191239
R23299 VGND.n1442 VGND.n1420 0.191
R23300 VGND VGND.n742 0.19025
R23301 VGND.n1524 VGND.n1523 0.1895
R23302 VGND VGND.n815 0.18875
R23303 VGND VGND.n1244 0.188
R23304 VGND VGND.n1121 0.188
R23305 VGND VGND.n1179 0.188
R23306 VGND VGND.n1141 0.188
R23307 VGND VGND.n996 0.188
R23308 VGND VGND.n976 0.188
R23309 VGND.n913 VGND.n912 0.18725
R23310 VGND.n3380 VGND.n208 0.1865
R23311 VGND.n1688 VGND 0.1835
R23312 VGND VGND.n614 0.1835
R23313 VGND VGND.n66 0.18275
R23314 VGND VGND.n91 0.18275
R23315 VGND.n103 VGND 0.18275
R23316 VGND VGND.n1705 0.18275
R23317 VGND VGND.n1803 0.18275
R23318 VGND.n1560 VGND.n1559 0.182
R23319 VGND.n1568 VGND 0.1805
R23320 VGND.n315 VGND 0.1805
R23321 VGND VGND.n1466 0.1805
R23322 VGND VGND.n1468 0.1805
R23323 VGND.n1541 VGND.n1540 0.1805
R23324 VGND.n1505 VGND 0.1805
R23325 VGND.n1679 VGND 0.1805
R23326 VGND VGND.n752 0.1805
R23327 VGND.n642 VGND 0.1805
R23328 VGND.n954 VGND.n953 0.1805
R23329 VGND.n2395 VGND.n2394 0.1805
R23330 VGND.n2883 VGND.n409 0.1805
R23331 VGND.n2788 VGND.n2787 0.1805
R23332 VGND.n2166 VGND.n2165 0.1805
R23333 VGND.n1459 VGND.n1458 0.1775
R23334 VGND.n2406 VGND.n2405 0.1775
R23335 VGND.n240 VGND 0.1745
R23336 VGND VGND.n81 0.1745
R23337 VGND VGND.n1289 0.1745
R23338 VGND.n296 VGND.n295 0.1745
R23339 VGND VGND.n318 0.1745
R23340 VGND.n1526 VGND 0.1745
R23341 VGND.n254 VGND.n253 0.1745
R23342 VGND.n1573 VGND.n1572 0.1715
R23343 VGND.n1381 VGND.n1380 0.1715
R23344 VGND.n3428 VGND.n3427 0.1715
R23345 VGND.n324 VGND.n323 0.1715
R23346 VGND.n1457 VGND.n1456 0.1715
R23347 VGND VGND.n1508 0.1715
R23348 VGND.n1506 VGND.n1505 0.1715
R23349 VGND.n1655 VGND.n1654 0.1715
R23350 VGND.n1964 VGND.n1963 0.1715
R23351 VGND.n1795 VGND.n1794 0.1715
R23352 VGND.n643 VGND.n642 0.1715
R23353 VGND.n2935 VGND.n2934 0.1715
R23354 VGND.n2410 VGND 0.17075
R23355 VGND VGND.n853 0.17
R23356 VGND VGND.n3446 0.17
R23357 VGND VGND.n1459 0.17
R23358 VGND.n1586 VGND.n1585 0.16925
R23359 VGND.n3450 VGND.n3449 0.1685
R23360 VGND.n129 VGND.n128 0.1685
R23361 VGND.n235 VGND.n234 0.1685
R23362 VGND.n234 VGND.n233 0.1685
R23363 VGND.n68 VGND.n67 0.1685
R23364 VGND.n70 VGND.n69 0.1685
R23365 VGND.n102 VGND.n101 0.1685
R23366 VGND.n101 VGND.n100 0.1685
R23367 VGND.n100 VGND.n99 0.1685
R23368 VGND.n98 VGND.n97 0.1685
R23369 VGND.n97 VGND.n96 0.1685
R23370 VGND.n96 VGND.n54 0.1685
R23371 VGND.n1325 VGND.n1324 0.1685
R23372 VGND.n1328 VGND.n1327 0.1685
R23373 VGND.n1330 VGND.n1329 0.1685
R23374 VGND.n1569 VGND.n1568 0.1685
R23375 VGND.n3689 VGND.n3688 0.1685
R23376 VGND.n1252 VGND.n1251 0.1685
R23377 VGND VGND.n1472 0.1685
R23378 VGND.n1520 VGND.n1519 0.1685
R23379 VGND.n3404 VGND.n3403 0.1685
R23380 VGND.n1231 VGND 0.1685
R23381 VGND.n1668 VGND.n1667 0.1685
R23382 VGND.n1735 VGND.n1734 0.1685
R23383 VGND.n752 VGND.n751 0.1685
R23384 VGND.n1089 VGND.n1088 0.1685
R23385 VGND.n1993 VGND 0.1685
R23386 VGND.n1902 VGND.n1901 0.1685
R23387 VGND.n2391 VGND.n2390 0.1685
R23388 VGND.n2193 VGND.n2192 0.1685
R23389 VGND.n495 VGND.n494 0.1685
R23390 VGND.n496 VGND.n495 0.1685
R23391 VGND.n497 VGND.n496 0.1685
R23392 VGND.n498 VGND.n497 0.1685
R23393 VGND.n499 VGND.n498 0.1685
R23394 VGND.n500 VGND.n499 0.1685
R23395 VGND.n501 VGND.n500 0.1685
R23396 VGND.n502 VGND.n501 0.1685
R23397 VGND.n504 VGND.n503 0.1685
R23398 VGND.n505 VGND.n504 0.1685
R23399 VGND.n506 VGND.n505 0.1685
R23400 VGND.n507 VGND.n506 0.1685
R23401 VGND.n2359 VGND.n2358 0.1685
R23402 VGND.n2550 VGND.n2549 0.1685
R23403 VGND.n2549 VGND.n2548 0.1685
R23404 VGND.n2548 VGND.n2547 0.1685
R23405 VGND.n2547 VGND.n2546 0.1685
R23406 VGND.n2546 VGND.n2545 0.1685
R23407 VGND.n2545 VGND.n2544 0.1685
R23408 VGND.n2543 VGND.n2542 0.1685
R23409 VGND.n2542 VGND.n2541 0.1685
R23410 VGND.n2541 VGND.n2540 0.1685
R23411 VGND.n2540 VGND.n2539 0.1685
R23412 VGND.n2539 VGND.n2538 0.1685
R23413 VGND.n2538 VGND.n2537 0.1685
R23414 VGND.n2537 VGND.n2536 0.1685
R23415 VGND.n2893 VGND.n2892 0.1685
R23416 VGND.n2894 VGND.n2893 0.1685
R23417 VGND.n2896 VGND.n2895 0.1685
R23418 VGND.n2897 VGND.n2896 0.1685
R23419 VGND.n2898 VGND.n2897 0.1685
R23420 VGND.n2899 VGND.n2898 0.1685
R23421 VGND.n2901 VGND.n2900 0.1685
R23422 VGND.n2902 VGND.n2901 0.1685
R23423 VGND.n2903 VGND.n2902 0.1685
R23424 VGND.n2904 VGND.n2903 0.1685
R23425 VGND.n2905 VGND.n2904 0.1685
R23426 VGND.n2906 VGND.n2905 0.1685
R23427 VGND.n2907 VGND.n2906 0.1685
R23428 VGND.n2024 VGND.n2023 0.1685
R23429 VGND.n2025 VGND.n2024 0.1685
R23430 VGND.n2026 VGND.n2025 0.1685
R23431 VGND.n2029 VGND.n2028 0.1685
R23432 VGND.n2030 VGND.n2029 0.1685
R23433 VGND.n2058 VGND 0.1685
R23434 VGND.n2966 VGND.n2965 0.1685
R23435 VGND.n2965 VGND.n2964 0.1685
R23436 VGND.n2964 VGND.n2963 0.1685
R23437 VGND.n2996 VGND.n2995 0.1685
R23438 VGND.n2995 VGND.n2994 0.1685
R23439 VGND.n2994 VGND.n2993 0.1685
R23440 VGND.n2984 VGND.n2983 0.1685
R23441 VGND.n2983 VGND.n2982 0.1685
R23442 VGND.n2982 VGND.n2981 0.1685
R23443 VGND.n2981 VGND.n2980 0.1685
R23444 VGND.n2980 VGND.n2979 0.1685
R23445 VGND.n3049 VGND.n3048 0.1685
R23446 VGND.n3050 VGND.n3049 0.1685
R23447 VGND.n3051 VGND.n3050 0.1685
R23448 VGND.n3052 VGND.n3051 0.1685
R23449 VGND.n3053 VGND.n3052 0.1685
R23450 VGND.n3054 VGND.n3053 0.1685
R23451 VGND.n3055 VGND.n3054 0.1685
R23452 VGND.n3072 VGND.n3071 0.1685
R23453 VGND.n3071 VGND.n3070 0.1685
R23454 VGND.n3070 VGND.n3069 0.1685
R23455 VGND.n3069 VGND.n3068 0.1685
R23456 VGND.n3068 VGND.n3067 0.1685
R23457 VGND.n3067 VGND.n3066 0.1685
R23458 VGND.n3066 VGND.n3065 0.1685
R23459 VGND.n3064 VGND.n3063 0.1685
R23460 VGND.n3063 VGND.n3062 0.1685
R23461 VGND.n3102 VGND.n3101 0.1685
R23462 VGND.n3101 VGND.n3100 0.1685
R23463 VGND.n3100 VGND.n3099 0.1685
R23464 VGND.n3089 VGND.n3088 0.1685
R23465 VGND.n3088 VGND.n3087 0.1685
R23466 VGND.n3087 VGND.n3086 0.1685
R23467 VGND.n3152 VGND.n3151 0.1685
R23468 VGND.n3153 VGND.n3152 0.1685
R23469 VGND.n3154 VGND.n3153 0.1685
R23470 VGND.n3155 VGND.n3154 0.1685
R23471 VGND.n3156 VGND.n3155 0.1685
R23472 VGND.n3157 VGND.n3156 0.1685
R23473 VGND.n3158 VGND.n3157 0.1685
R23474 VGND.n3160 VGND.n3159 0.1685
R23475 VGND.n3161 VGND.n3160 0.1685
R23476 VGND.n3178 VGND.n3177 0.1685
R23477 VGND.n3177 VGND.n3176 0.1685
R23478 VGND.n3176 VGND.n3175 0.1685
R23479 VGND.n3175 VGND.n3174 0.1685
R23480 VGND.n3174 VGND.n3173 0.1685
R23481 VGND.n3173 VGND.n3172 0.1685
R23482 VGND.n3172 VGND.n3171 0.1685
R23483 VGND.n3170 VGND.n3169 0.1685
R23484 VGND.n3169 VGND.n3168 0.1685
R23485 VGND.n3168 VGND.n3167 0.1685
R23486 VGND.n3167 VGND.n3166 0.1685
R23487 VGND.n3207 VGND.n3206 0.1685
R23488 VGND.n3206 VGND.n3205 0.1685
R23489 VGND.n3194 VGND.n3193 0.1685
R23490 VGND.n3279 VGND.n3278 0.1685
R23491 VGND.n3280 VGND.n3279 0.1685
R23492 VGND.n3281 VGND.n3280 0.1685
R23493 VGND.n3282 VGND.n3281 0.1685
R23494 VGND.n3283 VGND.n3282 0.1685
R23495 VGND.n3284 VGND.n3283 0.1685
R23496 VGND.n3285 VGND.n3284 0.1685
R23497 VGND.n3287 VGND.n3286 0.1685
R23498 VGND.n3288 VGND.n3287 0.1685
R23499 VGND.n3289 VGND.n3288 0.1685
R23500 VGND.n3290 VGND.n3289 0.1685
R23501 VGND.n3308 VGND.n3307 0.1685
R23502 VGND.n3307 VGND.n3306 0.1685
R23503 VGND.n3306 VGND.n3305 0.1685
R23504 VGND.n3305 VGND.n3304 0.1685
R23505 VGND.n3304 VGND.n3303 0.1685
R23506 VGND.n3303 VGND.n3302 0.1685
R23507 VGND.n3302 VGND.n3301 0.1685
R23508 VGND.n3300 VGND.n3299 0.1685
R23509 VGND.n3299 VGND.n3298 0.1685
R23510 VGND.n3298 VGND.n3297 0.1685
R23511 VGND.n3297 VGND.n3296 0.1685
R23512 VGND.n3296 VGND.n3295 0.1685
R23513 VGND.n3295 VGND.n3294 0.1685
R23514 VGND.n3752 VGND.n3751 0.1685
R23515 VGND.n3751 VGND.n3750 0.1685
R23516 VGND.n3750 VGND.n3749 0.1685
R23517 VGND.n3749 VGND.n3748 0.1685
R23518 VGND.n3748 VGND.n3747 0.1685
R23519 VGND.n3747 VGND.n3746 0.1685
R23520 VGND.n3746 VGND.n3745 0.1685
R23521 VGND.n3744 VGND.n3743 0.1685
R23522 VGND.n3743 VGND.n3742 0.1685
R23523 VGND.n3742 VGND.n3741 0.1685
R23524 VGND.n3741 VGND.n3740 0.1685
R23525 VGND.n3740 VGND.n3739 0.1685
R23526 VGND.n3739 VGND.n3738 0.1685
R23527 VGND.n3734 VGND.n3733 0.1685
R23528 VGND.n3733 VGND.n3732 0.1685
R23529 VGND.n3732 VGND.n3731 0.1685
R23530 VGND.n3731 VGND.n3730 0.1685
R23531 VGND.n3730 VGND.n3729 0.1685
R23532 VGND.n3729 VGND.n3728 0.1685
R23533 VGND.n3728 VGND.n3727 0.1685
R23534 VGND.n3726 VGND.n3725 0.1685
R23535 VGND.n3725 VGND.n3724 0.1685
R23536 VGND.n3724 VGND.n3723 0.1685
R23537 VGND.n3723 VGND.n3722 0.1685
R23538 VGND.n3722 VGND.n3721 0.1685
R23539 VGND.n3721 VGND.n3720 0.1685
R23540 VGND.n3720 VGND.n3719 0.1685
R23541 VGND.n111 VGND 0.167
R23542 VGND.n1395 VGND 0.167
R23543 VGND VGND.n1387 0.167
R23544 VGND.n928 VGND 0.1655
R23545 VGND.n194 VGND 0.1655
R23546 VGND.n1250 VGND.n1249 0.1655
R23547 VGND.n1507 VGND.n1506 0.1655
R23548 VGND.n3398 VGND.n3397 0.1655
R23549 VGND.n1913 VGND.n1912 0.1655
R23550 VGND.n2936 VGND.n2935 0.1655
R23551 VGND.n1512 VGND 0.16475
R23552 VGND.n914 VGND.n913 0.164
R23553 VGND.n1293 VGND.n1292 0.164
R23554 VGND.n1382 VGND 0.164
R23555 VGND.n3417 VGND 0.164
R23556 VGND.n1241 VGND.n1240 0.164
R23557 VGND.n1229 VGND.n1228 0.164
R23558 VGND.n1225 VGND.n1224 0.164
R23559 VGND.n1635 VGND.n1634 0.164
R23560 VGND.n1642 VGND.n1641 0.164
R23561 VGND.n1689 VGND.n1688 0.164
R23562 VGND.n1756 VGND 0.164
R23563 VGND.n1169 VGND.n1168 0.164
R23564 VGND.n1965 VGND 0.164
R23565 VGND.n1110 VGND.n1109 0.164
R23566 VGND.n1100 VGND.n1099 0.164
R23567 VGND.n1091 VGND.n1090 0.164
R23568 VGND.n1937 VGND.n614 0.164
R23569 VGND.n454 VGND.n453 0.164
R23570 VGND.n2438 VGND.n2437 0.164
R23571 VGND.n2460 VGND.n2459 0.164
R23572 VGND.n2454 VGND.n2453 0.164
R23573 VGND.n1039 VGND.n1038 0.164
R23574 VGND VGND.n3429 0.1625
R23575 VGND.n865 VGND.n864 0.161
R23576 VGND VGND.n2384 0.161
R23577 VGND.n3147 VGND 0.1595
R23578 VGND VGND.n168 0.15875
R23579 VGND.n1583 VGND.n1582 0.15875
R23580 VGND VGND.n292 0.15875
R23581 VGND.n1127 VGND 0.15875
R23582 VGND.n2389 VGND 0.15875
R23583 VGND VGND.n830 0.1565
R23584 VGND VGND.n859 0.1565
R23585 VGND.n124 VGND 0.1565
R23586 VGND.n1298 VGND 0.1565
R23587 VGND.n1577 VGND 0.1565
R23588 VGND VGND.n310 0.1565
R23589 VGND.n1458 VGND 0.1565
R23590 VGND VGND.n1556 0.1565
R23591 VGND VGND.n1548 0.1565
R23592 VGND VGND.n1534 0.1565
R23593 VGND VGND.n1504 0.1565
R23594 VGND VGND.n3395 0.1565
R23595 VGND VGND.n1784 0.1565
R23596 VGND VGND.n1768 0.1565
R23597 VGND.n1960 VGND 0.1565
R23598 VGND VGND.n1959 0.1565
R23599 VGND.n626 VGND 0.1565
R23600 VGND.n638 VGND 0.1565
R23601 VGND VGND.n641 0.1565
R23602 VGND.n1923 VGND 0.1565
R23603 VGND VGND.n1900 0.1565
R23604 VGND VGND.n956 0.1565
R23605 VGND VGND.n2386 0.1565
R23606 VGND.n2386 VGND.n2385 0.1565
R23607 VGND.n2655 VGND.n2654 0.1565
R23608 VGND.n514 VGND.n513 0.1565
R23609 VGND VGND.n2357 0.1565
R23610 VGND VGND.n162 0.15575
R23611 VGND.n225 VGND 0.15575
R23612 VGND VGND.n1300 0.15575
R23613 VGND VGND.n1309 0.15575
R23614 VGND.n1344 VGND 0.15575
R23615 VGND.n1585 VGND 0.15575
R23616 VGND.n3414 VGND 0.15575
R23617 VGND.n1467 VGND 0.15575
R23618 VGND VGND.n1471 0.15575
R23619 VGND.n3384 VGND 0.15575
R23620 VGND.n1691 VGND 0.15575
R23621 VGND VGND.n1692 0.15575
R23622 VGND.n1941 VGND 0.15575
R23623 VGND.n750 VGND 0.15575
R23624 VGND VGND.n2178 0.15575
R23625 VGND VGND.n2053 0.15575
R23626 VGND.n2056 VGND 0.15575
R23627 VGND.n852 VGND 0.15425
R23628 VGND VGND.n134 0.15425
R23629 VGND.n67 VGND 0.15425
R23630 VGND.n92 VGND 0.15425
R23631 VGND VGND.n102 0.15425
R23632 VGND VGND.n1323 0.15425
R23633 VGND.n1277 VGND 0.15425
R23634 VGND VGND.n1643 0.15425
R23635 VGND VGND.n1126 0.15425
R23636 VGND.n747 VGND 0.15425
R23637 VGND.n450 VGND 0.15425
R23638 VGND.n2429 VGND 0.15425
R23639 VGND VGND.n2022 0.15425
R23640 VGND.n1527 VGND 0.1535
R23641 VGND VGND.n1687 0.1535
R23642 VGND.n649 VGND 0.1535
R23643 VGND.n2191 VGND.n2190 0.1535
R23644 VGND.n1317 VGND 0.152
R23645 VGND.n322 VGND 0.1505
R23646 VGND VGND.n1476 0.1505
R23647 VGND.n1797 VGND 0.1505
R23648 VGND VGND.n1162 0.14975
R23649 VGND VGND.n1673 0.14825
R23650 VGND VGND.n1960 0.14825
R23651 VGND.n1982 VGND.n1981 0.1475
R23652 VGND.n815 VGND 0.14675
R23653 VGND.n1299 VGND 0.14675
R23654 VGND.n3412 VGND 0.14675
R23655 VGND VGND.n744 0.14675
R23656 VGND.n635 VGND 0.14675
R23657 VGND.n2394 VGND 0.14675
R23658 VGND.n1152 VGND.n1151 0.146
R23659 VGND.n2001 VGND.n576 0.146
R23660 VGND.n2384 VGND.n482 0.146
R23661 VGND.n754 VGND.n753 0.14525
R23662 VGND.n822 VGND 0.1445
R23663 VGND.n829 VGND 0.1445
R23664 VGND.n3438 VGND.n3437 0.1445
R23665 VGND.n3436 VGND.n3435 0.1445
R23666 VGND.n138 VGND.n137 0.1445
R23667 VGND.n301 VGND.n300 0.1445
R23668 VGND.n1613 VGND.n1612 0.1445
R23669 VGND.n1609 VGND.n1608 0.1445
R23670 VGND.n1464 VGND.n1463 0.1445
R23671 VGND.n1556 VGND 0.1445
R23672 VGND.n1549 VGND 0.1445
R23673 VGND.n3386 VGND.n3385 0.1445
R23674 VGND.n1215 VGND.n1214 0.1445
R23675 VGND.n1213 VGND.n1212 0.1445
R23676 VGND.n1703 VGND.n1702 0.1445
R23677 VGND.n1705 VGND.n1704 0.1445
R23678 VGND VGND.n1710 0.1445
R23679 VGND.n1773 VGND 0.1445
R23680 VGND.n1183 VGND.n1182 0.1445
R23681 VGND.n1985 VGND.n1984 0.1445
R23682 VGND.n1983 VGND.n1982 0.1445
R23683 VGND.n1972 VGND.n587 0.1445
R23684 VGND.n1936 VGND.n1935 0.1445
R23685 VGND.n990 VGND.n989 0.1445
R23686 VGND.n977 VGND 0.1445
R23687 VGND.n2401 VGND 0.1445
R23688 VGND.n2219 VGND.n2218 0.1445
R23689 VGND.n1054 VGND.n1053 0.1445
R23690 VGND.n1038 VGND.n1037 0.1445
R23691 VGND.n2050 VGND.n2049 0.1445
R23692 VGND.n1315 VGND.n1314 0.14375
R23693 VGND.t6400 VGND.t6697 0.143554
R23694 VGND.t3682 VGND.t6409 0.143554
R23695 VGND.t139 VGND.t137 0.143554
R23696 VGND VGND.n914 0.143
R23697 VGND.n923 VGND 0.143
R23698 VGND.n922 VGND 0.143
R23699 VGND.n810 VGND 0.143
R23700 VGND.n813 VGND 0.143
R23701 VGND VGND.n1290 0.143
R23702 VGND VGND.n1291 0.143
R23703 VGND.n1322 VGND 0.143
R23704 VGND.n1244 VGND 0.143
R23705 VGND VGND.n1241 0.143
R23706 VGND VGND.n1277 0.143
R23707 VGND.n1276 VGND 0.143
R23708 VGND VGND.n1617 0.143
R23709 VGND.n1228 VGND 0.143
R23710 VGND VGND.n1225 0.143
R23711 VGND VGND.n1222 0.143
R23712 VGND.n1641 VGND 0.143
R23713 VGND.n1646 VGND 0.143
R23714 VGND VGND.n1116 0.143
R23715 VGND VGND.n1115 0.143
R23716 VGND VGND.n1181 0.143
R23717 VGND.n1175 VGND 0.143
R23718 VGND.n1160 VGND 0.143
R23719 VGND.n1153 VGND 0.143
R23720 VGND.n1073 VGND 0.143
R23721 VGND VGND.n1068 0.143
R23722 VGND VGND.n1108 0.143
R23723 VGND VGND.n1107 0.143
R23724 VGND VGND.n1097 0.143
R23725 VGND.n1090 VGND 0.143
R23726 VGND.n2000 VGND 0.143
R23727 VGND.n1997 VGND 0.143
R23728 VGND VGND.n1996 0.143
R23729 VGND VGND.n980 0.143
R23730 VGND.n974 VGND 0.143
R23731 VGND VGND.n965 0.143
R23732 VGND VGND.n964 0.143
R23733 VGND.n461 VGND 0.143
R23734 VGND VGND.n456 0.143
R23735 VGND VGND.n452 0.143
R23736 VGND VGND.n428 0.143
R23737 VGND.n2437 VGND 0.143
R23738 VGND.n2434 VGND 0.143
R23739 VGND VGND.n2433 0.143
R23740 VGND.n2461 VGND 0.143
R23741 VGND VGND.n2452 0.143
R23742 VGND VGND.n2225 0.143
R23743 VGND.n2525 VGND 0.143
R23744 VGND.n1048 VGND 0.143
R23745 VGND VGND.n1036 0.143
R23746 VGND VGND.n2008 0.143
R23747 VGND VGND.n2015 0.143
R23748 VGND.n2016 VGND 0.143
R23749 VGND.n2021 VGND 0.143
R23750 VGND.n3448 VGND.n3447 0.1415
R23751 VGND.n1391 VGND.n1390 0.1415
R23752 VGND.n299 VGND.n298 0.1415
R23753 VGND.n1532 VGND 0.1415
R23754 VGND.n1514 VGND.n1513 0.1415
R23755 VGND.n1790 VGND.n1789 0.1415
R23756 VGND.n1788 VGND.n1787 0.1415
R23757 VGND VGND.n636 0.1415
R23758 VGND.n1013 VGND.n1012 0.1415
R23759 VGND.n2205 VGND.n2204 0.1415
R23760 VGND.n2621 VGND.n2620 0.1415
R23761 VGND.n2610 VGND.n2609 0.1415
R23762 VGND.n394 VGND.n393 0.1415
R23763 VGND.n2961 VGND.n2960 0.1415
R23764 VGND.n436 VGND.n435 0.1415
R23765 VGND.n2487 VGND.n2486 0.1415
R23766 VGND.n2998 VGND.n2997 0.1415
R23767 VGND.n3002 VGND.n3001 0.1415
R23768 VGND.n1389 VGND.n1388 0.14
R23769 VGND.n1387 VGND.n1386 0.14
R23770 VGND.n1617 VGND.n1616 0.14
R23771 VGND.n1197 VGND.n1196 0.14
R23772 VGND.n1195 VGND.n1194 0.14
R23773 VGND VGND.n1762 0.14
R23774 VGND.n1181 VGND.n1180 0.14
R23775 VGND.n1172 VGND.n1171 0.14
R23776 VGND.n1170 VGND.n1169 0.14
R23777 VGND.n980 VGND.n979 0.14
R23778 VGND.n1036 VGND.n1035 0.14
R23779 VGND.n1029 VGND.n1028 0.14
R23780 VGND.n1027 VGND.n1026 0.14
R23781 VGND VGND.n1344 0.13925
R23782 VGND.n1590 VGND 0.13925
R23783 VGND.n1208 VGND 0.13925
R23784 VGND VGND.n2046 0.13925
R23785 VGND.n3674 VGND 0.1385
R23786 VGND.n3486 VGND 0.1385
R23787 VGND.n3639 VGND 0.1385
R23788 VGND.n3654 VGND 0.1385
R23789 VGND.n3469 VGND 0.1385
R23790 VGND.n3576 VGND 0.1385
R23791 VGND.n3608 VGND 0.1385
R23792 VGND.n3624 VGND 0.1385
R23793 VGND.n3592 VGND 0.1385
R23794 VGND.n3560 VGND 0.1385
R23795 VGND.n3544 VGND 0.1385
R23796 VGND.n3705 VGND 0.1385
R23797 VGND.n25 VGND 0.1385
R23798 VGND.n3499 VGND 0.1385
R23799 VGND.n3514 VGND 0.1385
R23800 VGND.n3529 VGND 0.1385
R23801 VGND.n812 VGND 0.1385
R23802 VGND.n833 VGND.n832 0.1385
R23803 VGND.n831 VGND 0.1385
R23804 VGND VGND.n862 0.1385
R23805 VGND VGND.n1417 0.1385
R23806 VGND VGND.n3450 0.1385
R23807 VGND VGND.n3439 0.1385
R23808 VGND.n3437 VGND 0.1385
R23809 VGND VGND.n138 0.1385
R23810 VGND.n167 VGND.n166 0.1385
R23811 VGND.n168 VGND 0.1385
R23812 VGND VGND.n174 0.1385
R23813 VGND.n3453 VGND 0.1385
R23814 VGND VGND.n1294 0.1385
R23815 VGND VGND.n1326 0.1385
R23816 VGND.n1347 VGND.n1346 0.1385
R23817 VGND.n291 VGND.n290 0.1385
R23818 VGND.n295 VGND 0.1385
R23819 VGND.n300 VGND 0.1385
R23820 VGND.n44 VGND 0.1385
R23821 VGND.n1262 VGND 0.1385
R23822 VGND.n1625 VGND.n1624 0.1385
R23823 VGND VGND.n1611 0.1385
R23824 VGND.n1465 VGND 0.1385
R23825 VGND VGND.n1541 0.1385
R23826 VGND VGND.n1527 0.1385
R23827 VGND.n1509 VGND 0.1385
R23828 VGND VGND.n269 0.1385
R23829 VGND VGND.n799 0.1385
R23830 VGND.n1640 VGND.n1639 0.1385
R23831 VGND VGND.n1645 0.1385
R23832 VGND VGND.n1708 0.1385
R23833 VGND.n1774 VGND.n1773 0.1385
R23834 VGND VGND.n1757 0.1385
R23835 VGND.n3377 VGND 0.1385
R23836 VGND.n3360 VGND 0.1385
R23837 VGND VGND.n1183 0.1385
R23838 VGND.n1161 VGND 0.1385
R23839 VGND.n1147 VGND 0.1385
R23840 VGND VGND.n1127 0.1385
R23841 VGND.n1869 VGND 0.1385
R23842 VGND.n1824 VGND 0.1385
R23843 VGND.n1074 VGND 0.1385
R23844 VGND.n1098 VGND 0.1385
R23845 VGND VGND.n1923 0.1385
R23846 VGND.n1917 VGND 0.1385
R23847 VGND VGND.n1907 0.1385
R23848 VGND.n667 VGND 0.1385
R23849 VGND.n975 VGND 0.1385
R23850 VGND.n971 VGND 0.1385
R23851 VGND VGND.n968 0.1385
R23852 VGND.n2208 VGND 0.1385
R23853 VGND.n2863 VGND 0.1385
R23854 VGND.n2615 VGND 0.1385
R23855 VGND.n2604 VGND 0.1385
R23856 VGND VGND.n399 0.1385
R23857 VGND.n2955 VGND 0.1385
R23858 VGND.n2767 VGND 0.1385
R23859 VGND.n2635 VGND 0.1385
R23860 VGND.n462 VGND 0.1385
R23861 VGND VGND.n455 0.1385
R23862 VGND VGND.n451 0.1385
R23863 VGND.n2426 VGND 0.1385
R23864 VGND VGND.n2364 0.1385
R23865 VGND.n532 VGND 0.1385
R23866 VGND VGND.n2451 0.1385
R23867 VGND VGND.n2242 0.1385
R23868 VGND VGND.n2248 0.1385
R23869 VGND.n2333 VGND 0.1385
R23870 VGND VGND.n2910 0.1385
R23871 VGND.n2923 VGND 0.1385
R23872 VGND.n2020 VGND.n2019 0.1385
R23873 VGND.n2047 VGND 0.1385
R23874 VGND VGND.n3356 0.1385
R23875 VGND.n9 VGND 0.1385
R23876 VGND.n3778 VGND 0.1385
R23877 VGND.n3670 VGND 0.137
R23878 VGND VGND.n3485 0.137
R23879 VGND VGND.n3637 0.137
R23880 VGND VGND.n3652 0.137
R23881 VGND VGND.n3468 0.137
R23882 VGND.n3572 VGND 0.137
R23883 VGND.n3604 VGND 0.137
R23884 VGND.n3620 VGND 0.137
R23885 VGND.n3588 VGND 0.137
R23886 VGND.n3556 VGND 0.137
R23887 VGND VGND.n3542 0.137
R23888 VGND.n3701 VGND 0.137
R23889 VGND VGND.n24 0.137
R23890 VGND VGND.n3497 0.137
R23891 VGND VGND.n3512 0.137
R23892 VGND VGND.n3527 0.137
R23893 VGND.n920 VGND 0.137
R23894 VGND VGND.n857 0.137
R23895 VGND.n872 VGND 0.137
R23896 VGND VGND.n1408 0.137
R23897 VGND.n137 VGND 0.137
R23898 VGND.n229 VGND 0.137
R23899 VGND.n347 VGND 0.137
R23900 VGND.n1256 VGND 0.137
R23901 VGND.n1608 VGND 0.137
R23902 VGND VGND.n1455 0.137
R23903 VGND.n1555 VGND 0.137
R23904 VGND.n3407 VGND.n3406 0.137
R23905 VGND VGND.n1230 0.137
R23906 VGND.n1218 VGND 0.137
R23907 VGND VGND.n1653 0.137
R23908 VGND VGND.n1683 0.137
R23909 VGND.n1784 VGND 0.137
R23910 VGND.n1770 VGND 0.137
R23911 VGND.n3370 VGND 0.137
R23912 VGND.n1144 VGND 0.137
R23913 VGND.n1131 VGND 0.137
R23914 VGND VGND.n1798 0.137
R23915 VGND VGND.n1812 0.137
R23916 VGND.n1853 VGND 0.137
R23917 VGND.n1834 VGND 0.137
R23918 VGND.n1088 VGND 0.137
R23919 VGND VGND.n1079 0.137
R23920 VGND VGND.n1992 0.137
R23921 VGND VGND.n628 0.137
R23922 VGND.n1890 VGND 0.137
R23923 VGND.n714 VGND 0.137
R23924 VGND.n696 VGND 0.137
R23925 VGND.n677 VGND 0.137
R23926 VGND.n1009 VGND 0.137
R23927 VGND.n999 VGND 0.137
R23928 VGND.n959 VGND 0.137
R23929 VGND VGND.n2193 0.137
R23930 VGND.n2217 VGND 0.137
R23931 VGND.n2590 VGND 0.137
R23932 VGND.n2572 VGND 0.137
R23933 VGND VGND.n2837 0.137
R23934 VGND VGND.n2855 0.137
R23935 VGND.n2873 VGND 0.137
R23936 VGND VGND.n2741 0.137
R23937 VGND VGND.n2759 0.137
R23938 VGND.n2814 VGND 0.137
R23939 VGND.n2796 VGND 0.137
R23940 VGND.n2777 VGND 0.137
R23941 VGND.n2699 VGND 0.137
R23942 VGND.n2682 VGND 0.137
R23943 VGND.n2680 VGND 0.137
R23944 VGND VGND.n439 0.137
R23945 VGND VGND.n449 0.137
R23946 VGND.n2443 VGND 0.137
R23947 VGND VGND.n490 0.137
R23948 VGND VGND.n507 0.137
R23949 VGND.n542 VGND 0.137
R23950 VGND.n2483 VGND 0.137
R23951 VGND.n2465 VGND 0.137
R23952 VGND VGND.n2226 0.137
R23953 VGND.n2241 VGND 0.137
R23954 VGND VGND.n2246 0.137
R23955 VGND VGND.n2265 0.137
R23956 VGND VGND.n2283 0.137
R23957 VGND VGND.n2302 0.137
R23958 VGND VGND.n2320 0.137
R23959 VGND.n2343 VGND 0.137
R23960 VGND.n2553 VGND 0.137
R23961 VGND.n2536 VGND 0.137
R23962 VGND.n2534 VGND 0.137
R23963 VGND.n2505 VGND 0.137
R23964 VGND.n2503 VGND 0.137
R23965 VGND VGND.n2890 0.137
R23966 VGND VGND.n2907 0.137
R23967 VGND VGND.n2919 0.137
R23968 VGND.n2942 VGND 0.137
R23969 VGND.n2932 VGND 0.137
R23970 VGND VGND.n1016 0.137
R23971 VGND.n2162 VGND 0.137
R23972 VGND.n2142 VGND 0.137
R23973 VGND.n2125 VGND 0.137
R23974 VGND.n2123 VGND 0.137
R23975 VGND.n2993 VGND 0.137
R23976 VGND.n2979 VGND 0.137
R23977 VGND VGND.n3046 0.137
R23978 VGND VGND.n3056 0.137
R23979 VGND VGND.n3061 0.137
R23980 VGND.n3099 VGND 0.137
R23981 VGND.n3092 VGND 0.137
R23982 VGND.n3086 VGND 0.137
R23983 VGND VGND.n3149 0.137
R23984 VGND VGND.n3161 0.137
R23985 VGND VGND.n3165 0.137
R23986 VGND.n3205 VGND 0.137
R23987 VGND.n3197 VGND 0.137
R23988 VGND.n3193 VGND 0.137
R23989 VGND VGND.n3276 0.137
R23990 VGND VGND.n3290 0.137
R23991 VGND VGND.n3293 0.137
R23992 VGND.n3334 VGND 0.137
R23993 VGND.n3325 VGND 0.137
R23994 VGND.n3738 VGND 0.137
R23995 VGND.n3736 VGND 0.137
R23996 VGND VGND.n3004 0.137
R23997 VGND VGND.n3013 0.137
R23998 VGND.n3037 VGND 0.137
R23999 VGND.n3028 VGND 0.137
R24000 VGND VGND.n3108 0.137
R24001 VGND VGND.n3117 0.137
R24002 VGND.n3142 VGND 0.137
R24003 VGND.n3133 VGND 0.137
R24004 VGND VGND.n3213 0.137
R24005 VGND VGND.n3222 0.137
R24006 VGND.n3271 VGND 0.137
R24007 VGND.n3262 VGND 0.137
R24008 VGND.n3252 VGND 0.137
R24009 VGND.n3243 VGND 0.137
R24010 VGND VGND.n3766 0.137
R24011 VGND.n819 VGND.n818 0.1355
R24012 VGND.n3463 VGND.n54 0.1355
R24013 VGND.n904 VGND.n903 0.1355
R24014 VGND.n908 VGND.n907 0.1355
R24015 VGND.n3687 VGND.n3686 0.1355
R24016 VGND.n1270 VGND.n1269 0.1355
R24017 VGND.n1528 VGND 0.1355
R24018 VGND.n2232 VGND.n2231 0.1355
R24019 VGND.n3719 VGND.n3718 0.1355
R24020 VGND.n3767 VGND.n0 0.1355
R24021 VGND.n864 VGND.n863 0.13475
R24022 VGND.n744 VGND.n743 0.134
R24023 VGND VGND.n1819 0.13325
R24024 VGND VGND.n1978 0.13325
R24025 VGND VGND.n886 0.1325
R24026 VGND VGND.n1577 0.1325
R24027 VGND.n1476 VGND.n1475 0.1325
R24028 VGND VGND.n1542 0.1325
R24029 VGND VGND.n1525 0.1325
R24030 VGND VGND.n3391 0.1325
R24031 VGND VGND.n1215 0.1325
R24032 VGND VGND.n1780 0.1325
R24033 VGND.n1766 VGND.n1765 0.1325
R24034 VGND VGND.n1753 0.1325
R24035 VGND.n1739 VGND.n1738 0.1325
R24036 VGND.n1798 VGND.n1797 0.1325
R24037 VGND VGND.n1102 0.1325
R24038 VGND.n1986 VGND.n1985 0.1325
R24039 VGND.n627 VGND 0.1325
R24040 VGND.n1934 VGND.n1933 0.1325
R24041 VGND VGND.n2409 0.1325
R24042 VGND.n2185 VGND 0.1325
R24043 VGND VGND.n2198 0.1325
R24044 VGND.n2045 VGND 0.1325
R24045 VGND.n862 VGND.n861 0.13175
R24046 VGND.n1932 VGND 0.13175
R24047 VGND.n1211 VGND.n1210 0.13025
R24048 VGND.n1956 VGND 0.1295
R24049 VGND VGND.n1955 0.1295
R24050 VGND.n2410 VGND.n470 0.1295
R24051 VGND.n2190 VGND 0.1295
R24052 VGND.n1437 VGND 0.12875
R24053 VGND.n3445 VGND 0.12875
R24054 VGND VGND.n1336 0.12875
R24055 VGND.n1574 VGND 0.12875
R24056 VGND.n1377 VGND 0.12875
R24057 VGND.n3418 VGND 0.12875
R24058 VGND VGND.n303 0.12875
R24059 VGND VGND.n306 0.12875
R24060 VGND.n1539 VGND 0.12875
R24061 VGND.n1130 VGND 0.12875
R24062 VGND.n1961 VGND 0.12875
R24063 VGND.n1948 VGND 0.12875
R24064 VGND VGND.n1799 0.12875
R24065 VGND.n1980 VGND 0.12875
R24066 VGND.n998 VGND 0.12875
R24067 VGND VGND.n2181 0.12875
R24068 VGND VGND.n2044 0.12875
R24069 VGND.n2091 VGND 0.12875
R24070 VGND.n163 VGND 0.12725
R24071 VGND VGND.n1965 0.12725
R24072 VGND.n1804 VGND 0.12725
R24073 VGND.n2063 VGND.n2062 0.12725
R24074 VGND.n3416 VGND.n3415 0.1265
R24075 VGND.n259 VGND.n258 0.1265
R24076 VGND.n1769 VGND 0.1265
R24077 VGND.n1755 VGND.n1754 0.1265
R24078 VGND VGND.n1909 0.1265
R24079 VGND VGND.n514 0.1265
R24080 VGND VGND.n2069 0.1265
R24081 VGND.n2087 VGND 0.1265
R24082 VGND VGND.n851 0.12575
R24083 VGND.n1553 VGND 0.12575
R24084 VGND VGND.n2038 0.12575
R24085 VGND VGND.n317 0.125
R24086 VGND.n1742 VGND 0.125
R24087 VGND.n1307 VGND 0.1235
R24088 VGND VGND.n1391 0.1235
R24089 VGND VGND.n1454 0.1235
R24090 VGND.n1513 VGND 0.1235
R24091 VGND.n3397 VGND.n3396 0.1235
R24092 VGND.n1442 VGND.n1441 0.122
R24093 VGND.n3148 VGND.n3147 0.122
R24094 VGND.n3144 VGND.n3143 0.122
R24095 VGND VGND.n1436 0.12125
R24096 VGND VGND.n1313 0.12125
R24097 VGND VGND.n1947 0.12125
R24098 VGND.n2180 VGND 0.12125
R24099 VGND VGND.n1316 0.1205
R24100 VGND.n1374 VGND 0.1205
R24101 VGND VGND.n346 0.1205
R24102 VGND.n1628 VGND 0.1205
R24103 VGND.n1525 VGND.n1524 0.1205
R24104 VGND.n1782 VGND.n1781 0.1205
R24105 VGND.n957 VGND 0.1205
R24106 VGND.n1057 VGND 0.1205
R24107 VGND VGND.n3757 0.1205
R24108 VGND.n172 VGND.n171 0.11975
R24109 VGND.n836 VGND 0.119
R24110 VGND.n1300 VGND.n1299 0.119
R24111 VGND.n1629 VGND 0.119
R24112 VGND VGND.n757 0.119
R24113 VGND VGND.n1766 0.11825
R24114 VGND VGND.n2388 0.11825
R24115 VGND.n1416 VGND.n1415 0.1175
R24116 VGND.n3444 VGND.n3443 0.1175
R24117 VGND.n1146 VGND.n1145 0.1175
R24118 VGND.n970 VGND.n969 0.1175
R24119 VGND.n935 VGND.n917 0.116
R24120 VGND.n3407 VGND.n198 0.116
R24121 VGND.n1042 VGND 0.116
R24122 VGND.n3272 VGND.n364 0.116
R24123 VGND.n930 VGND 0.1145
R24124 VGND VGND.n927 0.1145
R24125 VGND.n827 VGND 0.1145
R24126 VGND.n1418 VGND 0.1145
R24127 VGND.n164 VGND 0.1145
R24128 VGND.n170 VGND 0.1145
R24129 VGND.n177 VGND 0.1145
R24130 VGND VGND.n193 0.1145
R24131 VGND.n188 VGND 0.1145
R24132 VGND VGND.n239 0.1145
R24133 VGND VGND.n235 0.1145
R24134 VGND VGND.n232 0.1145
R24135 VGND.n62 VGND 0.1145
R24136 VGND VGND.n65 0.1145
R24137 VGND.n69 VGND 0.1145
R24138 VGND VGND.n78 0.1145
R24139 VGND.n83 VGND 0.1145
R24140 VGND.n85 VGND 0.1145
R24141 VGND.n93 VGND 0.1145
R24142 VGND VGND.n98 0.1145
R24143 VGND VGND.n901 0.1145
R24144 VGND VGND.n905 0.1145
R24145 VGND.n906 VGND 0.1145
R24146 VGND.n1310 VGND 0.1145
R24147 VGND.n1326 VGND 0.1145
R24148 VGND.n1329 VGND 0.1145
R24149 VGND VGND.n1340 0.1145
R24150 VGND VGND.n1589 0.1145
R24151 VGND.n328 VGND 0.1145
R24152 VGND VGND.n3690 0.1145
R24153 VGND VGND.n3687 0.1145
R24154 VGND VGND.n1275 0.1145
R24155 VGND VGND.n1271 0.1145
R24156 VGND.n1265 VGND 0.1145
R24157 VGND VGND.n1261 0.1145
R24158 VGND.n1255 VGND.n1254 0.1145
R24159 VGND VGND.n1252 0.1145
R24160 VGND VGND.n1247 0.1145
R24161 VGND VGND.n1627 0.1145
R24162 VGND.n1624 VGND 0.1145
R24163 VGND VGND.n1623 0.1145
R24164 VGND VGND.n1618 0.1145
R24165 VGND VGND.n1610 0.1145
R24166 VGND.n1607 VGND.n1606 0.1145
R24167 VGND VGND.n1604 0.1145
R24168 VGND VGND.n1465 0.1145
R24169 VGND VGND.n1557 0.1145
R24170 VGND VGND.n1547 0.1145
R24171 VGND VGND.n1535 0.1145
R24172 VGND VGND.n1520 0.1145
R24173 VGND.n1518 VGND 0.1145
R24174 VGND VGND.n3398 0.1145
R24175 VGND VGND.n3381 0.1145
R24176 VGND VGND.n1199 0.1145
R24177 VGND VGND.n1221 0.1145
R24178 VGND.n1217 VGND.n1216 0.1145
R24179 VGND.n1683 VGND 0.1145
R24180 VGND.n1696 VGND 0.1145
R24181 VGND VGND.n1715 0.1145
R24182 VGND VGND.n1714 0.1145
R24183 VGND VGND.n1740 0.1145
R24184 VGND.n3369 VGND.n3368 0.1145
R24185 VGND VGND.n1174 0.1145
R24186 VGND.n1156 VGND 0.1145
R24187 VGND VGND.n1155 0.1145
R24188 VGND VGND.n1152 0.1145
R24189 VGND.n1143 VGND.n1142 0.1145
R24190 VGND VGND.n1137 0.1145
R24191 VGND.n1132 VGND 0.1145
R24192 VGND VGND.n1131 0.1145
R24193 VGND.n746 VGND 0.1145
R24194 VGND.n1822 VGND.n1821 0.1145
R24195 VGND VGND.n1820 0.1145
R24196 VGND VGND.n721 0.1145
R24197 VGND.n1870 VGND.n1869 0.1145
R24198 VGND VGND.n1868 0.1145
R24199 VGND.n1852 VGND.n1851 0.1145
R24200 VGND VGND.n1850 0.1145
R24201 VGND.n1833 VGND.n1832 0.1145
R24202 VGND.n1102 VGND 0.1145
R24203 VGND VGND.n1091 0.1145
R24204 VGND.n1083 VGND 0.1145
R24205 VGND VGND.n1082 0.1145
R24206 VGND VGND.n576 0.1145
R24207 VGND VGND.n1991 0.1145
R24208 VGND.n637 VGND 0.1145
R24209 VGND VGND.n1918 0.1145
R24210 VGND VGND.n1916 0.1145
R24211 VGND VGND.n1915 0.1145
R24212 VGND VGND.n1904 0.1145
R24213 VGND.n1889 VGND.n1888 0.1145
R24214 VGND VGND.n1887 0.1145
R24215 VGND.n713 VGND.n712 0.1145
R24216 VGND VGND.n711 0.1145
R24217 VGND.n695 VGND.n694 0.1145
R24218 VGND VGND.n693 0.1145
R24219 VGND.n676 VGND.n675 0.1145
R24220 VGND.n1008 VGND.n1007 0.1145
R24221 VGND VGND.n955 0.1145
R24222 VGND.n2183 VGND 0.1145
R24223 VGND VGND.n2185 0.1145
R24224 VGND VGND.n2216 0.1145
R24225 VGND.n2589 VGND.n2588 0.1145
R24226 VGND VGND.n2587 0.1145
R24227 VGND.n2571 VGND.n2570 0.1145
R24228 VGND VGND.n2569 0.1145
R24229 VGND.n2839 VGND.n2838 0.1145
R24230 VGND.n2840 VGND 0.1145
R24231 VGND.n2862 VGND.n2861 0.1145
R24232 VGND VGND.n2860 0.1145
R24233 VGND.n2872 VGND.n2871 0.1145
R24234 VGND.n2612 VGND 0.1145
R24235 VGND.n2601 VGND 0.1145
R24236 VGND.n390 VGND 0.1145
R24237 VGND VGND.n387 0.1145
R24238 VGND.n2743 VGND.n2742 0.1145
R24239 VGND.n2744 VGND 0.1145
R24240 VGND.n2766 VGND.n2765 0.1145
R24241 VGND VGND.n2764 0.1145
R24242 VGND.n2813 VGND.n2812 0.1145
R24243 VGND VGND.n2811 0.1145
R24244 VGND.n2795 VGND.n2794 0.1145
R24245 VGND VGND.n2793 0.1145
R24246 VGND.n2776 VGND.n2775 0.1145
R24247 VGND.n2698 VGND.n2697 0.1145
R24248 VGND.n2681 VGND.n2680 0.1145
R24249 VGND VGND.n2679 0.1145
R24250 VGND.n441 VGND.n440 0.1145
R24251 VGND.n442 VGND 0.1145
R24252 VGND VGND.n2443 0.1145
R24253 VGND VGND.n2440 0.1145
R24254 VGND.n2431 VGND 0.1145
R24255 VGND.n2427 VGND.n2426 0.1145
R24256 VGND VGND.n2425 0.1145
R24257 VGND.n492 VGND.n491 0.1145
R24258 VGND.n494 VGND 0.1145
R24259 VGND VGND.n2366 0.1145
R24260 VGND VGND.n2361 0.1145
R24261 VGND.n541 VGND.n540 0.1145
R24262 VGND.n2482 VGND.n2481 0.1145
R24263 VGND.n2464 VGND.n2463 0.1145
R24264 VGND.n2230 VGND 0.1145
R24265 VGND VGND.n2233 0.1145
R24266 VGND.n2234 VGND 0.1145
R24267 VGND VGND.n2237 0.1145
R24268 VGND.n2243 VGND 0.1145
R24269 VGND.n2248 VGND.n2247 0.1145
R24270 VGND.n2249 VGND 0.1145
R24271 VGND.n2267 VGND.n2266 0.1145
R24272 VGND.n2268 VGND 0.1145
R24273 VGND.n2285 VGND.n2284 0.1145
R24274 VGND.n2286 VGND 0.1145
R24275 VGND.n2304 VGND.n2303 0.1145
R24276 VGND.n2305 VGND 0.1145
R24277 VGND.n2331 VGND.n2330 0.1145
R24278 VGND VGND.n2329 0.1145
R24279 VGND.n2342 VGND.n2341 0.1145
R24280 VGND VGND.n2491 0.1145
R24281 VGND VGND.n2531 0.1145
R24282 VGND.n2520 VGND 0.1145
R24283 VGND.n2517 VGND 0.1145
R24284 VGND VGND.n2500 0.1145
R24285 VGND VGND.n1020 0.1145
R24286 VGND VGND.n1018 0.1145
R24287 VGND.n1061 VGND 0.1145
R24288 VGND VGND.n1060 0.1145
R24289 VGND.n1050 VGND.n1049 0.1145
R24290 VGND VGND.n1047 0.1145
R24291 VGND.n1044 VGND 0.1145
R24292 VGND VGND.n1040 0.1145
R24293 VGND VGND.n1032 0.1145
R24294 VGND.n1024 VGND 0.1145
R24295 VGND.n2006 VGND 0.1145
R24296 VGND.n2009 VGND 0.1145
R24297 VGND.n2023 VGND 0.1145
R24298 VGND.n2027 VGND 0.1145
R24299 VGND.n2028 VGND 0.1145
R24300 VGND.n2161 VGND.n2160 0.1145
R24301 VGND VGND.n2159 0.1145
R24302 VGND.n2141 VGND.n2140 0.1145
R24303 VGND.n2124 VGND.n2123 0.1145
R24304 VGND VGND.n2122 0.1145
R24305 VGND VGND.n2967 0.1145
R24306 VGND VGND.n2966 0.1145
R24307 VGND VGND.n2996 0.1145
R24308 VGND VGND.n2984 0.1145
R24309 VGND.n3059 VGND 0.1145
R24310 VGND VGND.n3089 0.1145
R24311 VGND.n3164 VGND 0.1145
R24312 VGND VGND.n3194 0.1145
R24313 VGND.n3293 VGND 0.1145
R24314 VGND VGND.n3734 0.1145
R24315 VGND VGND.n84 0.11375
R24316 VGND VGND.n90 0.11375
R24317 VGND.n104 VGND 0.11375
R24318 VGND VGND.n1579 0.11375
R24319 VGND.n503 VGND 0.11375
R24320 VGND VGND.n2543 0.11375
R24321 VGND.n2900 VGND 0.11375
R24322 VGND.n2033 VGND 0.11375
R24323 VGND.n3056 VGND 0.11375
R24324 VGND VGND.n3064 0.11375
R24325 VGND.n3159 VGND 0.11375
R24326 VGND VGND.n3170 0.11375
R24327 VGND.n3286 VGND 0.11375
R24328 VGND VGND.n3300 0.11375
R24329 VGND VGND.n3744 0.11375
R24330 VGND VGND.n3726 0.11375
R24331 VGND.n183 VGND 0.113
R24332 VGND.n1284 VGND.n1283 0.113
R24333 VGND.n1286 VGND.n1285 0.113
R24334 VGND.n1288 VGND.n1287 0.113
R24335 VGND VGND.n1337 0.113
R24336 VGND.n1575 VGND 0.113
R24337 VGND.n1105 VGND 0.113
R24338 VGND.n1101 VGND.n1100 0.113
R24339 VGND.n1094 VGND.n1093 0.113
R24340 VGND.n2430 VGND.n2429 0.113
R24341 VGND VGND.n2550 0.113
R24342 VGND.n2516 VGND.n2515 0.113
R24343 VGND.n2895 VGND 0.113
R24344 VGND VGND.n375 0.113
R24345 VGND VGND.n817 0.11225
R24346 VGND VGND.n1678 0.11225
R24347 VGND VGND.n634 0.11225
R24348 VGND VGND.n3433 0.1115
R24349 VGND.n218 VGND.n217 0.1115
R24350 VGND.n3426 VGND.n3425 0.1115
R24351 VGND.n1950 VGND.n1949 0.1115
R24352 VGND.n516 VGND.n515 0.1115
R24353 VGND.n2167 VGND.n2166 0.1115
R24354 VGND.n1469 VGND 0.11075
R24355 VGND.n1978 VGND.n1977 0.11075
R24356 VGND.n1230 VGND 0.11
R24357 VGND VGND.n1189 0.11
R24358 VGND VGND.n1187 0.11
R24359 VGND VGND.n1075 0.11
R24360 VGND.n1107 VGND 0.11
R24361 VGND.n1992 VGND 0.11
R24362 VGND VGND.n994 0.11
R24363 VGND VGND.n992 0.11
R24364 VGND.n987 VGND 0.11
R24365 VGND VGND.n986 0.11
R24366 VGND.n985 VGND 0.11
R24367 VGND.n964 VGND 0.11
R24368 VGND VGND.n463 0.11
R24369 VGND VGND.n2461 0.11
R24370 VGND.n2225 VGND 0.11
R24371 VGND VGND.n2241 0.11
R24372 VGND VGND.n1056 0.11
R24373 VGND.n1055 VGND 0.11
R24374 VGND VGND.n1052 0.11
R24375 VGND.n1051 VGND 0.11
R24376 VGND.n3208 VGND 0.11
R24377 VGND.n171 VGND.n170 0.10925
R24378 VGND.n226 VGND.n225 0.10925
R24379 VGND.n84 VGND.n83 0.10925
R24380 VGND.n90 VGND.n89 0.10925
R24381 VGND.n94 VGND.n93 0.10925
R24382 VGND.n105 VGND.n104 0.10925
R24383 VGND.n1309 VGND.n1308 0.10925
R24384 VGND.n1601 VGND.n1600 0.10925
R24385 VGND.n2053 VGND.n2052 0.10925
R24386 VGND VGND.n3672 0.1085
R24387 VGND.n3483 VGND 0.1085
R24388 VGND.n3635 VGND 0.1085
R24389 VGND.n3650 VGND 0.1085
R24390 VGND.n3466 VGND 0.1085
R24391 VGND VGND.n3574 0.1085
R24392 VGND VGND.n3606 0.1085
R24393 VGND VGND.n3622 0.1085
R24394 VGND VGND.n3590 0.1085
R24395 VGND VGND.n3558 0.1085
R24396 VGND.n3540 VGND 0.1085
R24397 VGND VGND.n3703 0.1085
R24398 VGND.n22 VGND 0.1085
R24399 VGND.n3495 VGND 0.1085
R24400 VGND.n3510 VGND 0.1085
R24401 VGND.n3525 VGND 0.1085
R24402 VGND.n809 VGND.n808 0.1085
R24403 VGND.n828 VGND.n827 0.1085
R24404 VGND.n1417 VGND 0.1085
R24405 VGND.n3441 VGND.n3440 0.1085
R24406 VGND.n134 VGND.n133 0.1085
R24407 VGND.n132 VGND.n131 0.1085
R24408 VGND.n130 VGND.n129 0.1085
R24409 VGND.n125 VGND.n124 0.1085
R24410 VGND VGND.n169 0.1085
R24411 VGND.n184 VGND.n183 0.1085
R24412 VGND.n232 VGND.n231 0.1085
R24413 VGND.n71 VGND.n70 0.1085
R24414 VGND.n1311 VGND.n1310 0.1085
R24415 VGND.n1321 VGND.n1320 0.1085
R24416 VGND.n1331 VGND.n1330 0.1085
R24417 VGND.n1333 VGND.n1332 0.1085
R24418 VGND.n1335 VGND.n1334 0.1085
R24419 VGND.n1594 VGND.n1593 0.1085
R24420 VGND VGND.n1567 0.1085
R24421 VGND.n310 VGND.n309 0.1085
R24422 VGND.n1243 VGND.n1242 0.1085
R24423 VGND VGND.n1262 0.1085
R24424 VGND.n1627 VGND.n1626 0.1085
R24425 VGND.n1614 VGND.n1613 0.1085
R24426 VGND.n1604 VGND.n1603 0.1085
R24427 VGND.n1478 VGND 0.1085
R24428 VGND.n1559 VGND.n1558 0.1085
R24429 VGND.n1537 VGND.n1536 0.1085
R24430 VGND.n253 VGND 0.1085
R24431 VGND.n255 VGND.n254 0.1085
R24432 VGND.n1233 VGND.n1232 0.1085
R24433 VGND.n1227 VGND.n1226 0.1085
R24434 VGND.n1638 VGND.n1637 0.1085
R24435 VGND.n1702 VGND.n1701 0.1085
R24436 VGND.n1707 VGND.n1706 0.1085
R24437 VGND.n1775 VGND.n1774 0.1085
R24438 VGND VGND.n1746 0.1085
R24439 VGND.n1736 VGND.n1735 0.1085
R24440 VGND.n1120 VGND.n1119 0.1085
R24441 VGND.n1118 VGND.n1117 0.1085
R24442 VGND.n1149 VGND.n1148 0.1085
R24443 VGND.n1072 VGND.n1071 0.1085
R24444 VGND.n1070 VGND.n1069 0.1085
R24445 VGND.n1096 VGND.n1095 0.1085
R24446 VGND VGND.n1085 0.1085
R24447 VGND.n1999 VGND.n1998 0.1085
R24448 VGND.n1995 VGND.n1994 0.1085
R24449 VGND.n641 VGND.n640 0.1085
R24450 VGND VGND.n1928 0.1085
R24451 VGND.n1926 VGND.n1925 0.1085
R24452 VGND VGND.n1920 0.1085
R24453 VGND.n1911 VGND.n1910 0.1085
R24454 VGND.n1903 VGND.n1902 0.1085
R24455 VGND VGND.n984 0.1085
R24456 VGND.n984 VGND.n983 0.1085
R24457 VGND.n973 VGND.n972 0.1085
R24458 VGND.n967 VGND.n966 0.1085
R24459 VGND.n2408 VGND 0.1085
R24460 VGND.n2397 VGND.n2396 0.1085
R24461 VGND.n2392 VGND.n2391 0.1085
R24462 VGND VGND.n2217 0.1085
R24463 VGND VGND.n2564 0.1085
R24464 VGND.n413 VGND 0.1085
R24465 VGND.n2624 VGND 0.1085
R24466 VGND.n460 VGND.n459 0.1085
R24467 VGND.n458 VGND.n457 0.1085
R24468 VGND.n2436 VGND.n2435 0.1085
R24469 VGND.n2432 VGND.n2431 0.1085
R24470 VGND.n512 VGND.n511 0.1085
R24471 VGND.n2366 VGND.n2365 0.1085
R24472 VGND.n2360 VGND.n2359 0.1085
R24473 VGND.n2458 VGND.n2457 0.1085
R24474 VGND.n2456 VGND.n2455 0.1085
R24475 VGND.n1016 VGND 0.1085
R24476 VGND.n1059 VGND 0.1085
R24477 VGND.n2014 VGND.n2013 0.1085
R24478 VGND.n2018 VGND.n2017 0.1085
R24479 VGND.n2031 VGND.n2030 0.1085
R24480 VGND.n196 VGND 0.107
R24481 VGND.n982 VGND.n981 0.107
R24482 VGND.n2446 VGND.n2445 0.107
R24483 VGND.n2524 VGND.n2523 0.107
R24484 VGND.n2078 VGND.n2077 0.107
R24485 VGND.n1385 VGND.n1384 0.1055
R24486 VGND.n1531 VGND.n1530 0.1055
R24487 VGND VGND.n1690 0.1055
R24488 VGND.n1957 VGND.n1956 0.1055
R24489 VGND.n1794 VGND.n767 0.1055
R24490 VGND VGND.n1048 0.104
R24491 VGND VGND.n1034 0.104
R24492 VGND.n294 VGND.n293 0.1025
R24493 VGND VGND.n256 0.1025
R24494 VGND.n1781 VGND 0.1025
R24495 VGND.n2372 VGND.n2371 0.1025
R24496 VGND.n2165 VGND 0.1025
R24497 VGND.n3339 VGND.n3338 0.1025
R24498 VGND.n3335 VGND.n3334 0.1025
R24499 VGND.n3253 VGND.n3252 0.1025
R24500 VGND VGND.n911 0.101
R24501 VGND.n241 VGND 0.101
R24502 VGND.n1643 VGND 0.101
R24503 VGND.n1943 VGND.n1942 0.101
R24504 VGND.n1906 VGND 0.101
R24505 VGND.n2363 VGND 0.101
R24506 VGND.n1579 VGND 0.0995
R24507 VGND VGND.n1691 0.0995
R24508 VGND.n1874 VGND.n1873 0.0995
R24509 VGND.n817 VGND 0.09875
R24510 VGND.n820 VGND 0.09875
R24511 VGND VGND.n64 0.09875
R24512 VGND VGND.n85 0.09875
R24513 VGND.n1379 VGND 0.09875
R24514 VGND VGND.n328 0.09875
R24515 VGND.n1247 VGND 0.09875
R24516 VGND.n1534 VGND 0.09875
R24517 VGND.n1504 VGND 0.09875
R24518 VGND VGND.n1647 0.09875
R24519 VGND VGND.n1669 0.09875
R24520 VGND.n3376 VGND 0.09875
R24521 VGND.n1159 VGND 0.09875
R24522 VGND VGND.n746 0.09875
R24523 VGND.n748 VGND.n747 0.09875
R24524 VGND VGND.n1103 0.09875
R24525 VGND.n1086 VGND 0.09875
R24526 VGND VGND.n638 0.09875
R24527 VGND.n1929 VGND 0.09875
R24528 VGND.n1900 VGND 0.09875
R24529 VGND VGND.n2188 0.09875
R24530 VGND.n519 VGND 0.09875
R24531 VGND.n2357 VGND 0.09875
R24532 VGND VGND.n2228 0.09875
R24533 VGND VGND.n2061 0.09875
R24534 VGND.n1587 VGND 0.09725
R24535 VGND.n2178 VGND.n2177 0.09725
R24536 VGND.n859 VGND 0.0965
R24537 VGND.n885 VGND.n867 0.0965
R24538 VGND VGND.n1404 0.0965
R24539 VGND.n1411 VGND.n1410 0.0965
R24540 VGND.n165 VGND.n164 0.0965
R24541 VGND.n243 VGND 0.0965
R24542 VGND.n242 VGND.n241 0.0965
R24543 VGND.n1316 VGND 0.0965
R24544 VGND VGND.n1588 0.0965
R24545 VGND.n320 VGND.n319 0.0965
R24546 VGND VGND.n1628 0.0965
R24547 VGND VGND.n1622 0.0965
R24548 VGND.n1602 VGND 0.0965
R24549 VGND.n3401 VGND.n3400 0.0965
R24550 VGND VGND.n3380 0.0965
R24551 VGND.n1212 VGND 0.0965
R24552 VGND VGND.n1209 0.0965
R24553 VGND VGND.n1758 0.0965
R24554 VGND.n1752 VGND.n1751 0.0965
R24555 VGND VGND.n749 0.0965
R24556 VGND.n1991 VGND 0.0965
R24557 VGND VGND.n637 0.0965
R24558 VGND.n1907 VGND.n1906 0.0965
R24559 VGND.n2656 VGND.n2655 0.0965
R24560 VGND.n511 VGND.n510 0.0965
R24561 VGND.n2364 VGND.n2363 0.0965
R24562 VGND VGND.n2032 0.0965
R24563 VGND VGND.n2081 0.0965
R24564 VGND.n3103 VGND.n375 0.0965
R24565 VGND.n3106 VGND.n373 0.0965
R24566 VGND.t2010 VGND.t5880 0.0958694
R24567 VGND.t34 VGND.n55 0.0958694
R24568 VGND.t5706 VGND.t2 0.0958694
R24569 VGND.t3072 VGND.t1059 0.0958694
R24570 VGND.t6697 VGND.t3682 0.0958694
R24571 VGND.n3338 VGND 0.09575
R24572 VGND VGND.n1394 0.095
R24573 VGND.n1692 VGND 0.095
R24574 VGND.n2062 VGND 0.095
R24575 VGND.n867 VGND.n866 0.09425
R24576 VGND VGND.n3442 0.09425
R24577 VGND.n65 VGND 0.09425
R24578 VGND.n1319 VGND 0.09425
R24579 VGND VGND.n1578 0.09425
R24580 VGND.n302 VGND 0.09425
R24581 VGND.n316 VGND.n315 0.09425
R24582 VGND VGND.n3386 0.09425
R24583 VGND VGND.n1235 0.09425
R24584 VGND.n639 VGND 0.09425
R24585 VGND VGND.n2517 0.09425
R24586 VGND.n917 VGND.n916 0.09275
R24587 VGND.n3429 VGND 0.09275
R24588 VGND.n823 VGND.n822 0.09125
R24589 VGND.n636 VGND.n635 0.09125
R24590 VGND.n1922 VGND.n1921 0.09125
R24591 VGND.n220 VGND.n219 0.0905
R24592 VGND.n222 VGND.n221 0.0905
R24593 VGND.n325 VGND 0.0905
R24594 VGND.n1273 VGND 0.0905
R24595 VGND VGND.n1621 0.0905
R24596 VGND.n3388 VGND.n3387 0.0905
R24597 VGND VGND.n1682 0.0905
R24598 VGND VGND.n1750 0.0905
R24599 VGND.n956 VGND 0.0905
R24600 VGND.n2369 VGND.n2368 0.0905
R24601 VGND VGND.n2163 0.0905
R24602 VGND.n1189 VGND.n1188 0.089
R24603 VGND.n1187 VGND.n1186 0.089
R24604 VGND.n1179 VGND.n1178 0.089
R24605 VGND.n1168 VGND.n1167 0.089
R24606 VGND.n1141 VGND.n1140 0.089
R24607 VGND.n996 VGND.n995 0.089
R24608 VGND.n994 VGND.n993 0.089
R24609 VGND.n992 VGND.n991 0.089
R24610 VGND.n988 VGND.n987 0.089
R24611 VGND.n2529 VGND.n2528 0.089
R24612 VGND VGND.n931 0.0875
R24613 VGND.n929 VGND.n928 0.0875
R24614 VGND VGND.n924 0.0875
R24615 VGND.n195 VGND.n194 0.0875
R24616 VGND.n3431 VGND.n3430 0.0875
R24617 VGND VGND.n321 0.0875
R24618 VGND.n1463 VGND.n1462 0.0875
R24619 VGND VGND.n3402 0.0875
R24620 VGND.n1238 VGND.n1192 0.0875
R24621 VGND.n1667 VGND 0.0875
R24622 VGND.n1699 VGND.n1698 0.0875
R24623 VGND.n1771 VGND.n1770 0.0875
R24624 VGND VGND.n1974 0.0875
R24625 VGND.n950 VGND.n470 0.0875
R24626 VGND.n2368 VGND 0.0875
R24627 VGND.n2038 VGND 0.0875
R24628 VGND VGND.n176 0.08675
R24629 VGND.n1438 VGND 0.086
R24630 VGND.n1949 VGND 0.086
R24631 VGND VGND.n2449 0.086
R24632 VGND.n751 VGND.n750 0.08525
R24633 VGND.n2034 VGND.n2033 0.08525
R24634 VGND.n927 VGND.n926 0.0845
R24635 VGND VGND.n816 0.0845
R24636 VGND.n857 VGND.n856 0.0845
R24637 VGND.n1419 VGND.n1418 0.0845
R24638 VGND.n216 VGND.n215 0.0845
R24639 VGND VGND.n61 0.0845
R24640 VGND.n77 VGND.n76 0.0845
R24641 VGND.n87 VGND.n86 0.0845
R24642 VGND.n89 VGND.n88 0.0845
R24643 VGND.n110 VGND 0.0845
R24644 VGND.n108 VGND.n107 0.0845
R24645 VGND.n106 VGND.n105 0.0845
R24646 VGND.n901 VGND.n900 0.0845
R24647 VGND.n903 VGND.n902 0.0845
R24648 VGND.n1312 VGND.n1311 0.0845
R24649 VGND VGND.n1318 0.0845
R24650 VGND.n1346 VGND.n1345 0.0845
R24651 VGND.n309 VGND.n308 0.0845
R24652 VGND.n332 VGND.n331 0.0845
R24653 VGND.n337 VGND.n336 0.0845
R24654 VGND.n339 VGND.n338 0.0845
R24655 VGND.n1275 VGND.n1274 0.0845
R24656 VGND.n1268 VGND.n1267 0.0845
R24657 VGND.n1266 VGND.n1265 0.0845
R24658 VGND.n1264 VGND.n1263 0.0845
R24659 VGND.n1261 VGND.n1260 0.0845
R24660 VGND.n1257 VGND.n1256 0.0845
R24661 VGND.n1615 VGND.n1614 0.0845
R24662 VGND VGND.n1479 0.0845
R24663 VGND.n1515 VGND.n1514 0.0845
R24664 VGND.n3406 VGND.n3405 0.0845
R24665 VGND.n1201 VGND.n1200 0.0845
R24666 VGND.n1199 VGND.n1198 0.0845
R24667 VGND.n1193 VGND.n1192 0.0845
R24668 VGND.n1237 VGND.n1236 0.0845
R24669 VGND.n1221 VGND.n1220 0.0845
R24670 VGND.n1219 VGND.n1218 0.0845
R24671 VGND.n1681 VGND.n1680 0.0845
R24672 VGND.n1701 VGND.n1700 0.0845
R24673 VGND.n1785 VGND 0.0845
R24674 VGND.n1776 VGND.n1775 0.0845
R24675 VGND.n3375 VGND.n3374 0.0845
R24676 VGND.n3373 VGND.n3372 0.0845
R24677 VGND.n3371 VGND.n3370 0.0845
R24678 VGND.n1185 VGND.n1184 0.0845
R24679 VGND.n1177 VGND.n1176 0.0845
R24680 VGND.n1174 VGND.n1173 0.0845
R24681 VGND.n1166 VGND.n1165 0.0845
R24682 VGND.n1163 VGND 0.0845
R24683 VGND.n1139 VGND.n1138 0.0845
R24684 VGND.n1868 VGND.n1867 0.0845
R24685 VGND.n1866 VGND.n1865 0.0845
R24686 VGND.n1864 VGND.n1863 0.0845
R24687 VGND.n1862 VGND.n1861 0.0845
R24688 VGND.n1860 VGND.n1859 0.0845
R24689 VGND.n1858 VGND.n1857 0.0845
R24690 VGND.n1856 VGND.n1855 0.0845
R24691 VGND.n1854 VGND.n1853 0.0845
R24692 VGND.n1850 VGND.n1849 0.0845
R24693 VGND.n1848 VGND.n1847 0.0845
R24694 VGND.n1846 VGND.n1845 0.0845
R24695 VGND.n1844 VGND.n1843 0.0845
R24696 VGND.n1841 VGND.n1840 0.0845
R24697 VGND.n1839 VGND.n1838 0.0845
R24698 VGND.n1837 VGND.n1836 0.0845
R24699 VGND.n1835 VGND.n1834 0.0845
R24700 VGND.n1104 VGND 0.0845
R24701 VGND VGND.n629 0.0845
R24702 VGND.n1928 VGND.n1927 0.0845
R24703 VGND.n1920 VGND.n1919 0.0845
R24704 VGND.n1918 VGND.n1917 0.0845
R24705 VGND.n1899 VGND.n1898 0.0845
R24706 VGND.n1897 VGND.n1896 0.0845
R24707 VGND.n1895 VGND.n1894 0.0845
R24708 VGND.n1893 VGND.n1892 0.0845
R24709 VGND.n1891 VGND.n1890 0.0845
R24710 VGND.n1887 VGND.n1886 0.0845
R24711 VGND.n1885 VGND.n1884 0.0845
R24712 VGND.n1883 VGND.n1882 0.0845
R24713 VGND.n1881 VGND.n1880 0.0845
R24714 VGND.n719 VGND.n718 0.0845
R24715 VGND.n717 VGND.n716 0.0845
R24716 VGND.n715 VGND.n714 0.0845
R24717 VGND.n711 VGND.n710 0.0845
R24718 VGND.n709 VGND.n708 0.0845
R24719 VGND.n707 VGND.n706 0.0845
R24720 VGND.n705 VGND.n704 0.0845
R24721 VGND.n703 VGND.n702 0.0845
R24722 VGND.n701 VGND.n700 0.0845
R24723 VGND.n699 VGND.n698 0.0845
R24724 VGND.n697 VGND.n696 0.0845
R24725 VGND.n693 VGND.n692 0.0845
R24726 VGND.n691 VGND.n690 0.0845
R24727 VGND.n689 VGND.n688 0.0845
R24728 VGND.n687 VGND.n686 0.0845
R24729 VGND.n684 VGND.n683 0.0845
R24730 VGND.n682 VGND.n681 0.0845
R24731 VGND.n680 VGND.n679 0.0845
R24732 VGND.n678 VGND.n677 0.0845
R24733 VGND.n939 VGND.n938 0.0845
R24734 VGND.n937 VGND.n936 0.0845
R24735 VGND.n1010 VGND.n1009 0.0845
R24736 VGND.n960 VGND.n959 0.0845
R24737 VGND.n2563 VGND.n2562 0.0845
R24738 VGND.n2561 VGND.n2560 0.0845
R24739 VGND.n2597 VGND.n2596 0.0845
R24740 VGND.n2595 VGND.n2594 0.0845
R24741 VGND.n2593 VGND.n2592 0.0845
R24742 VGND.n2591 VGND.n2590 0.0845
R24743 VGND.n2587 VGND.n2586 0.0845
R24744 VGND.n2585 VGND.n2584 0.0845
R24745 VGND.n2583 VGND.n2582 0.0845
R24746 VGND.n2581 VGND.n2580 0.0845
R24747 VGND.n2579 VGND.n2578 0.0845
R24748 VGND.n2577 VGND.n2576 0.0845
R24749 VGND.n2575 VGND.n2574 0.0845
R24750 VGND.n2573 VGND.n2572 0.0845
R24751 VGND.n2569 VGND.n2568 0.0845
R24752 VGND.n2567 VGND.n2566 0.0845
R24753 VGND.n2565 VGND.n410 0.0845
R24754 VGND.n2829 VGND.n2828 0.0845
R24755 VGND.n2831 VGND.n2830 0.0845
R24756 VGND.n2833 VGND.n2832 0.0845
R24757 VGND.n2835 VGND.n2834 0.0845
R24758 VGND.n2837 VGND.n2836 0.0845
R24759 VGND.n2841 VGND.n2840 0.0845
R24760 VGND.n2843 VGND.n2842 0.0845
R24761 VGND.n2845 VGND.n2844 0.0845
R24762 VGND.n2847 VGND.n2846 0.0845
R24763 VGND.n2849 VGND.n2848 0.0845
R24764 VGND.n2851 VGND.n2850 0.0845
R24765 VGND.n2853 VGND.n2852 0.0845
R24766 VGND.n2855 VGND.n2854 0.0845
R24767 VGND.n2860 VGND.n2859 0.0845
R24768 VGND.n2858 VGND.n2857 0.0845
R24769 VGND.n2856 VGND.n409 0.0845
R24770 VGND.n2882 VGND.n2881 0.0845
R24771 VGND.n2880 VGND.n2879 0.0845
R24772 VGND.n2878 VGND.n2877 0.0845
R24773 VGND.n2876 VGND.n2875 0.0845
R24774 VGND.n2874 VGND.n2873 0.0845
R24775 VGND.n415 VGND.n414 0.0845
R24776 VGND.n417 VGND.n416 0.0845
R24777 VGND.n2735 VGND.n2734 0.0845
R24778 VGND.n2737 VGND.n2736 0.0845
R24779 VGND.n2739 VGND.n2738 0.0845
R24780 VGND.n2741 VGND.n2740 0.0845
R24781 VGND.n2745 VGND.n2744 0.0845
R24782 VGND.n2747 VGND.n2746 0.0845
R24783 VGND.n2749 VGND.n2748 0.0845
R24784 VGND.n2751 VGND.n2750 0.0845
R24785 VGND.n2753 VGND.n2752 0.0845
R24786 VGND.n2755 VGND.n2754 0.0845
R24787 VGND.n2757 VGND.n2756 0.0845
R24788 VGND.n2759 VGND.n2758 0.0845
R24789 VGND.n2764 VGND.n2763 0.0845
R24790 VGND.n2762 VGND.n2761 0.0845
R24791 VGND.n2760 VGND.n412 0.0845
R24792 VGND.n2823 VGND.n2822 0.0845
R24793 VGND.n2821 VGND.n2820 0.0845
R24794 VGND.n2819 VGND.n2818 0.0845
R24795 VGND.n2817 VGND.n2816 0.0845
R24796 VGND.n2815 VGND.n2814 0.0845
R24797 VGND.n2811 VGND.n2810 0.0845
R24798 VGND.n2809 VGND.n2808 0.0845
R24799 VGND.n2807 VGND.n2806 0.0845
R24800 VGND.n2805 VGND.n2804 0.0845
R24801 VGND.n2803 VGND.n2802 0.0845
R24802 VGND.n2801 VGND.n2800 0.0845
R24803 VGND.n2799 VGND.n2798 0.0845
R24804 VGND.n2797 VGND.n2796 0.0845
R24805 VGND.n2793 VGND.n2792 0.0845
R24806 VGND.n2791 VGND.n2790 0.0845
R24807 VGND.n2789 VGND.n2788 0.0845
R24808 VGND.n2786 VGND.n2785 0.0845
R24809 VGND.n2784 VGND.n2783 0.0845
R24810 VGND.n2782 VGND.n2781 0.0845
R24811 VGND.n2780 VGND.n2779 0.0845
R24812 VGND.n2778 VGND.n2777 0.0845
R24813 VGND.n2627 VGND.n2626 0.0845
R24814 VGND.n2625 VGND.n2623 0.0845
R24815 VGND.n2726 VGND.n2725 0.0845
R24816 VGND.n2724 VGND.n2723 0.0845
R24817 VGND.n2722 VGND.n2721 0.0845
R24818 VGND.n2720 VGND.n2719 0.0845
R24819 VGND.n2717 VGND.n2716 0.0845
R24820 VGND.n2714 VGND.n2713 0.0845
R24821 VGND.n2712 VGND.n2711 0.0845
R24822 VGND.n2710 VGND.n2709 0.0845
R24823 VGND.n2708 VGND.n2707 0.0845
R24824 VGND.n2706 VGND.n2705 0.0845
R24825 VGND.n2704 VGND.n2703 0.0845
R24826 VGND.n2702 VGND.n2701 0.0845
R24827 VGND.n2696 VGND.n2695 0.0845
R24828 VGND.n2694 VGND.n2693 0.0845
R24829 VGND.n2691 VGND.n2690 0.0845
R24830 VGND.n2687 VGND.n2686 0.0845
R24831 VGND.n2685 VGND.n2684 0.0845
R24832 VGND.n2683 VGND.n2682 0.0845
R24833 VGND.n2678 VGND.n2677 0.0845
R24834 VGND.n2676 VGND.n2675 0.0845
R24835 VGND.n2674 VGND.n2673 0.0845
R24836 VGND.n2670 VGND.n2669 0.0845
R24837 VGND.n2668 VGND.n2667 0.0845
R24838 VGND.n2666 VGND.n2665 0.0845
R24839 VGND.n2664 VGND.n2663 0.0845
R24840 VGND.n2661 VGND.n2660 0.0845
R24841 VGND.n2659 VGND.n2658 0.0845
R24842 VGND.n2657 VGND.n2656 0.0845
R24843 VGND.n2654 VGND.n2653 0.0845
R24844 VGND.n2652 VGND.n2651 0.0845
R24845 VGND.n2650 VGND.n2649 0.0845
R24846 VGND.n2648 VGND.n2647 0.0845
R24847 VGND.n2646 VGND.n2645 0.0845
R24848 VGND.n432 VGND.n431 0.0845
R24849 VGND.n434 VGND.n433 0.0845
R24850 VGND.n439 VGND.n438 0.0845
R24851 VGND.n2425 VGND.n2424 0.0845
R24852 VGND.n2423 VGND.n2422 0.0845
R24853 VGND.n2421 VGND.n2420 0.0845
R24854 VGND.n2419 VGND.n2418 0.0845
R24855 VGND.n2417 VGND.n2416 0.0845
R24856 VGND.n2415 VGND.n2414 0.0845
R24857 VGND.n488 VGND.n468 0.0845
R24858 VGND.n490 VGND.n489 0.0845
R24859 VGND.n518 VGND.n517 0.0845
R24860 VGND.n2356 VGND.n2355 0.0845
R24861 VGND.n2354 VGND.n2353 0.0845
R24862 VGND.n547 VGND.n546 0.0845
R24863 VGND.n545 VGND.n544 0.0845
R24864 VGND.n543 VGND.n542 0.0845
R24865 VGND.n423 VGND.n422 0.0845
R24866 VGND.n421 VGND.n420 0.0845
R24867 VGND.n2484 VGND.n2483 0.0845
R24868 VGND.n2478 VGND.n2477 0.0845
R24869 VGND.n2476 VGND.n2475 0.0845
R24870 VGND.n2474 VGND.n2473 0.0845
R24871 VGND.n2472 VGND.n2471 0.0845
R24872 VGND.n2468 VGND.n2467 0.0845
R24873 VGND.n2466 VGND.n2465 0.0845
R24874 VGND.n2237 VGND.n2236 0.0845
R24875 VGND.n2239 VGND.n2238 0.0845
R24876 VGND.n2244 VGND.n2243 0.0845
R24877 VGND.n2250 VGND.n2249 0.0845
R24878 VGND.n2252 VGND.n2251 0.0845
R24879 VGND.n2254 VGND.n2253 0.0845
R24880 VGND.n2256 VGND.n2255 0.0845
R24881 VGND.n2258 VGND.n2257 0.0845
R24882 VGND.n2260 VGND.n2259 0.0845
R24883 VGND.n2263 VGND.n2262 0.0845
R24884 VGND.n2265 VGND.n2264 0.0845
R24885 VGND.n2269 VGND.n2268 0.0845
R24886 VGND.n2271 VGND.n2270 0.0845
R24887 VGND.n2273 VGND.n2272 0.0845
R24888 VGND.n2275 VGND.n2274 0.0845
R24889 VGND.n2277 VGND.n2276 0.0845
R24890 VGND.n2279 VGND.n2278 0.0845
R24891 VGND.n2281 VGND.n2280 0.0845
R24892 VGND.n2283 VGND.n2282 0.0845
R24893 VGND.n2287 VGND.n2286 0.0845
R24894 VGND.n2289 VGND.n2288 0.0845
R24895 VGND.n2291 VGND.n2290 0.0845
R24896 VGND.n2293 VGND.n2292 0.0845
R24897 VGND.n2295 VGND.n2294 0.0845
R24898 VGND.n2300 VGND.n2299 0.0845
R24899 VGND.n2302 VGND.n2301 0.0845
R24900 VGND.n2306 VGND.n2305 0.0845
R24901 VGND.n2308 VGND.n2307 0.0845
R24902 VGND.n2310 VGND.n2309 0.0845
R24903 VGND.n2312 VGND.n2311 0.0845
R24904 VGND.n2314 VGND.n2313 0.0845
R24905 VGND.n2316 VGND.n2315 0.0845
R24906 VGND.n2318 VGND.n2317 0.0845
R24907 VGND.n2320 VGND.n2319 0.0845
R24908 VGND.n2329 VGND.n2328 0.0845
R24909 VGND.n2327 VGND.n2326 0.0845
R24910 VGND.n2325 VGND.n2324 0.0845
R24911 VGND.n2323 VGND.n2322 0.0845
R24912 VGND.n2321 VGND.n2222 0.0845
R24913 VGND.n2348 VGND.n2347 0.0845
R24914 VGND.n2346 VGND.n2345 0.0845
R24915 VGND.n2344 VGND.n2343 0.0845
R24916 VGND.n2527 VGND.n2526 0.0845
R24917 VGND.n2523 VGND.n2522 0.0845
R24918 VGND.n2521 VGND.n2520 0.0845
R24919 VGND.n2519 VGND.n2518 0.0845
R24920 VGND.n1064 VGND.n1063 0.0845
R24921 VGND.n1047 VGND.n1046 0.0845
R24922 VGND.n1045 VGND.n1044 0.0845
R24923 VGND.n1043 VGND.n1042 0.0845
R24924 VGND.n1034 VGND.n1033 0.0845
R24925 VGND.n1032 VGND.n1031 0.0845
R24926 VGND.n1025 VGND.n1024 0.0845
R24927 VGND.n2007 VGND.n2006 0.0845
R24928 VGND.n2010 VGND.n2009 0.0845
R24929 VGND VGND.n2012 0.0845
R24930 VGND.n2051 VGND 0.0845
R24931 VGND VGND.n2057 0.0845
R24932 VGND.n2075 VGND.n2074 0.0845
R24933 VGND.n2083 VGND.n2082 0.0845
R24934 VGND.n2085 VGND.n2084 0.0845
R24935 VGND.n2157 VGND.n2156 0.0845
R24936 VGND.n2155 VGND.n2154 0.0845
R24937 VGND.n2153 VGND.n2152 0.0845
R24938 VGND.n2151 VGND.n2150 0.0845
R24939 VGND.n2149 VGND.n2148 0.0845
R24940 VGND.n2147 VGND.n2146 0.0845
R24941 VGND.n2145 VGND.n2144 0.0845
R24942 VGND.n2139 VGND.n2138 0.0845
R24943 VGND.n2137 VGND.n2136 0.0845
R24944 VGND.n2135 VGND.n2134 0.0845
R24945 VGND.n2130 VGND.n2129 0.0845
R24946 VGND.n2128 VGND.n2127 0.0845
R24947 VGND.n2126 VGND.n2125 0.0845
R24948 VGND.n2121 VGND.n2120 0.0845
R24949 VGND.n2119 VGND.n2118 0.0845
R24950 VGND.n2117 VGND.n2116 0.0845
R24951 VGND.n2113 VGND.n2112 0.0845
R24952 VGND.n2111 VGND.n2110 0.0845
R24953 VGND.n2109 VGND.n2108 0.0845
R24954 VGND.n2107 VGND.n2106 0.0845
R24955 VGND.n2104 VGND.n2103 0.0845
R24956 VGND.n2102 VGND.n2101 0.0845
R24957 VGND.n2100 VGND.n2099 0.0845
R24958 VGND.n2098 VGND.n2097 0.0845
R24959 VGND.n3340 VGND.n3339 0.0845
R24960 VGND.n3342 VGND.n3341 0.0845
R24961 VGND.n3344 VGND.n3343 0.0845
R24962 VGND.n3346 VGND.n3345 0.0845
R24963 VGND.n3735 VGND 0.0845
R24964 VGND.n1921 VGND 0.08375
R24965 VGND VGND.n1303 0.083
R24966 VGND.n2644 VGND 0.083
R24967 VGND VGND.n3347 0.083
R24968 VGND VGND.n1376 0.08225
R24969 VGND.n257 VGND 0.08225
R24970 VGND VGND.n1979 0.08225
R24971 VGND.n3683 VGND.n3465 0.0815
R24972 VGND.n3667 VGND.n3666 0.0815
R24973 VGND.n3648 VGND.n3638 0.0815
R24974 VGND.n3663 VGND.n3653 0.0815
R24975 VGND.n3479 VGND.n3478 0.0815
R24976 VGND.n3585 VGND.n3571 0.0815
R24977 VGND.n3617 VGND.n3603 0.0815
R24978 VGND.n3633 VGND.n3619 0.0815
R24979 VGND.n3601 VGND.n3587 0.0815
R24980 VGND.n3569 VGND.n3555 0.0815
R24981 VGND.n3553 VGND.n3543 0.0815
R24982 VGND.n3714 VGND.n20 0.0815
R24983 VGND.n35 VGND.n34 0.0815
R24984 VGND.n3508 VGND.n3498 0.0815
R24985 VGND.n3523 VGND.n3513 0.0815
R24986 VGND.n3538 VGND.n3528 0.0815
R24987 VGND VGND.n933 0.0815
R24988 VGND VGND.n163 0.0815
R24989 VGND.n1282 VGND.n1281 0.0815
R24990 VGND VGND.n1378 0.0815
R24991 VGND VGND.n1511 0.0815
R24992 VGND VGND.n1666 0.0815
R24993 VGND.n1112 VGND.n1111 0.0815
R24994 VGND VGND.n2404 0.0815
R24995 VGND.n1482 VGND.n1481 0.08075
R24996 VGND.n1378 VGND 0.08
R24997 VGND.n1511 VGND 0.08
R24998 VGND VGND.n1670 0.08
R24999 VGND.n1176 VGND.n1175 0.08
R25000 VGND.n1165 VGND.n1164 0.08
R25001 VGND.n1158 VGND.n1157 0.08
R25002 VGND.n1085 VGND.n1084 0.08
R25003 VGND.n1081 VGND.n1080 0.08
R25004 VGND.n2236 VGND.n2235 0.08
R25005 VGND.n2240 VGND.n2239 0.08
R25006 VGND.n2526 VGND.n2525 0.08
R25007 VGND.n1063 VGND.n1062 0.08
R25008 VGND.n2011 VGND.n2010 0.08
R25009 VGND.n1955 VGND.n1954 0.0785
R25010 VGND.n634 VGND.n633 0.0785
R25011 VGND VGND.n3444 0.0755
R25012 VGND.n1394 VGND.n1393 0.0755
R25013 VGND.n1431 VGND 0.07475
R25014 VGND.n135 VGND 0.07475
R25015 VGND.n1626 VGND 0.07475
R25016 VGND.n1516 VGND 0.07475
R25017 VGND.n1080 VGND 0.07475
R25018 VGND VGND.n2240 0.07475
R25019 VGND VGND.n831 0.0725
R25020 VGND.n1414 VGND.n1413 0.0725
R25021 VGND.n174 VGND 0.0725
R25022 VGND.n189 VGND.n188 0.0725
R25023 VGND VGND.n184 0.0725
R25024 VGND.n224 VGND.n223 0.0725
R25025 VGND VGND.n1312 0.0725
R25026 VGND.n1595 VGND.n886 0.0725
R25027 VGND.n1593 VGND 0.0725
R25028 VGND.n1397 VGND.n1396 0.0725
R25029 VGND VGND.n3420 0.0725
R25030 VGND VGND.n1599 0.0725
R25031 VGND VGND.n1515 0.0725
R25032 VGND.n1700 VGND 0.0725
R25033 VGND VGND.n1777 0.0725
R25034 VGND VGND.n1747 0.0725
R25035 VGND VGND.n1967 0.0725
R25036 VGND.n761 VGND.n760 0.0725
R25037 VGND.n1803 VGND 0.0725
R25038 VGND.n1806 VGND.n1805 0.0725
R25039 VGND VGND.n639 0.0725
R25040 VGND.n952 VGND.n951 0.0725
R25041 VGND.n2398 VGND.n2397 0.0725
R25042 VGND.n2177 VGND.n482 0.0725
R25043 VGND.n2186 VGND 0.0725
R25044 VGND.n2883 VGND.n2882 0.0725
R25045 VGND.n2787 VGND.n2786 0.0725
R25046 VGND.n2887 VGND.n2886 0.0725
R25047 VGND.n2041 VGND.n2040 0.0725
R25048 VGND.n2052 VGND.n2051 0.0725
R25049 VGND.n2082 VGND 0.0725
R25050 VGND.n3103 VGND.n3102 0.0725
R25051 VGND.n916 VGND.n915 0.07175
R25052 VGND.n1190 VGND 0.07175
R25053 VGND VGND.n934 0.07025
R25054 VGND.n73 VGND 0.07025
R25055 VGND VGND.n109 0.07025
R25056 VGND VGND.n1592 0.07025
R25057 VGND.n307 VGND 0.07025
R25058 VGND.n1236 VGND 0.07025
R25059 VGND VGND.n1158 0.07025
R25060 VGND.n1154 VGND 0.07025
R25061 VGND VGND.n1144 0.07025
R25062 VGND VGND.n1129 0.07025
R25063 VGND VGND.n1106 0.07025
R25064 VGND VGND.n997 0.07025
R25065 VGND VGND.n963 0.07025
R25066 VGND VGND.n2428 0.07025
R25067 VGND.n2242 VGND 0.07025
R25068 VGND.n2518 VGND 0.07025
R25069 VGND.n2070 VGND 0.07025
R25070 VGND VGND.n1590 0.0695
R25071 VGND.n3431 VGND 0.0695
R25072 VGND.n1764 VGND.n1763 0.0695
R25073 VGND VGND.n756 0.0695
R25074 VGND.n1297 VGND.n1296 0.06875
R25075 VGND.n1471 VGND 0.06875
R25076 VGND VGND.n2184 0.06875
R25077 VGND.n1296 VGND.n1295 0.0665
R25078 VGND.n1398 VGND.n1397 0.0665
R25079 VGND VGND.n1276 0.06575
R25080 VGND VGND.n1201 0.06575
R25081 VGND.n1269 VGND 0.065
R25082 VGND.n1529 VGND.n1528 0.0635
R25083 VGND.n1674 VGND 0.0635
R25084 VGND.n1479 VGND.n1478 0.06275
R25085 VGND.n2057 VGND.n2056 0.06125
R25086 VGND.n934 VGND 0.0605
R25087 VGND.n128 VGND.n127 0.0605
R25088 VGND.n126 VGND.n125 0.0605
R25089 VGND.n239 VGND.n238 0.0605
R25090 VGND.n231 VGND.n230 0.0605
R25091 VGND.n72 VGND.n71 0.0605
R25092 VGND.n109 VGND 0.0605
R25093 VGND.n1306 VGND.n1305 0.0605
R25094 VGND.n1320 VGND.n1319 0.0605
R25095 VGND.n1592 VGND 0.0605
R25096 VGND VGND.n307 0.0605
R25097 VGND VGND.n314 0.0605
R25098 VGND.n1603 VGND.n1602 0.0605
R25099 VGND.n1547 VGND.n1546 0.0605
R25100 VGND.n3383 VGND.n3382 0.0605
R25101 VGND.n1645 VGND.n1644 0.0605
R25102 VGND.n1708 VGND.n1707 0.0605
R25103 VGND.n1710 VGND.n1709 0.0605
R25104 VGND.n1119 VGND.n1118 0.0605
R25105 VGND.n1180 VGND 0.0605
R25106 VGND.n1148 VGND.n1147 0.0605
R25107 VGND.n1142 VGND 0.0605
R25108 VGND.n1129 VGND 0.0605
R25109 VGND.n1962 VGND.n1961 0.0605
R25110 VGND.n1071 VGND.n1070 0.0605
R25111 VGND.n1099 VGND.n1098 0.0605
R25112 VGND.n628 VGND.n627 0.0605
R25113 VGND.n1912 VGND.n1911 0.0605
R25114 VGND.n997 VGND 0.0605
R25115 VGND.n972 VGND.n971 0.0605
R25116 VGND.n968 VGND.n967 0.0605
R25117 VGND.n963 VGND 0.0605
R25118 VGND.n459 VGND.n458 0.0605
R25119 VGND.n510 VGND 0.0605
R25120 VGND.n1020 VGND 0.0605
R25121 VGND.n1049 VGND 0.0605
R25122 VGND.n1035 VGND 0.0605
R25123 VGND.n2032 VGND.n2031 0.0605
R25124 VGND VGND.n2070 0.0605
R25125 VGND.n3275 VGND 0.0605
R25126 VGND.n95 VGND.n94 0.05975
R25127 VGND.n1588 VGND.n1587 0.05975
R25128 VGND.n1209 VGND.n1208 0.05975
R25129 VGND.n2046 VGND.n2045 0.05975
R25130 VGND.n902 VGND 0.059
R25131 VGND VGND.n1264 0.059
R25132 VGND.n1200 VGND 0.059
R25133 VGND.n1196 VGND 0.059
R25134 VGND VGND.n1195 0.059
R25135 VGND VGND.n1237 0.059
R25136 VGND VGND.n1234 0.059
R25137 VGND.n1121 VGND 0.059
R25138 VGND.n1171 VGND 0.059
R25139 VGND VGND.n1170 0.059
R25140 VGND.n2238 VGND 0.059
R25141 VGND VGND.n2519 0.059
R25142 VGND VGND.n1043 0.059
R25143 VGND.n1033 VGND 0.059
R25144 VGND.n1028 VGND 0.059
R25145 VGND VGND.n1027 0.059
R25146 VGND VGND.n574 0.059
R25147 VGND.n926 VGND.n925 0.0575
R25148 VGND.n853 VGND.n852 0.0575
R25149 VGND.n855 VGND.n854 0.0575
R25150 VGND.n1432 VGND.n1431 0.0575
R25151 VGND.n162 VGND.n60 0.0575
R25152 VGND VGND.n1317 0.0575
R25153 VGND.n297 VGND 0.0575
R25154 VGND.n298 VGND 0.0575
R25155 VGND.n1768 VGND.n1767 0.0575
R25156 VGND.n1164 VGND 0.0575
R25157 VGND.n1128 VGND 0.0575
R25158 VGND.n756 VGND 0.0575
R25159 VGND.n1818 VGND 0.0575
R25160 VGND.n1112 VGND 0.0575
R25161 VGND.n1910 VGND 0.0575
R25162 VGND.n1013 VGND 0.0575
R25163 VGND.n2188 VGND.n2187 0.0575
R25164 VGND.n2220 VGND 0.0575
R25165 VGND.n2599 VGND.n2598 0.0575
R25166 VGND.n2733 VGND.n2732 0.0575
R25167 VGND.n2729 VGND.n2728 0.0575
R25168 VGND.n435 VGND 0.0575
R25169 VGND.n2487 VGND 0.0575
R25170 VGND.n1066 VGND.n1065 0.0575
R25171 VGND VGND.n2011 0.0575
R25172 VGND VGND.n2079 0.0575
R25173 VGND VGND.n550 0.0575
R25174 VGND.n1452 VGND.n845 0.05675
R25175 VGND.n1819 VGND.n1818 0.05675
R25176 VGND.n931 VGND.n930 0.056
R25177 VGND.n179 VGND.n178 0.056
R25178 VGND.n3461 VGND 0.056
R25179 VGND.n1234 VGND.n1233 0.056
R25180 VGND.n1647 VGND.n1646 0.056
R25181 VGND.n1851 VGND 0.056
R25182 VGND.n1097 VGND.n1096 0.056
R25183 VGND.n1998 VGND.n1997 0.056
R25184 VGND.n1996 VGND.n1995 0.056
R25185 VGND.n1888 VGND 0.056
R25186 VGND.n712 VGND 0.056
R25187 VGND.n694 VGND 0.056
R25188 VGND.n2588 VGND 0.056
R25189 VGND.n2570 VGND 0.056
R25190 VGND VGND.n2839 0.056
R25191 VGND.n2861 VGND 0.056
R25192 VGND VGND.n2743 0.056
R25193 VGND.n2765 VGND 0.056
R25194 VGND.n2812 VGND 0.056
R25195 VGND.n2794 VGND 0.056
R25196 VGND.n2700 VGND 0.056
R25197 VGND.n2435 VGND.n2434 0.056
R25198 VGND.n2433 VGND.n2432 0.056
R25199 VGND VGND.n2267 0.056
R25200 VGND VGND.n2285 0.056
R25201 VGND VGND.n2304 0.056
R25202 VGND.n2330 VGND 0.056
R25203 VGND.n2551 VGND 0.056
R25204 VGND VGND.n2894 0.056
R25205 VGND.n2015 VGND.n2014 0.056
R25206 VGND.n2017 VGND.n2016 0.056
R25207 VGND.n2143 VGND 0.056
R25208 VGND.n2972 VGND 0.056
R25209 VGND.n3062 VGND 0.056
R25210 VGND.n3078 VGND 0.056
R25211 VGND.n3166 VGND 0.056
R25212 VGND.n3184 VGND 0.056
R25213 VGND.n3294 VGND 0.056
R25214 VGND.n17 VGND 0.056
R25215 VGND.n3678 VGND 0.05525
R25216 VGND.n3490 VGND 0.05525
R25217 VGND.n3643 VGND 0.05525
R25218 VGND.n3658 VGND 0.05525
R25219 VGND.n3473 VGND 0.05525
R25220 VGND.n3580 VGND 0.05525
R25221 VGND.n3612 VGND 0.05525
R25222 VGND.n3628 VGND 0.05525
R25223 VGND.n3596 VGND 0.05525
R25224 VGND.n3564 VGND 0.05525
R25225 VGND.n3548 VGND 0.05525
R25226 VGND.n3709 VGND 0.05525
R25227 VGND.n29 VGND 0.05525
R25228 VGND.n3503 VGND 0.05525
R25229 VGND.n3518 VGND 0.05525
R25230 VGND.n3533 VGND 0.05525
R25231 VGND.n874 VGND 0.05525
R25232 VGND VGND.n1416 0.05525
R25233 VGND.n3457 VGND 0.05525
R25234 VGND VGND.n341 0.05525
R25235 VGND.n351 VGND 0.05525
R25236 VGND.n3693 VGND 0.05525
R25237 VGND.n48 VGND 0.05525
R25238 VGND VGND.n264 0.05525
R25239 VGND.n1677 VGND 0.05525
R25240 VGND.n3364 VGND 0.05525
R25241 VGND.n1137 VGND 0.05525
R25242 VGND.n1861 VGND 0.05525
R25243 VGND.n1828 VGND 0.05525
R25244 VGND.n1092 VGND 0.05525
R25245 VGND.n671 VGND 0.05525
R25246 VGND.n1003 VGND 0.05525
R25247 VGND.n1001 VGND 0.05525
R25248 VGND.n2212 VGND 0.05525
R25249 VGND.n2598 VGND 0.05525
R25250 VGND.n2867 VGND 0.05525
R25251 VGND.n2619 VGND 0.05525
R25252 VGND.n2608 VGND 0.05525
R25253 VGND VGND.n395 0.05525
R25254 VGND.n2959 VGND 0.05525
R25255 VGND VGND.n2733 0.05525
R25256 VGND.n2771 VGND 0.05525
R25257 VGND.n2728 VGND 0.05525
R25258 VGND.n2725 VGND 0.05525
R25259 VGND.n2707 VGND 0.05525
R25260 VGND.n2689 VGND 0.05525
R25261 VGND.n2672 VGND 0.05525
R25262 VGND.n2653 VGND 0.05525
R25263 VGND.n2639 VGND 0.05525
R25264 VGND VGND.n445 0.05525
R25265 VGND VGND.n446 0.05525
R25266 VGND.n2418 VGND 0.05525
R25267 VGND VGND.n502 0.05525
R25268 VGND.n536 VGND 0.05525
R25269 VGND.n2473 VGND 0.05525
R25270 VGND.n2470 VGND 0.05525
R25271 VGND VGND.n2256 0.05525
R25272 VGND.n2337 VGND 0.05525
R25273 VGND.n2544 VGND 0.05525
R25274 VGND.n2509 VGND 0.05525
R25275 VGND.n2508 VGND 0.05525
R25276 VGND.n2498 VGND 0.05525
R25277 VGND VGND.n2899 0.05525
R25278 VGND VGND.n2914 0.05525
R25279 VGND.n2946 VGND 0.05525
R25280 VGND.n2937 VGND 0.05525
R25281 VGND.n2927 VGND 0.05525
R25282 VGND.n2150 VGND 0.05525
R25283 VGND.n2115 VGND 0.05525
R25284 VGND.n2097 VGND 0.05525
R25285 VGND VGND.n3352 0.05525
R25286 VGND.n2991 VGND 0.05525
R25287 VGND.n2987 VGND 0.05525
R25288 VGND.n2973 VGND 0.05525
R25289 VGND VGND.n3055 0.05525
R25290 VGND.n3065 VGND 0.05525
R25291 VGND.n3093 VGND 0.05525
R25292 VGND.n3080 VGND 0.05525
R25293 VGND VGND.n3158 0.05525
R25294 VGND.n3171 VGND 0.05525
R25295 VGND.n3199 VGND 0.05525
R25296 VGND.n3187 VGND 0.05525
R25297 VGND VGND.n3285 0.05525
R25298 VGND.n3301 VGND 0.05525
R25299 VGND.n3328 VGND 0.05525
R25300 VGND.n3317 VGND 0.05525
R25301 VGND.n3745 VGND 0.05525
R25302 VGND.n3727 VGND 0.05525
R25303 VGND.n13 VGND 0.05525
R25304 VGND VGND.n3009 0.05525
R25305 VGND.n3014 VGND 0.05525
R25306 VGND.n3032 VGND 0.05525
R25307 VGND.n3023 VGND 0.05525
R25308 VGND VGND.n3113 0.05525
R25309 VGND.n3119 VGND 0.05525
R25310 VGND.n3137 VGND 0.05525
R25311 VGND.n3128 VGND 0.05525
R25312 VGND VGND.n3218 0.05525
R25313 VGND.n3225 VGND 0.05525
R25314 VGND.n3266 VGND 0.05525
R25315 VGND.n3257 VGND 0.05525
R25316 VGND.n3247 VGND 0.05525
R25317 VGND.n3238 VGND 0.05525
R25318 VGND VGND.n3762 0.05525
R25319 VGND.n3771 VGND 0.05525
R25320 VGND.n3782 VGND 0.05525
R25321 VGND.n3672 VGND 0.0545
R25322 VGND.n3671 VGND 0.0545
R25323 VGND VGND.n3483 0.0545
R25324 VGND VGND.n3484 0.0545
R25325 VGND VGND.n3635 0.0545
R25326 VGND VGND.n3636 0.0545
R25327 VGND VGND.n3650 0.0545
R25328 VGND VGND.n3651 0.0545
R25329 VGND VGND.n3466 0.0545
R25330 VGND VGND.n3467 0.0545
R25331 VGND.n3574 VGND 0.0545
R25332 VGND.n3573 VGND 0.0545
R25333 VGND.n3606 VGND 0.0545
R25334 VGND.n3605 VGND 0.0545
R25335 VGND.n3622 VGND 0.0545
R25336 VGND.n3621 VGND 0.0545
R25337 VGND.n3590 VGND 0.0545
R25338 VGND.n3589 VGND 0.0545
R25339 VGND.n3558 VGND 0.0545
R25340 VGND.n3557 VGND 0.0545
R25341 VGND VGND.n3540 0.0545
R25342 VGND VGND.n3541 0.0545
R25343 VGND.n3703 VGND 0.0545
R25344 VGND.n3702 VGND 0.0545
R25345 VGND VGND.n22 0.0545
R25346 VGND VGND.n23 0.0545
R25347 VGND VGND.n3495 0.0545
R25348 VGND VGND.n3496 0.0545
R25349 VGND VGND.n3510 0.0545
R25350 VGND VGND.n3511 0.0545
R25351 VGND VGND.n3525 0.0545
R25352 VGND VGND.n3526 0.0545
R25353 VGND VGND.n3436 0.0545
R25354 VGND.n136 VGND.n135 0.0545
R25355 VGND VGND.n126 0.0545
R25356 VGND.n191 VGND 0.0545
R25357 VGND.n186 VGND 0.0545
R25358 VGND VGND.n214 0.0545
R25359 VGND VGND.n220 0.0545
R25360 VGND.n236 VGND 0.0545
R25361 VGND.n233 VGND 0.0545
R25362 VGND.n230 VGND 0.0545
R25363 VGND VGND.n62 0.0545
R25364 VGND VGND.n68 0.0545
R25365 VGND VGND.n72 0.0545
R25366 VGND VGND.n74 0.0545
R25367 VGND VGND.n87 0.0545
R25368 VGND VGND.n92 0.0545
R25369 VGND VGND.n95 0.0545
R25370 VGND.n107 VGND 0.0545
R25371 VGND.n99 VGND 0.0545
R25372 VGND VGND.n1306 0.0545
R25373 VGND VGND.n1325 0.0545
R25374 VGND VGND.n1328 0.0545
R25375 VGND.n1571 VGND 0.0545
R25376 VGND VGND.n1383 0.0545
R25377 VGND VGND.n299 0.0545
R25378 VGND VGND.n301 0.0545
R25379 VGND VGND.n304 0.0545
R25380 VGND VGND.n305 0.0545
R25381 VGND VGND.n329 0.0545
R25382 VGND VGND.n334 0.0545
R25383 VGND VGND.n339 0.0545
R25384 VGND.n3688 VGND 0.0545
R25385 VGND.n1260 VGND 0.0545
R25386 VGND.n1259 VGND 0.0545
R25387 VGND.n1253 VGND 0.0545
R25388 VGND.n1618 VGND 0.0545
R25389 VGND.n1616 VGND 0.0545
R25390 VGND.n1612 VGND 0.0545
R25391 VGND.n1605 VGND 0.0545
R25392 VGND VGND.n1464 0.0545
R25393 VGND.n1477 VGND 0.0545
R25394 VGND.n1558 VGND 0.0545
R25395 VGND.n1551 VGND 0.0545
R25396 VGND.n1536 VGND 0.0545
R25397 VGND.n1503 VGND 0.0545
R25398 VGND.n3403 VGND 0.0545
R25399 VGND VGND.n3389 0.0545
R25400 VGND VGND.n3383 0.0545
R25401 VGND.n3381 VGND 0.0545
R25402 VGND VGND.n208 0.0545
R25403 VGND.n256 VGND.n255 0.0545
R25404 VGND VGND.n268 0.0545
R25405 VGND.n1216 VGND 0.0545
R25406 VGND VGND.n1633 0.0545
R25407 VGND VGND.n1636 0.0545
R25408 VGND.n1644 VGND 0.0545
R25409 VGND VGND.n1648 0.0545
R25410 VGND.n1695 VGND.n1694 0.0545
R25411 VGND VGND.n1703 0.0545
R25412 VGND.n1704 VGND 0.0545
R25413 VGND.n1709 VGND 0.0545
R25414 VGND.n1714 VGND 0.0545
R25415 VGND.n1712 VGND 0.0545
R25416 VGND.n1711 VGND 0.0545
R25417 VGND.n1777 VGND 0.0545
R25418 VGND VGND.n1772 0.0545
R25419 VGND.n1761 VGND 0.0545
R25420 VGND VGND.n1752 0.0545
R25421 VGND.n1747 VGND 0.0545
R25422 VGND.n1745 VGND 0.0545
R25423 VGND.n3372 VGND 0.0545
R25424 VGND.n1188 VGND 0.0545
R25425 VGND.n1186 VGND 0.0545
R25426 VGND.n1182 VGND 0.0545
R25427 VGND.n1178 VGND 0.0545
R25428 VGND.n1167 VGND 0.0545
R25429 VGND.n1140 VGND 0.0545
R25430 VGND.n1136 VGND 0.0545
R25431 VGND.n1133 VGND 0.0545
R25432 VGND VGND.n1132 0.0545
R25433 VGND VGND.n762 0.0545
R25434 VGND VGND.n1796 0.0545
R25435 VGND VGND.n1801 0.0545
R25436 VGND VGND.n1809 0.0545
R25437 VGND.n1816 VGND 0.0545
R25438 VGND.n1872 VGND 0.0545
R25439 VGND.n1078 VGND 0.0545
R25440 VGND VGND.n626 0.0545
R25441 VGND.n630 VGND 0.0545
R25442 VGND.n1930 VGND 0.0545
R25443 VGND.n1919 VGND 0.0545
R25444 VGND.n1894 VGND 0.0545
R25445 VGND.n941 VGND 0.0545
R25446 VGND.n936 VGND 0.0545
R25447 VGND.n1012 VGND 0.0545
R25448 VGND.n1006 VGND 0.0545
R25449 VGND.n995 VGND 0.0545
R25450 VGND.n993 VGND 0.0545
R25451 VGND.n991 VGND 0.0545
R25452 VGND VGND.n990 0.0545
R25453 VGND.n989 VGND 0.0545
R25454 VGND VGND.n988 0.0545
R25455 VGND.n981 VGND 0.0545
R25456 VGND.n962 VGND 0.0545
R25457 VGND.n961 VGND 0.0545
R25458 VGND.n2399 VGND 0.0545
R25459 VGND VGND.n2395 0.0545
R25460 VGND VGND.n2182 0.0545
R25461 VGND VGND.n2189 0.0545
R25462 VGND VGND.n2200 0.0545
R25463 VGND VGND.n2219 0.0545
R25464 VGND VGND.n429 0.0545
R25465 VGND VGND.n434 0.0545
R25466 VGND VGND.n436 0.0545
R25467 VGND.n464 VGND 0.0545
R25468 VGND.n2444 VGND 0.0545
R25469 VGND.n2440 VGND 0.0545
R25470 VGND.n2439 VGND 0.0545
R25471 VGND.n2428 VGND 0.0545
R25472 VGND VGND.n493 0.0545
R25473 VGND.n515 VGND 0.0545
R25474 VGND.n2375 VGND 0.0545
R25475 VGND.n546 VGND 0.0545
R25476 VGND.n425 VGND 0.0545
R25477 VGND.n420 VGND 0.0545
R25478 VGND.n2486 VGND 0.0545
R25479 VGND.n2480 VGND 0.0545
R25480 VGND.n2462 VGND 0.0545
R25481 VGND VGND.n2224 0.0545
R25482 VGND VGND.n2244 0.0545
R25483 VGND VGND.n2245 0.0545
R25484 VGND.n2490 VGND 0.0545
R25485 VGND.n2555 VGND 0.0545
R25486 VGND.n2528 VGND 0.0545
R25487 VGND.n2513 VGND 0.0545
R25488 VGND.n1065 VGND 0.0545
R25489 VGND.n1058 VGND.n1057 0.0545
R25490 VGND VGND.n1054 0.0545
R25491 VGND.n1053 VGND 0.0545
R25492 VGND.n1037 VGND 0.0545
R25493 VGND.n1030 VGND.n1029 0.0545
R25494 VGND VGND.n2007 0.0545
R25495 VGND VGND.n2026 0.0545
R25496 VGND VGND.n2027 0.0545
R25497 VGND VGND.n2042 0.0545
R25498 VGND VGND.n2072 0.0545
R25499 VGND VGND.n2075 0.0545
R25500 VGND VGND.n2080 0.0545
R25501 VGND VGND.n2083 0.0545
R25502 VGND.n2090 VGND 0.0545
R25503 VGND VGND.n2164 0.0545
R25504 VGND.n2968 VGND 0.0545
R25505 VGND.n2967 VGND 0.0545
R25506 VGND.n2997 VGND 0.0545
R25507 VGND.n2985 VGND 0.0545
R25508 VGND.n3090 VGND 0.0545
R25509 VGND.n3195 VGND 0.0545
R25510 VGND.n3323 VGND 0.0545
R25511 VGND VGND.n381 0.0545
R25512 VGND VGND.n3002 0.0545
R25513 VGND.n818 VGND 0.05375
R25514 VGND.n835 VGND 0.05375
R25515 VGND VGND.n865 0.05375
R25516 VGND VGND.n2067 0.05375
R25517 VGND.n178 VGND.n177 0.053
R25518 VGND.n3410 VGND.n157 0.053
R25519 VGND VGND.n332 0.053
R25520 VGND.n1274 VGND 0.053
R25521 VGND.n1621 VGND.n1620 0.053
R25522 VGND.n1184 VGND 0.053
R25523 VGND.n1878 VGND.n720 0.053
R25524 VGND VGND.n2624 0.053
R25525 VGND.n2719 VGND 0.053
R25526 VGND.n2716 VGND 0.053
R25527 VGND.n2663 VGND 0.053
R25528 VGND.n2645 VGND 0.053
R25529 VGND.n1031 VGND 0.053
R25530 VGND VGND.n2034 0.053
R25531 VGND VGND.n2085 0.053
R25532 VGND.n2159 VGND 0.053
R25533 VGND.n2106 VGND 0.053
R25534 VGND VGND.n3346 0.053
R25535 VGND.n1676 VGND.n1675 0.05225
R25536 VGND.n933 VGND.n932 0.0515
R25537 VGND.n1439 VGND.n1438 0.0515
R25538 VGND.n1285 VGND.n1284 0.0515
R25539 VGND.n1115 VGND.n1114 0.0515
R25540 VGND.n1967 VGND.n1966 0.0515
R25541 VGND.n1953 VGND.n1952 0.0515
R25542 VGND.n2449 VGND.n426 0.0515
R25543 VGND.n2005 VGND.n2004 0.0515
R25544 VGND.n1313 VGND 0.05
R25545 VGND.n2077 VGND 0.04925
R25546 VGND.n885 VGND 0.0485
R25547 VGND.n1407 VGND.n1406 0.0485
R25548 VGND VGND.n3438 0.0485
R25549 VGND.n900 VGND 0.0485
R25550 VGND.n1567 VGND.n1566 0.0485
R25551 VGND.n1376 VGND 0.0485
R25552 VGND.n326 VGND.n325 0.0485
R25553 VGND VGND.n1272 0.0485
R25554 VGND.n1543 VGND 0.0485
R25555 VGND VGND.n257 0.0485
R25556 VGND.n1969 VGND 0.0485
R25557 VGND.n764 VGND.n763 0.0485
R25558 VGND.n1809 VGND.n1808 0.0485
R25559 VGND.n1989 VGND.n1988 0.0485
R25560 VGND.n1979 VGND 0.0485
R25561 VGND.n2409 VGND.n2408 0.0485
R25562 VGND VGND.n1019 0.0485
R25563 VGND VGND.n1041 0.0485
R25564 VGND.t4514 VGND.t3209 0.0481847
R25565 VGND.t102 VGND.t2010 0.0481847
R25566 VGND.t80 VGND.t34 0.0481847
R25567 VGND.t71 VGND.t5706 0.0481847
R25568 VGND.t199 VGND.t71 0.0481847
R25569 VGND.t38 VGND.t199 0.0481847
R25570 VGND.n3451 VGND.t38 0.0481847
R25571 VGND.t325 VGND.t108 0.0481847
R25572 VGND.t108 VGND.t3072 0.0481847
R25573 VGND.t6409 VGND.t3612 0.0481847
R25574 VGND.t3612 VGND.t2052 0.0481847
R25575 VGND.t2052 VGND.t139 0.0481847
R25576 VGND.t137 VGND.t6224 0.0481847
R25577 VGND.n1966 VGND 0.04775
R25578 VGND.n1560 VGND.n1443 0.047
R25579 VGND.n2297 VGND.n2296 0.047
R25580 VGND.n2916 VGND.n2915 0.047
R25581 VGND.n1470 VGND.n1469 0.04625
R25582 VGND.n1977 VGND 0.0455
R25583 VGND VGND.n1304 0.04475
R25584 VGND.n2643 VGND 0.04475
R25585 VGND VGND.n3348 0.04475
R25586 VGND.n1678 VGND.n1677 0.044
R25587 VGND.n1670 VGND 0.04325
R25588 VGND VGND.n1946 0.04325
R25589 VGND.n830 VGND.n829 0.0425
R25590 VGND VGND.n858 0.0425
R25591 VGND.n1434 VGND.n1433 0.0425
R25592 VGND.n243 VGND.n242 0.0425
R25593 VGND.n1595 VGND 0.0425
R25594 VGND.n1591 VGND 0.0425
R25595 VGND VGND.n1570 0.0425
R25596 VGND VGND.n1598 0.0425
R25597 VGND.n1460 VGND 0.0425
R25598 VGND.n1805 VGND 0.0425
R25599 VGND.n958 VGND 0.0425
R25600 VGND VGND.n2203 0.0425
R25601 VGND.n2371 VGND 0.0425
R25602 VGND.n2367 VGND 0.0425
R25603 VGND.n925 VGND 0.04175
R25604 VGND.n1767 VGND 0.04175
R25605 VGND.n1942 VGND.n1941 0.04175
R25606 VGND.n2037 VGND.n2036 0.04175
R25607 VGND VGND.n165 0.041
R25608 VGND VGND.n1470 0.041
R25609 VGND.n1472 VGND 0.041
R25610 VGND.n3400 VGND 0.041
R25611 VGND.n640 VGND 0.04025
R25612 VGND VGND.n80 0.0395
R25613 VGND VGND.n1531 0.0395
R25614 VGND.n1660 VGND.n1659 0.0395
R25615 VGND.n2179 VGND 0.0395
R25616 VGND.n3754 VGND 0.0395
R25617 VGND.n176 VGND.n175 0.03875
R25618 VGND.n314 VGND.n313 0.03875
R25619 VGND.n3387 VGND 0.03875
R25620 VGND.n836 VGND.n824 0.038
R25621 VGND.n1629 VGND.n838 0.038
R25622 VGND.n1632 VGND.n799 0.038
R25623 VGND.n983 VGND.n982 0.038
R25624 VGND.n2298 VGND.n2297 0.038
R25625 VGND VGND.n809 0.0365
R25626 VGND.n832 VGND 0.0365
R25627 VGND VGND.n172 0.0365
R25628 VGND.n190 VGND.n189 0.0365
R25629 VGND.n1578 VGND 0.0365
R25630 VGND.n319 VGND 0.0365
R25631 VGND VGND.n1552 0.0365
R25632 VGND.n1550 VGND.n1549 0.0365
R25633 VGND.n262 VGND.n261 0.0365
R25634 VGND.n1235 VGND 0.0365
R25635 VGND.n1653 VGND.n1652 0.0365
R25636 VGND.n1976 VGND 0.0365
R25637 VGND.n2380 VGND 0.0365
R25638 VGND VGND.n2377 0.0365
R25639 VGND.n1564 VGND.n1563 0.035
R25640 VGND.n3683 VGND.n3682 0.0335
R25641 VGND.n3666 VGND.n3494 0.0335
R25642 VGND.n3648 VGND.n3647 0.0335
R25643 VGND.n3663 VGND.n3662 0.0335
R25644 VGND.n3478 VGND.n3477 0.0335
R25645 VGND.n3585 VGND.n3584 0.0335
R25646 VGND.n3617 VGND.n3616 0.0335
R25647 VGND.n3633 VGND.n3632 0.0335
R25648 VGND.n3601 VGND.n3600 0.0335
R25649 VGND.n3569 VGND.n3568 0.0335
R25650 VGND.n3553 VGND.n3552 0.0335
R25651 VGND.n3714 VGND.n3713 0.0335
R25652 VGND.n34 VGND.n33 0.0335
R25653 VGND.n3508 VGND.n3507 0.0335
R25654 VGND.n3523 VGND.n3522 0.0335
R25655 VGND.n3538 VGND.n3537 0.0335
R25656 VGND.n875 VGND.n874 0.0335
R25657 VGND.n873 VGND.n872 0.0335
R25658 VGND.n1308 VGND.n1307 0.0335
R25659 VGND.n1383 VGND.n1382 0.0335
R25660 VGND.n1757 VGND.n1756 0.0335
R25661 VGND.n986 VGND.n985 0.0335
R25662 VGND.n2402 VGND.n2401 0.0335
R25663 VGND.n2388 VGND.n2387 0.0335
R25664 VGND.n2446 VGND.n428 0.0335
R25665 VGND.n1056 VGND.n1055 0.0335
R25666 VGND.n1052 VGND.n1051 0.0335
R25667 VGND.n2004 VGND.n574 0.0335
R25668 VGND.n1190 VGND.n1114 0.032
R25669 VGND.n1875 VGND.n721 0.032
R25670 VGND.n1103 VGND 0.032
R25671 VGND.n1879 VGND.n1878 0.032
R25672 VGND.n1066 VGND.n1015 0.032
R25673 VGND.n2133 VGND.n2132 0.032
R25674 VGND VGND.n3670 0.0305
R25675 VGND.n3485 VGND 0.0305
R25676 VGND.n3637 VGND 0.0305
R25677 VGND.n3652 VGND 0.0305
R25678 VGND.n3468 VGND 0.0305
R25679 VGND VGND.n3572 0.0305
R25680 VGND VGND.n3604 0.0305
R25681 VGND VGND.n3620 0.0305
R25682 VGND VGND.n3588 0.0305
R25683 VGND VGND.n3556 0.0305
R25684 VGND.n3542 VGND 0.0305
R25685 VGND VGND.n3701 0.0305
R25686 VGND.n24 VGND 0.0305
R25687 VGND.n3497 VGND 0.0305
R25688 VGND.n3512 VGND 0.0305
R25689 VGND.n3527 VGND 0.0305
R25690 VGND.n808 VGND.n57 0.0305
R25691 VGND.n854 VGND 0.0305
R25692 VGND VGND.n882 0.0305
R25693 VGND.n1430 VGND 0.0305
R25694 VGND.n3442 VGND 0.0305
R25695 VGND.n3439 VGND 0.0305
R25696 VGND.n139 VGND 0.0305
R25697 VGND.n133 VGND 0.0305
R25698 VGND VGND.n130 0.0305
R25699 VGND.n214 VGND.n213 0.0305
R25700 VGND.n215 VGND 0.0305
R25701 VGND.n64 VGND.n63 0.0305
R25702 VGND.n66 VGND 0.0305
R25703 VGND.n75 VGND 0.0305
R25704 VGND.n91 VGND 0.0305
R25705 VGND VGND.n103 0.0305
R25706 VGND.n3462 VGND.n3461 0.0305
R25707 VGND VGND.n1282 0.0305
R25708 VGND.n1283 VGND 0.0305
R25709 VGND VGND.n1286 0.0305
R25710 VGND.n1287 VGND 0.0305
R25711 VGND.n1292 VGND 0.0305
R25712 VGND VGND.n1321 0.0305
R25713 VGND.n1327 VGND 0.0305
R25714 VGND.n1332 VGND 0.0305
R25715 VGND VGND.n1333 0.0305
R25716 VGND.n1345 VGND 0.0305
R25717 VGND VGND.n1342 0.0305
R25718 VGND VGND.n1594 0.0305
R25719 VGND.n1584 VGND 0.0305
R25720 VGND.n1580 VGND 0.0305
R25721 VGND.n1388 VGND 0.0305
R25722 VGND.n1386 VGND 0.0305
R25723 VGND.n293 VGND 0.0305
R25724 VGND.n308 VGND 0.0305
R25725 VGND.n329 VGND 0.0305
R25726 VGND.n330 VGND 0.0305
R25727 VGND.n335 VGND 0.0305
R25728 VGND.n53 VGND.n52 0.0305
R25729 VGND VGND.n1268 0.0305
R25730 VGND VGND.n1258 0.0305
R25731 VGND VGND.n1250 0.0305
R25732 VGND.n1619 VGND 0.0305
R25733 VGND.n1611 VGND 0.0305
R25734 VGND.n1466 VGND 0.0305
R25735 VGND.n1521 VGND 0.0305
R25736 VGND VGND.n1503 0.0305
R25737 VGND VGND.n198 0.0305
R25738 VGND VGND.n1640 0.0305
R25739 VGND.n1648 VGND 0.0305
R25740 VGND.n1649 VGND 0.0305
R25741 VGND.n1664 VGND.n1663 0.0305
R25742 VGND VGND.n1697 0.0305
R25743 VGND VGND.n1776 0.0305
R25744 VGND VGND.n3375 0.0305
R25745 VGND VGND.n1120 0.0305
R25746 VGND.n1117 VGND 0.0305
R25747 VGND VGND.n1159 0.0305
R25748 VGND VGND.n1149 0.0305
R25749 VGND.n749 VGND 0.0305
R25750 VGND.n753 VGND 0.0305
R25751 VGND VGND.n1072 0.0305
R25752 VGND.n1069 VGND 0.0305
R25753 VGND.n1109 VGND 0.0305
R25754 VGND VGND.n1101 0.0305
R25755 VGND VGND.n1094 0.0305
R25756 VGND VGND.n1089 0.0305
R25757 VGND.n1087 VGND.n1086 0.0305
R25758 VGND VGND.n1929 0.0305
R25759 VGND.n1915 VGND.n1914 0.0305
R25760 VGND VGND.n1899 0.0305
R25761 VGND VGND.n941 0.0305
R25762 VGND VGND.n940 0.0305
R25763 VGND VGND.n1011 0.0305
R25764 VGND.n978 VGND.n977 0.0305
R25765 VGND VGND.n973 0.0305
R25766 VGND.n966 VGND 0.0305
R25767 VGND VGND.n961 0.0305
R25768 VGND.n2184 VGND.n2183 0.0305
R25769 VGND VGND.n2717 0.0305
R25770 VGND.n429 VGND 0.0305
R25771 VGND.n430 VGND 0.0305
R25772 VGND.n437 VGND 0.0305
R25773 VGND VGND.n460 0.0305
R25774 VGND.n457 VGND 0.0305
R25775 VGND.n453 VGND 0.0305
R25776 VGND.n2442 VGND.n2441 0.0305
R25777 VGND VGND.n2430 0.0305
R25778 VGND.n520 VGND.n519 0.0305
R25779 VGND VGND.n2356 0.0305
R25780 VGND VGND.n425 0.0305
R25781 VGND VGND.n424 0.0305
R25782 VGND VGND.n2485 0.0305
R25783 VGND VGND.n2479 0.0305
R25784 VGND VGND.n2460 0.0305
R25785 VGND.n2457 VGND 0.0305
R25786 VGND VGND.n2456 0.0305
R25787 VGND.n2453 VGND 0.0305
R25788 VGND.n2226 VGND 0.0305
R25789 VGND.n2228 VGND.n2227 0.0305
R25790 VGND.n2246 VGND 0.0305
R25791 VGND.n2535 VGND.n2534 0.0305
R25792 VGND VGND.n2516 0.0305
R25793 VGND.n2514 VGND.n2513 0.0305
R25794 VGND.n2502 VGND.n2501 0.0305
R25795 VGND.n2909 VGND.n2908 0.0305
R25796 VGND VGND.n2020 0.0305
R25797 VGND.n2039 VGND 0.0305
R25798 VGND.n2061 VGND.n2060 0.0305
R25799 VGND.n2072 VGND 0.0305
R25800 VGND.n2073 VGND 0.0305
R25801 VGND.n2080 VGND 0.0305
R25802 VGND.n2084 VGND 0.0305
R25803 VGND.n2992 VGND.n2991 0.0305
R25804 VGND.n2978 VGND.n2977 0.0305
R25805 VGND.n3058 VGND.n3057 0.0305
R25806 VGND.n3098 VGND.n3097 0.0305
R25807 VGND.n3085 VGND.n3084 0.0305
R25808 VGND.n3163 VGND.n3162 0.0305
R25809 VGND.n3204 VGND.n3203 0.0305
R25810 VGND.n3192 VGND.n3191 0.0305
R25811 VGND.n3292 VGND.n3291 0.0305
R25812 VGND.n3333 VGND.n3332 0.0305
R25813 VGND.n3322 VGND.n3321 0.0305
R25814 VGND.n3737 VGND.n3736 0.0305
R25815 VGND.n18 VGND.n17 0.0305
R25816 VGND VGND.n1576 0.02975
R25817 VGND.n1600 VGND 0.02975
R25818 VGND VGND.n2727 0.02975
R25819 VGND VGND.n2688 0.02975
R25820 VGND VGND.n2671 0.02975
R25821 VGND VGND.n2469 0.02975
R25822 VGND VGND.n2131 0.02975
R25823 VGND VGND.n2114 0.02975
R25824 VGND.n834 VGND 0.029
R25825 VGND.n1429 VGND 0.029
R25826 VGND.n905 VGND.n904 0.029
R25827 VGND.n907 VGND.n906 0.029
R25828 VGND VGND.n1335 0.029
R25829 VGND VGND.n302 0.029
R25830 VGND.n1271 VGND.n1270 0.029
R25831 VGND.n1232 VGND 0.029
R25832 VGND VGND.n1638 0.029
R25833 VGND.n1690 VGND.n1689 0.029
R25834 VGND.n1157 VGND.n1156 0.029
R25835 VGND.n1155 VGND.n1154 0.029
R25836 VGND.n1084 VGND.n1083 0.029
R25837 VGND.n1082 VGND.n1081 0.029
R25838 VGND.n1994 VGND 0.029
R25839 VGND.n1937 VGND.n1936 0.029
R25840 VGND VGND.n2699 0.029
R25841 VGND.n2231 VGND.n2230 0.029
R25842 VGND.n2233 VGND.n2232 0.029
R25843 VGND.n2235 VGND.n2234 0.029
R25844 VGND.n2531 VGND.n2530 0.029
R25845 VGND.n1018 VGND.n1017 0.029
R25846 VGND.n1062 VGND.n1061 0.029
R25847 VGND.n1060 VGND.n1059 0.029
R25848 VGND.n1040 VGND.n1039 0.029
R25849 VGND VGND.n2018 0.029
R25850 VGND VGND.n2047 0.029
R25851 VGND VGND.n2063 0.029
R25852 VGND VGND.n2068 0.029
R25853 VGND VGND.n2142 0.029
R25854 VGND.n935 VGND 0.0275
R25855 VGND.n924 VGND.n923 0.0275
R25856 VGND.n1380 VGND.n1379 0.0275
R25857 VGND.n1545 VGND.n1544 0.0275
R25858 VGND.n1523 VGND.n1522 0.0275
R25859 VGND.n1508 VGND.n1507 0.0275
R25860 VGND.n1238 VGND 0.0275
R25861 VGND VGND.n1771 0.0275
R25862 VGND VGND.n1128 0.0275
R25863 VGND.n2400 VGND.n2399 0.0275
R25864 VGND.n2599 VGND.n2559 0.0275
R25865 VGND.n2732 VGND.n418 0.0275
R25866 VGND.n2557 VGND.n2489 0.0275
R25867 VGND.n2089 VGND.n2088 0.0275
R25868 VGND.n2998 VGND.n2963 0.0275
R25869 VGND.n2055 VGND.n2054 0.02675
R25870 VGND.n3447 VGND 0.026
R25871 VGND.n1291 VGND 0.026
R25872 VGND VGND.n1322 0.026
R25873 VGND.n1116 VGND 0.026
R25874 VGND VGND.n1160 0.026
R25875 VGND VGND.n1146 0.026
R25876 VGND.n1145 VGND 0.026
R25877 VGND VGND.n1073 0.026
R25878 VGND.n1068 VGND 0.026
R25879 VGND.n1108 VGND 0.026
R25880 VGND VGND.n974 0.026
R25881 VGND VGND.n970 0.026
R25882 VGND.n969 VGND 0.026
R25883 VGND.n965 VGND 0.026
R25884 VGND VGND.n461 0.026
R25885 VGND.n456 VGND 0.026
R25886 VGND.n452 VGND 0.026
R25887 VGND.n2452 VGND 0.026
R25888 VGND.n2008 VGND 0.026
R25889 VGND VGND.n2021 0.026
R25890 VGND.n1576 VGND.n1575 0.02525
R25891 VGND VGND.n828 0.0245
R25892 VGND.n1420 VGND.n1419 0.0245
R25893 VGND.n1441 VGND.n1440 0.0245
R25894 VGND.n3435 VGND.n3434 0.0245
R25895 VGND.n140 VGND.n139 0.0245
R25896 VGND.n187 VGND.n186 0.0245
R25897 VGND VGND.n229 0.0245
R25898 VGND.n78 VGND.n77 0.0245
R25899 VGND.n82 VGND 0.0245
R25900 VGND VGND.n1288 0.0245
R25901 VGND.n1324 VGND 0.0245
R25902 VGND.n1342 VGND.n1341 0.0245
R25903 VGND.n1267 VGND.n1266 0.0245
R25904 VGND.n1519 VGND.n1518 0.0245
R25905 VGND.n1517 VGND.n1516 0.0245
R25906 VGND.n267 VGND 0.0245
R25907 VGND.n1198 VGND.n1197 0.0245
R25908 VGND.n1194 VGND.n1193 0.0245
R25909 VGND VGND.n1229 0.0245
R25910 VGND.n1697 VGND.n1696 0.0245
R25911 VGND.n1706 VGND 0.0245
R25912 VGND.n1787 VGND.n1786 0.0245
R25913 VGND.n1780 VGND.n1779 0.0245
R25914 VGND.n1750 VGND.n1749 0.0245
R25915 VGND.n1173 VGND.n1172 0.0245
R25916 VGND.n1959 VGND.n1958 0.0245
R25917 VGND.n1801 VGND.n1800 0.0245
R25918 VGND.n1812 VGND.n1811 0.0245
R25919 VGND.n1106 VGND.n1105 0.0245
R25920 VGND VGND.n1092 0.0245
R25921 VGND VGND.n1078 0.0245
R25922 VGND.n1914 VGND 0.0245
R25923 VGND.n2224 VGND 0.0245
R25924 VGND.n2522 VGND.n2521 0.0245
R25925 VGND.n1046 VGND.n1045 0.0245
R25926 VGND.n1026 VGND.n1025 0.0245
R25927 VGND.n2013 VGND 0.0245
R25928 VGND.n2059 VGND.n2058 0.0245
R25929 VGND VGND.n2090 0.0245
R25930 VGND.n2163 VGND.n2162 0.0245
R25931 VGND.n631 VGND.n630 0.02375
R25932 VGND.n2132 VGND 0.02375
R25933 VGND.n811 VGND.n810 0.023
R25934 VGND.n814 VGND.n813 0.023
R25935 VGND.n1633 VGND.n1632 0.023
R25936 VGND.n2828 VGND.n2827 0.023
R25937 VGND.n2824 VGND.n2823 0.023
R25938 VGND.n2692 VGND.n2691 0.023
R25939 VGND.n3044 VGND.n3043 0.023
R25940 VGND.n3040 VGND.n3039 0.023
R25941 VGND.n169 VGND 0.02225
R25942 VGND VGND.n922 0.0215
R25943 VGND.n1462 VGND.n1461 0.0215
R25944 VGND.n2220 VGND.n2169 0.0215
R25945 VGND.n866 VGND 0.02075
R25946 VGND.n317 VGND.n316 0.02075
R25947 VGND.n633 VGND 0.02075
R25948 VGND.n1290 VGND 0.02
R25949 VGND VGND.n1153 0.02
R25950 VGND.n2381 VGND.n485 0.02
R25951 VGND VGND.n908 0.01925
R25952 VGND.n3390 VGND 0.0185
R25953 VGND.n3377 VGND.n3376 0.0185
R25954 VGND.n1151 VGND.n1150 0.0185
R25955 VGND.n1842 VGND.n1841 0.0185
R25956 VGND.n2001 VGND.n2000 0.0185
R25957 VGND.n685 VGND.n684 0.0185
R25958 VGND VGND.n954 0.0185
R25959 VGND VGND.n2374 0.0185
R25960 VGND.n3273 VGND 0.017375
R25961 VGND.n3000 VGND 0.017375
R25962 VGND.n3041 VGND 0.017375
R25963 VGND.n3105 VGND 0.017375
R25964 VGND.n3145 VGND 0.017375
R25965 VGND.n3210 VGND 0.017375
R25966 VGND.n360 VGND 0.017375
R25967 VGND.n3716 VGND 0.017375
R25968 VGND.n3756 VGND 0.017375
R25969 VGND.n346 VGND.n345 0.017
R25970 VGND.n1540 VGND 0.017
R25971 VGND.n1150 VGND 0.017
R25972 VGND.n3754 VGND.n4 0.017
R25973 VGND.n3757 VGND.n2 0.017
R25974 VGND.n1598 VGND.n845 0.0155
R25975 VGND.n1657 VGND.n1656 0.0155
R25976 VGND.n2203 VGND.n2202 0.0155
R25977 VGND.n3682 VGND 0.01475
R25978 VGND.n3494 VGND 0.01475
R25979 VGND.n3647 VGND 0.01475
R25980 VGND.n3662 VGND 0.01475
R25981 VGND.n3477 VGND 0.01475
R25982 VGND.n3584 VGND 0.01475
R25983 VGND.n3616 VGND 0.01475
R25984 VGND.n3632 VGND 0.01475
R25985 VGND.n3600 VGND 0.01475
R25986 VGND.n3568 VGND 0.01475
R25987 VGND.n3552 VGND 0.01475
R25988 VGND.n3713 VGND 0.01475
R25989 VGND.n33 VGND 0.01475
R25990 VGND.n3507 VGND 0.01475
R25991 VGND.n3522 VGND 0.01475
R25992 VGND.n3537 VGND 0.01475
R25993 VGND.n3443 VGND 0.01475
R25994 VGND VGND.n79 0.01475
R25995 VGND.n1323 VGND 0.01475
R25996 VGND.n1340 VGND 0.01475
R25997 VGND.n312 VGND.n311 0.01475
R25998 VGND.n3690 VGND 0.01475
R25999 VGND.n1254 VGND 0.01475
R26000 VGND.n1606 VGND 0.01475
R26001 VGND.n3405 VGND 0.01475
R26002 VGND.n1715 VGND 0.01475
R26003 VGND.n3368 VGND 0.01475
R26004 VGND.n1138 VGND 0.01475
R26005 VGND.n1820 VGND 0.01475
R26006 VGND.n1832 VGND 0.01475
R26007 VGND.n675 VGND 0.01475
R26008 VGND.n1007 VGND 0.01475
R26009 VGND.n979 VGND 0.01475
R26010 VGND.n2216 VGND 0.01475
R26011 VGND.n2871 VGND 0.01475
R26012 VGND VGND.n2612 0.01475
R26013 VGND VGND.n2601 0.01475
R26014 VGND VGND.n390 0.01475
R26015 VGND.n387 VGND 0.01475
R26016 VGND.n2775 VGND 0.01475
R26017 VGND VGND.n441 0.01475
R26018 VGND.n2445 VGND 0.01475
R26019 VGND VGND.n492 0.01475
R26020 VGND.n540 VGND 0.01475
R26021 VGND.n2463 VGND 0.01475
R26022 VGND.n2341 VGND 0.01475
R26023 VGND.n2022 VGND 0.01475
R26024 VGND VGND.n2041 0.01475
R26025 VGND.n1563 VGND.n1400 0.014
R26026 VGND.n1434 VGND 0.0137353
R26027 VGND.n1301 VGND 0.0137353
R26028 VGND.n1531 VGND 0.0137353
R26029 VGND.n1873 VGND 0.0137353
R26030 VGND.n2190 VGND 0.0137353
R26031 VGND.n1281 VGND 0.01325
R26032 VGND VGND.n1315 0.01325
R26033 VGND.n3415 VGND.n3414 0.01325
R26034 VGND.n743 VGND 0.01325
R26035 VGND VGND.n884 0.0125
R26036 VGND.n880 VGND.n879 0.0125
R26037 VGND.n877 VGND.n876 0.0125
R26038 VGND.n1405 VGND 0.0125
R26039 VGND VGND.n173 0.0125
R26040 VGND.n193 VGND.n192 0.0125
R26041 VGND.n185 VGND 0.0125
R26042 VGND.n237 VGND 0.0125
R26043 VGND VGND.n1298 0.0125
R26044 VGND.n1314 VGND 0.0125
R26045 VGND.n1589 VGND 0.0125
R26046 VGND VGND.n1586 0.0125
R26047 VGND VGND.n1584 0.0125
R26048 VGND VGND.n1580 0.0125
R26049 VGND.n1399 VGND 0.0125
R26050 VGND.n1392 VGND 0.0125
R26051 VGND.n3430 VGND 0.0125
R26052 VGND.n3419 VGND 0.0125
R26053 VGND VGND.n157 0.0125
R26054 VGND.n292 VGND 0.0125
R26055 VGND VGND.n327 0.0125
R26056 VGND.n1623 VGND 0.0125
R26057 VGND.n1557 VGND 0.0125
R26058 VGND.n1544 VGND 0.0125
R26059 VGND.n1535 VGND 0.0125
R26060 VGND VGND.n1521 0.0125
R26061 VGND.n3392 VGND 0.0125
R26062 VGND.n3385 VGND 0.0125
R26063 VGND VGND.n266 0.0125
R26064 VGND VGND.n1650 0.0125
R26065 VGND.n1651 VGND 0.0125
R26066 VGND.n1680 VGND 0.0125
R26067 VGND.n1778 VGND 0.0125
R26068 VGND.n1759 VGND 0.0125
R26069 VGND.n1748 VGND 0.0125
R26070 VGND.n1743 VGND.n1742 0.0125
R26071 VGND.n1734 VGND 0.0125
R26072 VGND VGND.n1968 0.0125
R26073 VGND VGND.n1795 0.0125
R26074 VGND VGND.n1802 0.0125
R26075 VGND.n1821 VGND 0.0125
R26076 VGND VGND.n1990 0.0125
R26077 VGND VGND.n1986 0.0125
R26078 VGND.n1973 VGND.n1972 0.0125
R26079 VGND.n1901 VGND 0.0125
R26080 VGND VGND.n957 0.0125
R26081 VGND VGND.n952 0.0125
R26082 VGND.n2390 VGND 0.0125
R26083 VGND VGND.n2389 0.0125
R26084 VGND.n2200 VGND.n2199 0.0125
R26085 VGND.n2218 VGND 0.0125
R26086 VGND.n2414 VGND.n2413 0.0125
R26087 VGND VGND.n2379 0.0125
R26088 VGND.n2378 VGND 0.0125
R26089 VGND.n2358 VGND 0.0125
R26090 VGND.n2261 VGND.n2260 0.0125
R26091 VGND.n2040 VGND.n2039 0.0125
R26092 VGND VGND.n2059 0.0125
R26093 VGND VGND.n2076 0.0125
R26094 VGND.n2160 VGND 0.0125
R26095 VGND.n912 VGND 0.01175
R26096 VGND.n1946 VGND.n1945 0.011
R26097 VGND.n3335 VGND 0.011
R26098 VGND.n1337 VGND 0.01025
R26099 VGND VGND.n1343 0.01025
R26100 VGND.n1582 VGND.n1581 0.01025
R26101 VGND VGND.n838 0.01025
R26102 VGND.n2229 VGND 0.01025
R26103 VGND VGND.n2532 0.01025
R26104 VGND.n1665 VGND.n1664 0.0095
R26105 VGND.n1947 VGND 0.0095
R26106 VGND.n196 VGND.n179 0.008
R26107 VGND VGND.n2524 0.008
R26108 VGND.n883 VGND 0.0065
R26109 VGND.n1223 VGND 0.0065
R26110 VGND.n1662 VGND.n1661 0.0065
R26111 VGND VGND.n1760 0.0065
R26112 VGND.n1988 VGND 0.0065
R26113 VGND.n2404 VGND.n2403 0.0065
R26114 VGND VGND.n2392 0.0065
R26115 VGND.n2533 VGND 0.0065
R26116 VGND.n2066 VGND.n2065 0.0065
R26117 VGND VGND.n2071 0.0065
R26118 VGND.n265 VGND 0.00575
R26119 VGND.n1294 VGND.n1293 0.005
R26120 VGND.n1636 VGND.n1635 0.005
R26121 VGND.n1162 VGND.n1161 0.005
R26122 VGND.n1075 VGND.n1074 0.005
R26123 VGND.n1111 VGND.n1110 0.005
R26124 VGND.n976 VGND.n975 0.005
R26125 VGND.n463 VGND.n462 0.005
R26126 VGND.n455 VGND.n454 0.005
R26127 VGND.n451 VGND.n450 0.005
R26128 VGND.n2459 VGND.n2458 0.005
R26129 VGND.n2455 VGND.n2454 0.005
R26130 VGND.n2451 VGND.n2450 0.005
R26131 VGND VGND.n56 0.0035
R26132 VGND VGND.n921 0.0035
R26133 VGND VGND.n811 0.0035
R26134 VGND VGND.n814 0.0035
R26135 VGND.n851 VGND.n58 0.0035
R26136 VGND.n1436 VGND 0.0035
R26137 VGND.n3433 VGND.n140 0.0035
R26138 VGND.n217 VGND 0.0035
R26139 VGND VGND.n3452 0.0035
R26140 VGND.n1301 VGND 0.0035
R26141 VGND.n340 VGND 0.0035
R26142 VGND.n3691 VGND 0.0035
R26143 VGND.n1278 VGND.n1240 0.0035
R26144 VGND.n1249 VGND.n1248 0.0035
R26145 VGND.n1454 VGND 0.0035
R26146 VGND VGND.n1457 0.0035
R26147 VGND.n1554 VGND.n1553 0.0035
R26148 VGND.n3394 VGND.n3393 0.0035
R26149 VGND.n1693 VGND 0.0035
R26150 VGND.n1791 VGND.n1790 0.0035
R26151 VGND VGND.n1744 0.0035
R26152 VGND.n1951 VGND 0.0035
R26153 VGND.n759 VGND.n758 0.0035
R26154 VGND.n767 VGND.n766 0.0035
R26155 VGND VGND.n1804 0.0035
R26156 VGND.n2352 VGND.n547 0.0035
R26157 VGND.n2349 VGND.n2348 0.0035
R26158 VGND.n2911 VGND 0.0035
R26159 VGND.n3208 VGND.n3207 0.0035
R26160 VGND.n3212 VGND.n3211 0.0035
R26161 VGND.n80 VGND 0.00275
R26162 VGND VGND.n259 0.00275
R26163 VGND.n1754 VGND 0.00275
R26164 VGND VGND.n3465 0.002
R26165 VGND.n3667 VGND 0.002
R26166 VGND.n3638 VGND 0.002
R26167 VGND.n3653 VGND 0.002
R26168 VGND.n3479 VGND 0.002
R26169 VGND VGND.n3571 0.002
R26170 VGND VGND.n3603 0.002
R26171 VGND VGND.n3619 0.002
R26172 VGND VGND.n3587 0.002
R26173 VGND VGND.n3555 0.002
R26174 VGND.n3543 VGND 0.002
R26175 VGND VGND.n20 0.002
R26176 VGND.n35 VGND 0.002
R26177 VGND.n3498 VGND 0.002
R26178 VGND.n3513 VGND 0.002
R26179 VGND.n3528 VGND 0.002
R26180 VGND VGND.n929 0.002
R26181 VGND VGND.n57 0.002
R26182 VGND.n816 VGND 0.002
R26183 VGND VGND.n833 0.002
R26184 VGND VGND.n58 0.002
R26185 VGND.n858 VGND 0.002
R26186 VGND VGND.n881 0.002
R26187 VGND VGND.n59 0.002
R26188 VGND.n1409 VGND 0.002
R26189 VGND VGND.n1437 0.002
R26190 VGND.n3446 VGND 0.002
R26191 VGND VGND.n3445 0.002
R26192 VGND VGND.n136 0.002
R26193 VGND VGND.n60 0.002
R26194 VGND.n166 VGND 0.002
R26195 VGND VGND.n195 0.002
R26196 VGND.n213 VGND 0.002
R26197 VGND VGND.n240 0.002
R26198 VGND VGND.n61 0.002
R26199 VGND.n63 VGND 0.002
R26200 VGND.n81 VGND 0.002
R26201 VGND.n111 VGND 0.002
R26202 VGND VGND.n110 0.002
R26203 VGND.n3463 VGND 0.002
R26204 VGND VGND.n3462 0.002
R26205 VGND.n1289 VGND 0.002
R26206 VGND.n1303 VGND 0.002
R26207 VGND.n1304 VGND 0.002
R26208 VGND.n1318 VGND 0.002
R26209 VGND.n1336 VGND 0.002
R26210 VGND.n1347 VGND 0.002
R26211 VGND VGND.n1591 0.002
R26212 VGND VGND.n1574 0.002
R26213 VGND VGND.n1573 0.002
R26214 VGND VGND.n1398 0.002
R26215 VGND VGND.n1381 0.002
R26216 VGND VGND.n1377 0.002
R26217 VGND VGND.n3428 0.002
R26218 VGND VGND.n3418 0.002
R26219 VGND VGND.n3416 0.002
R26220 VGND.n290 VGND 0.002
R26221 VGND.n303 VGND 0.002
R26222 VGND.n306 VGND 0.002
R26223 VGND.n318 VGND 0.002
R26224 VGND.n333 VGND 0.002
R26225 VGND.n355 VGND 0.002
R26226 VGND.n3697 VGND 0.002
R26227 VGND.n3686 VGND 0.002
R26228 VGND VGND.n53 0.002
R26229 VGND VGND.n1273 0.002
R26230 VGND VGND.n1255 0.002
R26231 VGND VGND.n1625 0.002
R26232 VGND VGND.n1607 0.002
R26233 VGND.n1456 VGND 0.002
R26234 VGND.n1482 VGND 0.002
R26235 VGND VGND.n1554 0.002
R26236 VGND VGND.n1539 0.002
R26237 VGND VGND.n1526 0.002
R26238 VGND VGND.n1510 0.002
R26239 VGND VGND.n3399 0.002
R26240 VGND VGND.n3388 0.002
R26241 VGND.n258 VGND 0.002
R26242 VGND VGND.n1231 0.002
R26243 VGND VGND.n1217 0.002
R26244 VGND.n1639 VGND 0.002
R26245 VGND.n1654 VGND 0.002
R26246 VGND.n1671 VGND 0.002
R26247 VGND.n1684 VGND 0.002
R26248 VGND.n1694 VGND 0.002
R26249 VGND VGND.n1783 0.002
R26250 VGND VGND.n1769 0.002
R26251 VGND VGND.n1755 0.002
R26252 VGND VGND.n1741 0.002
R26253 VGND VGND.n3369 0.002
R26254 VGND VGND.n1163 0.002
R26255 VGND VGND.n1143 0.002
R26256 VGND VGND.n1130 0.002
R26257 VGND VGND.n1964 0.002
R26258 VGND VGND.n1948 0.002
R26259 VGND.n745 VGND 0.002
R26260 VGND.n758 VGND 0.002
R26261 VGND.n1799 VGND 0.002
R26262 VGND.n1822 VGND 0.002
R26263 VGND VGND.n1870 0.002
R26264 VGND VGND.n1852 0.002
R26265 VGND VGND.n1833 0.002
R26266 VGND VGND.n1104 0.002
R26267 VGND VGND.n1087 0.002
R26268 VGND VGND.n1993 0.002
R26269 VGND VGND.n1980 0.002
R26270 VGND.n629 VGND 0.002
R26271 VGND VGND.n644 0.002
R26272 VGND.n653 VGND 0.002
R26273 VGND VGND.n1931 0.002
R26274 VGND VGND.n1922 0.002
R26275 VGND VGND.n1905 0.002
R26276 VGND VGND.n1889 0.002
R26277 VGND VGND.n713 0.002
R26278 VGND VGND.n695 0.002
R26279 VGND VGND.n676 0.002
R26280 VGND VGND.n1008 0.002
R26281 VGND VGND.n998 0.002
R26282 VGND VGND.n978 0.002
R26283 VGND VGND.n958 0.002
R26284 VGND VGND.n2407 0.002
R26285 VGND VGND.n2393 0.002
R26286 VGND VGND.n2180 0.002
R26287 VGND.n2181 VGND 0.002
R26288 VGND VGND.n2589 0.002
R26289 VGND VGND.n2571 0.002
R26290 VGND.n2838 VGND 0.002
R26291 VGND.n2862 VGND 0.002
R26292 VGND VGND.n2872 0.002
R26293 VGND.n2742 VGND 0.002
R26294 VGND.n2766 VGND 0.002
R26295 VGND VGND.n2813 0.002
R26296 VGND VGND.n2795 0.002
R26297 VGND VGND.n2776 0.002
R26298 VGND.n2628 VGND 0.002
R26299 VGND VGND.n2718 0.002
R26300 VGND VGND.n2715 0.002
R26301 VGND VGND.n2698 0.002
R26302 VGND VGND.n2681 0.002
R26303 VGND VGND.n2662 0.002
R26304 VGND.n2662 VGND 0.002
R26305 VGND VGND.n2644 0.002
R26306 VGND VGND.n2643 0.002
R26307 VGND.n440 VGND 0.002
R26308 VGND.n465 VGND 0.002
R26309 VGND VGND.n2442 0.002
R26310 VGND VGND.n2427 0.002
R26311 VGND.n491 VGND 0.002
R26312 VGND.n520 VGND 0.002
R26313 VGND VGND.n2376 0.002
R26314 VGND VGND.n2362 0.002
R26315 VGND VGND.n541 0.002
R26316 VGND VGND.n2482 0.002
R26317 VGND VGND.n2464 0.002
R26318 VGND.n2227 VGND 0.002
R26319 VGND.n2247 VGND 0.002
R26320 VGND.n2266 VGND 0.002
R26321 VGND.n2284 VGND 0.002
R26322 VGND.n2303 VGND 0.002
R26323 VGND.n2331 VGND 0.002
R26324 VGND VGND.n2342 0.002
R26325 VGND VGND.n2552 0.002
R26326 VGND VGND.n2535 0.002
R26327 VGND VGND.n2533 0.002
R26328 VGND VGND.n2514 0.002
R26329 VGND VGND.n2504 0.002
R26330 VGND VGND.n2502 0.002
R26331 VGND.n2891 VGND 0.002
R26332 VGND.n2908 VGND 0.002
R26333 VGND.n2950 VGND 0.002
R26334 VGND VGND.n2941 0.002
R26335 VGND VGND.n2931 0.002
R26336 VGND VGND.n1058 0.002
R26337 VGND VGND.n1050 0.002
R26338 VGND VGND.n1030 0.002
R26339 VGND.n2012 VGND 0.002
R26340 VGND.n2019 VGND 0.002
R26341 VGND.n2035 VGND 0.002
R26342 VGND.n2044 VGND 0.002
R26343 VGND.n2048 VGND 0.002
R26344 VGND.n2060 VGND 0.002
R26345 VGND.n2069 VGND 0.002
R26346 VGND.n2071 VGND 0.002
R26347 VGND.n2091 VGND 0.002
R26348 VGND VGND.n2161 0.002
R26349 VGND VGND.n2158 0.002
R26350 VGND VGND.n2141 0.002
R26351 VGND VGND.n2124 0.002
R26352 VGND VGND.n2105 0.002
R26353 VGND.n2105 VGND 0.002
R26354 VGND.n3347 VGND 0.002
R26355 VGND.n3348 VGND 0.002
R26356 VGND VGND.n2992 0.002
R26357 VGND VGND.n2986 0.002
R26358 VGND VGND.n2978 0.002
R26359 VGND.n3047 VGND 0.002
R26360 VGND.n3057 VGND 0.002
R26361 VGND.n3073 VGND 0.002
R26362 VGND VGND.n3098 0.002
R26363 VGND VGND.n3091 0.002
R26364 VGND VGND.n3085 0.002
R26365 VGND.n3150 VGND 0.002
R26366 VGND.n3162 VGND 0.002
R26367 VGND.n3179 VGND 0.002
R26368 VGND VGND.n3204 0.002
R26369 VGND VGND.n3196 0.002
R26370 VGND VGND.n3192 0.002
R26371 VGND.n3277 VGND 0.002
R26372 VGND.n3291 VGND 0.002
R26373 VGND.n3309 VGND 0.002
R26374 VGND VGND.n3333 0.002
R26375 VGND VGND.n3324 0.002
R26376 VGND VGND.n3322 0.002
R26377 VGND VGND.n3753 0.002
R26378 VGND VGND.n3737 0.002
R26379 VGND VGND.n3735 0.002
R26380 VGND.n3718 VGND 0.002
R26381 VGND VGND.n18 0.002
R26382 VGND.n3005 VGND 0.002
R26383 VGND.n3018 VGND 0.002
R26384 VGND VGND.n3036 0.002
R26385 VGND VGND.n3027 0.002
R26386 VGND.n3109 VGND 0.002
R26387 VGND.n3123 VGND 0.002
R26388 VGND VGND.n3141 0.002
R26389 VGND VGND.n3132 0.002
R26390 VGND.n3214 VGND 0.002
R26391 VGND.n3229 VGND 0.002
R26392 VGND VGND.n3270 0.002
R26393 VGND VGND.n3261 0.002
R26394 VGND VGND.n3251 0.002
R26395 VGND VGND.n3242 0.002
R26396 VGND.n3758 VGND 0.002
R26397 VGND.n3775 VGND 0.002
R26398 VGND VGND.n0 0.002
R26399 VGND VGND.n3786 0.002
R26400 VGND.n1468 VGND.n1467 0.00125
R26401 VGND.n1940 VGND.n611 0.00125
R26402 VGND.n1925 VGND.n1924 0.00125
R26403 a_44296_24393.n13 a_44296_24393.t38 15.4765
R26404 a_44296_24393.n14 a_44296_24393.t36 15.4765
R26405 a_44296_24393.n15 a_44296_24393.t40 15.4765
R26406 a_44296_24393.n16 a_44296_24393.t14 15.4765
R26407 a_44296_24393.n17 a_44296_24393.t18 15.4765
R26408 a_44296_24393.n18 a_44296_24393.t23 15.4765
R26409 a_44296_24393.n19 a_44296_24393.t19 15.4765
R26410 a_44296_24393.n20 a_44296_24393.t24 15.4765
R26411 a_44296_24393.n21 a_44296_24393.t32 15.4765
R26412 a_44296_24393.n22 a_44296_24393.t28 15.4765
R26413 a_44296_24393.n23 a_44296_24393.t33 15.4765
R26414 a_44296_24393.n26 a_44296_24393.t29 15.4765
R26415 a_44296_24393.n10 a_44296_24393.t16 15.4765
R26416 a_44296_24393.n11 a_44296_24393.t42 15.4765
R26417 a_44296_24393.n12 a_44296_24393.t15 15.4765
R26418 a_44296_24393.n27 a_44296_24393.t41 15.4765
R26419 a_44296_24393.n13 a_44296_24393.t25 11.863
R26420 a_44296_24393.n14 a_44296_24393.t34 11.863
R26421 a_44296_24393.n15 a_44296_24393.t37 11.863
R26422 a_44296_24393.n16 a_44296_24393.t43 11.863
R26423 a_44296_24393.n17 a_44296_24393.t35 11.863
R26424 a_44296_24393.n18 a_44296_24393.t20 11.863
R26425 a_44296_24393.n19 a_44296_24393.t17 11.863
R26426 a_44296_24393.n20 a_44296_24393.t21 11.863
R26427 a_44296_24393.n21 a_44296_24393.t22 11.863
R26428 a_44296_24393.n22 a_44296_24393.t26 11.863
R26429 a_44296_24393.n10 a_44296_24393.t45 11.863
R26430 a_44296_24393.n11 a_44296_24393.t39 11.863
R26431 a_44296_24393.n12 a_44296_24393.t44 11.863
R26432 a_44296_24393.n27 a_44296_24393.t31 11.863
R26433 a_44296_24393.n24 a_44296_24393.t30 11.8022
R26434 a_44296_24393.n25 a_44296_24393.t27 11.8022
R26435 a_44296_24393.n7 a_44296_24393.t8 11.3584
R26436 a_44296_24393.n14 a_44296_24393.n13 10.5449
R26437 a_44296_24393.n15 a_44296_24393.n14 10.5449
R26438 a_44296_24393.n16 a_44296_24393.n15 10.5449
R26439 a_44296_24393.n17 a_44296_24393.n16 10.5449
R26440 a_44296_24393.n18 a_44296_24393.n17 10.5449
R26441 a_44296_24393.n19 a_44296_24393.n18 10.5449
R26442 a_44296_24393.n20 a_44296_24393.n19 10.5449
R26443 a_44296_24393.n21 a_44296_24393.n20 10.5449
R26444 a_44296_24393.n22 a_44296_24393.n21 10.5449
R26445 a_44296_24393.n23 a_44296_24393.n22 10.5449
R26446 a_44296_24393.n11 a_44296_24393.n10 10.5449
R26447 a_44296_24393.n12 a_44296_24393.n11 10.5449
R26448 a_44296_24393.n27 a_44296_24393.n12 10.5449
R26449 a_44296_24393.n27 a_44296_24393.n26 10.5449
R26450 a_44296_24393.n9 a_44296_24393.t1 10.4819
R26451 a_44296_24393.n25 a_44296_24393.n24 10.26
R26452 a_44296_24393.n8 a_44296_24393.n5 6.43746
R26453 a_44296_24393.n7 a_44296_24393.n6 6.43746
R26454 a_44296_24393.n3 a_44296_24393.n2 6.25311
R26455 a_44296_24393.n3 a_44296_24393.n1 5.37659
R26456 a_44296_24393.n4 a_44296_24393.n0 5.37659
R26457 a_44296_24393.n30 a_44296_24393.n29 5.37659
R26458 a_44296_24393.n5 a_44296_24393.t6 4.04494
R26459 a_44296_24393.n5 a_44296_24393.t3 4.04494
R26460 a_44296_24393.n6 a_44296_24393.t10 4.04494
R26461 a_44296_24393.n6 a_44296_24393.t9 4.04494
R26462 a_44296_24393.n2 a_44296_24393.t2 3.07367
R26463 a_44296_24393.n1 a_44296_24393.t4 3.07367
R26464 a_44296_24393.n0 a_44296_24393.t13 3.07367
R26465 a_44296_24393.t0 a_44296_24393.n30 3.07367
R26466 a_44296_24393.n2 a_44296_24393.t11 2.22001
R26467 a_44296_24393.n1 a_44296_24393.t5 2.22001
R26468 a_44296_24393.n0 a_44296_24393.t7 2.22001
R26469 a_44296_24393.n30 a_44296_24393.t12 2.22001
R26470 a_44296_24393.n28 a_44296_24393.n27 1.9195
R26471 a_44296_24393.n8 a_44296_24393.n7 0.877022
R26472 a_44296_24393.n9 a_44296_24393.n8 0.877022
R26473 a_44296_24393.n4 a_44296_24393.n3 0.877022
R26474 a_44296_24393.n29 a_44296_24393.n4 0.877022
R26475 a_44296_24393.n29 a_44296_24393.n28 0.430935
R26476 a_44296_24393.n28 a_44296_24393.n9 0.313543
R26477 a_44296_24393.n24 a_44296_24393.n23 0.0613333
R26478 a_44296_24393.n26 a_44296_24393.n25 0.0613333
R26479 clkbuf_1_0__f_clk.I.n6 clkbuf_1_0__f_clk.I.t33 31.7717
R26480 clkbuf_1_0__f_clk.I.n9 clkbuf_1_0__f_clk.I.t47 31.7717
R26481 clkbuf_1_0__f_clk.I.n3 clkbuf_1_0__f_clk.I.t56 29.7439
R26482 clkbuf_1_0__f_clk.I.n11 clkbuf_1_0__f_clk.I.t54 29.7439
R26483 clkbuf_1_0__f_clk.I.n6 clkbuf_1_0__f_clk.I.t40 18.7615
R26484 clkbuf_1_0__f_clk.I.n7 clkbuf_1_0__f_clk.I.t46 18.7615
R26485 clkbuf_1_0__f_clk.I.n3 clkbuf_1_0__f_clk.I.t59 18.7615
R26486 clkbuf_1_0__f_clk.I.n4 clkbuf_1_0__f_clk.I.t48 18.7615
R26487 clkbuf_1_0__f_clk.I.n5 clkbuf_1_0__f_clk.I.t51 18.7615
R26488 clkbuf_1_0__f_clk.I.n8 clkbuf_1_0__f_clk.I.t50 18.7615
R26489 clkbuf_1_0__f_clk.I.n11 clkbuf_1_0__f_clk.I.t57 18.7615
R26490 clkbuf_1_0__f_clk.I.n12 clkbuf_1_0__f_clk.I.t55 18.7615
R26491 clkbuf_1_0__f_clk.I.n13 clkbuf_1_0__f_clk.I.t39 18.7615
R26492 clkbuf_1_0__f_clk.I.n9 clkbuf_1_0__f_clk.I.t41 18.7615
R26493 clkbuf_1_0__f_clk.I.n10 clkbuf_1_0__f_clk.I.t34 18.7615
R26494 clkbuf_1_0__f_clk.I.n14 clkbuf_1_0__f_clk.I.t44 18.7615
R26495 clkbuf_1_0__f_clk.I.n15 clkbuf_1_0__f_clk.I 17.5834
R26496 clkbuf_1_0__f_clk.I.n11 clkbuf_1_0__f_clk.I.t35 11.133
R26497 clkbuf_1_0__f_clk.I.n12 clkbuf_1_0__f_clk.I.t32 11.133
R26498 clkbuf_1_0__f_clk.I.n13 clkbuf_1_0__f_clk.I.t36 11.133
R26499 clkbuf_1_0__f_clk.I.n9 clkbuf_1_0__f_clk.I.t49 11.133
R26500 clkbuf_1_0__f_clk.I.n10 clkbuf_1_0__f_clk.I.t45 11.133
R26501 clkbuf_1_0__f_clk.I.n14 clkbuf_1_0__f_clk.I.t52 11.133
R26502 clkbuf_1_0__f_clk.I.n6 clkbuf_1_0__f_clk.I.t58 11.0722
R26503 clkbuf_1_0__f_clk.I.n7 clkbuf_1_0__f_clk.I.t37 11.0722
R26504 clkbuf_1_0__f_clk.I.n3 clkbuf_1_0__f_clk.I.t53 11.0722
R26505 clkbuf_1_0__f_clk.I.n4 clkbuf_1_0__f_clk.I.t38 11.0722
R26506 clkbuf_1_0__f_clk.I.n5 clkbuf_1_0__f_clk.I.t43 11.0722
R26507 clkbuf_1_0__f_clk.I.n8 clkbuf_1_0__f_clk.I.t42 11.0722
R26508 clkbuf_1_0__f_clk.I.n7 clkbuf_1_0__f_clk.I.n6 10.5449
R26509 clkbuf_1_0__f_clk.I.n4 clkbuf_1_0__f_clk.I.n3 10.5449
R26510 clkbuf_1_0__f_clk.I.n5 clkbuf_1_0__f_clk.I.n4 10.5449
R26511 clkbuf_1_0__f_clk.I.n8 clkbuf_1_0__f_clk.I.n5 10.5449
R26512 clkbuf_1_0__f_clk.I.n8 clkbuf_1_0__f_clk.I.n7 10.5449
R26513 clkbuf_1_0__f_clk.I.n12 clkbuf_1_0__f_clk.I.n11 10.5449
R26514 clkbuf_1_0__f_clk.I.n13 clkbuf_1_0__f_clk.I.n12 10.5449
R26515 clkbuf_1_0__f_clk.I.n10 clkbuf_1_0__f_clk.I.n9 10.5449
R26516 clkbuf_1_0__f_clk.I.n14 clkbuf_1_0__f_clk.I.n10 10.5449
R26517 clkbuf_1_0__f_clk.I.n14 clkbuf_1_0__f_clk.I.n13 10.5449
R26518 clkbuf_1_0__f_clk.I.n15 clkbuf_1_0__f_clk.I 7.2005
R26519 clkbuf_1_0__f_clk.I.n40 clkbuf_1_0__f_clk.I.n39 7.0655
R26520 clkbuf_1_0__f_clk.I.n33 clkbuf_1_0__f_clk.I.n32 7.0655
R26521 clkbuf_1_0__f_clk.I.n42 clkbuf_1_0__f_clk.I.n36 6.4355
R26522 clkbuf_1_0__f_clk.I.n41 clkbuf_1_0__f_clk.I.n37 6.4355
R26523 clkbuf_1_0__f_clk.I.n40 clkbuf_1_0__f_clk.I.n38 6.4355
R26524 clkbuf_1_0__f_clk.I.n33 clkbuf_1_0__f_clk.I.n31 6.4355
R26525 clkbuf_1_0__f_clk.I.n34 clkbuf_1_0__f_clk.I.n30 6.4355
R26526 clkbuf_1_0__f_clk.I.n35 clkbuf_1_0__f_clk.I.n29 6.4355
R26527 clkbuf_1_0__f_clk.I.n16 clkbuf_1_0__f_clk.I.n15 4.5005
R26528 clkbuf_1_0__f_clk.I.n36 clkbuf_1_0__f_clk.I.t26 3.37782
R26529 clkbuf_1_0__f_clk.I.n36 clkbuf_1_0__f_clk.I.t28 3.37782
R26530 clkbuf_1_0__f_clk.I.n37 clkbuf_1_0__f_clk.I.t25 3.37782
R26531 clkbuf_1_0__f_clk.I.n37 clkbuf_1_0__f_clk.I.t24 3.37782
R26532 clkbuf_1_0__f_clk.I.n38 clkbuf_1_0__f_clk.I.t17 3.37782
R26533 clkbuf_1_0__f_clk.I.n38 clkbuf_1_0__f_clk.I.t23 3.37782
R26534 clkbuf_1_0__f_clk.I.n39 clkbuf_1_0__f_clk.I.t16 3.37782
R26535 clkbuf_1_0__f_clk.I.n39 clkbuf_1_0__f_clk.I.t19 3.37782
R26536 clkbuf_1_0__f_clk.I.n32 clkbuf_1_0__f_clk.I.t22 3.37782
R26537 clkbuf_1_0__f_clk.I.n32 clkbuf_1_0__f_clk.I.t27 3.37782
R26538 clkbuf_1_0__f_clk.I.n31 clkbuf_1_0__f_clk.I.t18 3.37782
R26539 clkbuf_1_0__f_clk.I.n31 clkbuf_1_0__f_clk.I.t20 3.37782
R26540 clkbuf_1_0__f_clk.I.n30 clkbuf_1_0__f_clk.I.t30 3.37782
R26541 clkbuf_1_0__f_clk.I.n30 clkbuf_1_0__f_clk.I.t21 3.37782
R26542 clkbuf_1_0__f_clk.I.n29 clkbuf_1_0__f_clk.I.t29 3.37782
R26543 clkbuf_1_0__f_clk.I.n29 clkbuf_1_0__f_clk.I.t31 3.37782
R26544 clkbuf_1_0__f_clk.I.n23 clkbuf_1_0__f_clk.I.n21 2.94809
R26545 clkbuf_1_0__f_clk.I.n2 clkbuf_1_0__f_clk.I.n0 2.93257
R26546 clkbuf_1_0__f_clk.I.n2 clkbuf_1_0__f_clk.I.n1 2.6005
R26547 clkbuf_1_0__f_clk.I.n18 clkbuf_1_0__f_clk.I.n17 2.6005
R26548 clkbuf_1_0__f_clk.I.n20 clkbuf_1_0__f_clk.I.n19 2.6005
R26549 clkbuf_1_0__f_clk.I.n27 clkbuf_1_0__f_clk.I.n26 2.6005
R26550 clkbuf_1_0__f_clk.I.n25 clkbuf_1_0__f_clk.I.n24 2.6005
R26551 clkbuf_1_0__f_clk.I.n23 clkbuf_1_0__f_clk.I.n22 2.6005
R26552 clkbuf_1_0__f_clk.I.n21 clkbuf_1_0__f_clk.I.t3 2.06607
R26553 clkbuf_1_0__f_clk.I.n24 clkbuf_1_0__f_clk.I.t12 2.06607
R26554 clkbuf_1_0__f_clk.I.n26 clkbuf_1_0__f_clk.I.t11 2.06607
R26555 clkbuf_1_0__f_clk.I.n19 clkbuf_1_0__f_clk.I.t6 2.06607
R26556 clkbuf_1_0__f_clk.I.n17 clkbuf_1_0__f_clk.I.t5 2.06607
R26557 clkbuf_1_0__f_clk.I.n1 clkbuf_1_0__f_clk.I.t1 2.06607
R26558 clkbuf_1_0__f_clk.I.n0 clkbuf_1_0__f_clk.I.t13 2.06607
R26559 clkbuf_1_0__f_clk.I.n22 clkbuf_1_0__f_clk.I.t2 2.06607
R26560 clkbuf_1_0__f_clk.I.n21 clkbuf_1_0__f_clk.I.t4 1.4923
R26561 clkbuf_1_0__f_clk.I.n24 clkbuf_1_0__f_clk.I.t10 1.4923
R26562 clkbuf_1_0__f_clk.I.n26 clkbuf_1_0__f_clk.I.t9 1.4923
R26563 clkbuf_1_0__f_clk.I.n19 clkbuf_1_0__f_clk.I.t8 1.4923
R26564 clkbuf_1_0__f_clk.I.n17 clkbuf_1_0__f_clk.I.t7 1.4923
R26565 clkbuf_1_0__f_clk.I.n1 clkbuf_1_0__f_clk.I.t14 1.4923
R26566 clkbuf_1_0__f_clk.I.n0 clkbuf_1_0__f_clk.I.t0 1.4923
R26567 clkbuf_1_0__f_clk.I.n22 clkbuf_1_0__f_clk.I.t15 1.4923
R26568 clkbuf_1_0__f_clk.I.n35 clkbuf_1_0__f_clk.I.n34 0.6305
R26569 clkbuf_1_0__f_clk.I.n34 clkbuf_1_0__f_clk.I.n33 0.6305
R26570 clkbuf_1_0__f_clk.I.n41 clkbuf_1_0__f_clk.I.n40 0.6305
R26571 clkbuf_1_0__f_clk.I.n42 clkbuf_1_0__f_clk.I.n41 0.6305
R26572 clkbuf_1_0__f_clk.I clkbuf_1_0__f_clk.I.n8 0.552085
R26573 clkbuf_1_0__f_clk.I clkbuf_1_0__f_clk.I.n14 0.552085
R26574 clkbuf_1_0__f_clk.I.n20 clkbuf_1_0__f_clk.I.n18 0.348086
R26575 clkbuf_1_0__f_clk.I.n27 clkbuf_1_0__f_clk.I.n25 0.348086
R26576 clkbuf_1_0__f_clk.I.n25 clkbuf_1_0__f_clk.I.n23 0.348086
R26577 clkbuf_1_0__f_clk.I.n18 clkbuf_1_0__f_clk.I.n16 0.199121
R26578 clkbuf_1_0__f_clk.I.n43 clkbuf_1_0__f_clk.I.n35 0.195969
R26579 clkbuf_1_0__f_clk.I.n43 clkbuf_1_0__f_clk.I.n42 0.181906
R26580 clkbuf_1_0__f_clk.I.n16 clkbuf_1_0__f_clk.I.n2 0.149466
R26581 clkbuf_1_0__f_clk.I.n28 clkbuf_1_0__f_clk.I.n20 0.116103
R26582 clkbuf_1_0__f_clk.I.n28 clkbuf_1_0__f_clk.I.n27 0.0928276
R26583 clkbuf_1_0__f_clk.I clkbuf_1_0__f_clk.I.n28 0.0755
R26584 clkbuf_1_0__f_clk.I clkbuf_1_0__f_clk.I.n43 0.059
R26585 _304_.ZN.n6 _304_.ZN.t11 16.5107
R26586 _304_.ZN.n9 _304_.ZN.t16 16.5107
R26587 _304_.ZN.n5 _304_.ZN.t15 16.5107
R26588 _304_.ZN.n13 _304_.ZN.t14 16.5107
R26589 _304_.ZN.n7 _304_.ZN.t17 13.5663
R26590 _304_.ZN.n8 _304_.ZN.t13 13.5663
R26591 _304_.ZN.n11 _304_.ZN.t10 13.5663
R26592 _304_.ZN.n12 _304_.ZN.t12 13.5663
R26593 _304_.ZN.n8 _304_.ZN.n7 13.3198
R26594 _304_.ZN.n12 _304_.ZN.n11 13.3198
R26595 _304_.ZN.n16 _304_.ZN.n15 11.5655
R26596 _304_.ZN.n10 _304_.ZN.n6 8.28737
R26597 _304_.ZN.n15 _304_.ZN.n5 8.02581
R26598 _304_.ZN.n14 _304_.ZN.n13 8.0005
R26599 _304_.ZN.n10 _304_.ZN.n9 8.0005
R26600 _304_.ZN.n2 _304_.ZN.n0 7.17702
R26601 _304_.ZN.n19 _304_.ZN.n17 6.72659
R26602 _304_.ZN.n2 _304_.ZN.n1 6.3005
R26603 _304_.ZN.n4 _304_.ZN.n3 6.3005
R26604 _304_.ZN.n0 _304_.ZN.t0 3.83001
R26605 _304_.ZN.n3 _304_.ZN.t1 3.83001
R26606 _304_.ZN.n19 _304_.ZN.n18 3.02702
R26607 _304_.ZN.n1 _304_.ZN.t6 1.99806
R26608 _304_.ZN.n1 _304_.ZN.t5 1.99806
R26609 _304_.ZN.n0 _304_.ZN.t9 1.70267
R26610 _304_.ZN.n3 _304_.ZN.t8 1.70267
R26611 _304_.ZN.n18 _304_.ZN.t2 1.68569
R26612 _304_.ZN.n18 _304_.ZN.t3 1.68569
R26613 _304_.ZN.n17 _304_.ZN.t4 1.6626
R26614 _304_.ZN.n17 _304_.ZN.t7 1.6626
R26615 _304_.ZN.n7 _304_.ZN.n6 1.03467
R26616 _304_.ZN.n9 _304_.ZN.n8 1.03467
R26617 _304_.ZN.n11 _304_.ZN.n5 1.03467
R26618 _304_.ZN.n13 _304_.ZN.n12 1.03467
R26619 _304_.ZN.n4 _304_.ZN.n2 0.877022
R26620 _304_.ZN.n16 _304_.ZN.n4 0.576512
R26621 _304_.ZN _304_.ZN.n10 0.492688
R26622 _304_.ZN.n14 _304_.ZN 0.368937
R26623 _304_.ZN _304_.ZN.n16 0.3155
R26624 _304_.ZN.n15 _304_.ZN.n14 0.262062
R26625 _304_.ZN _304_.ZN.n19 0.0356562
R26626 uio_oe[5] uio_oe[5].t0 4.13855
R26627 _324_.C.n30 _324_.C.n28 25.9205
R26628 _324_.C.n18 _324_.C.t28 22.7765
R26629 _324_.C.n17 _324_.C.t15 22.7765
R26630 _324_.C.n8 _324_.C.t14 22.7765
R26631 _324_.C.n7 _324_.C.t23 22.7765
R26632 _324_.C.n29 _324_.C.t10 19.7835
R26633 _324_.C.n14 _324_.C.t29 18.9805
R26634 _324_.C.n16 _324_.C.t18 18.9805
R26635 _324_.C.n27 _324_.C.t33 18.9805
R26636 _324_.C.n20 _324_.C 18.878
R26637 _324_.C.n15 _324_.C 18.6755
R26638 _324_.C.n31 _324_.C.n30 18.5405
R26639 _324_.C.n21 _324_.C.t20 18.141
R26640 _324_.C.n6 _324_.C.t26 16.3768
R26641 _324_.C.n26 _324_.C.n10 16.3355
R26642 _324_.C.n19 _324_.C.t24 16.3038
R26643 _324_.C.n12 _324_.C.t27 15.8415
R26644 _324_.C.n11 _324_.C.t31 15.8415
R26645 _324_.C.n10 _324_.C 15.4805
R26646 _324_.C.n19 _324_.C.t11 14.7222
R26647 _324_.C.n6 _324_.C.t19 14.7222
R26648 _324_.C.n29 _324_.C.t25 14.3085
R26649 _324_.C.n23 _324_.C.n20 14.2205
R26650 _324_.C.n21 _324_.C.t12 11.863
R26651 _324_.C.n14 _324_.C.t22 11.4372
R26652 _324_.C.n16 _324_.C.t32 11.4372
R26653 _324_.C.n27 _324_.C.t17 11.4372
R26654 _324_.C.n12 _324_.C.t9 11.3763
R26655 _324_.C.n11 _324_.C.t13 11.3763
R26656 _324_.C.n26 _324_.C.n25 10.2605
R26657 _324_.C.n28 _324_.C 9.67858
R26658 _324_.C.n30 _324_.C 9.67313
R26659 _324_.C.n13 _324_.C.n11 9.1255
R26660 _324_.C.n18 _324_.C.t16 8.73617
R26661 _324_.C.n17 _324_.C.t21 8.73617
R26662 _324_.C.n8 _324_.C.t30 8.73617
R26663 _324_.C.n7 _324_.C.t8 8.73617
R26664 _324_.C _324_.C.n17 8.27191
R26665 _324_.C _324_.C.n19 8.24092
R26666 _324_.C _324_.C.n6 8.21104
R26667 _324_.C _324_.C.n27 8.11576
R26668 _324_.C _324_.C.n14 8.11457
R26669 _324_.C _324_.C.n16 8.11457
R26670 _324_.C.n9 _324_.C.n7 8.11441
R26671 _324_.C _324_.C.n18 8.03566
R26672 _324_.C _324_.C.n8 8.03566
R26673 _324_.C _324_.C.n29 8.00997
R26674 _324_.C.n22 _324_.C.n21 8.0005
R26675 _324_.C.n28 _324_.C.n26 7.9205
R26676 _324_.C.n2 _324_.C.n1 7.33746
R26677 _324_.C.n25 _324_.C.n15 7.2005
R26678 _324_.C.n2 _324_.C.n0 6.46093
R26679 _324_.C.n15 _324_.C 6.2555
R26680 _324_.C.n24 _324_.C.n23 6.0755
R26681 _324_.C.n31 _324_.C.n5 5.49618
R26682 _324_.C.n4 _324_.C.n3 5.4118
R26683 _324_.C.n24 _324_.C 4.77358
R26684 _324_.C.n23 _324_.C.n22 4.67072
R26685 _324_.C.n20 _324_.C 4.5005
R26686 _324_.C.n25 _324_.C.n24 4.5005
R26687 _324_.C.n10 _324_.C.n9 4.5005
R26688 _324_.C.n0 _324_.C.t5 3.6005
R26689 _324_.C.n0 _324_.C.t6 3.6005
R26690 _324_.C.n1 _324_.C.t4 3.6005
R26691 _324_.C.n1 _324_.C.t7 3.6005
R26692 _324_.C _324_.C.n13 2.69288
R26693 _324_.C.n5 _324_.C.t0 2.06607
R26694 _324_.C.n3 _324_.C.t2 2.06607
R26695 _324_.C.n5 _324_.C.t1 1.4923
R26696 _324_.C.n3 _324_.C.t3 1.4923
R26697 _324_.C.n13 _324_.C.n12 1.41994
R26698 _324_.C.n4 _324_.C.n2 0.439189
R26699 _324_.C _324_.C.n31 0.3155
R26700 _324_.C _324_.C.n4 0.203
R26701 _324_.C.n9 _324_.C 0.158
R26702 _324_.C.n22 _324_.C 0.0878134
R26703 _359_.B _359_.B.n11 24.1205
R26704 _359_.B.n10 _359_.B.t8 18.6885
R26705 _359_.B.n7 _359_.B.t4 17.8003
R26706 _359_.B.n2 _359_.B.t5 17.6422
R26707 _359_.B.n0 _359_.B.t9 17.119
R26708 _359_.B.n9 _359_.B.n8 15.5894
R26709 _359_.B.n5 _359_.B.t3 15.3305
R26710 _359_.B.n5 _359_.B.t10 15.0872
R26711 _359_.B.n2 _359_.B.t11 14.8925
R26712 _359_.B.n7 _359_.B.t6 14.7465
R26713 _359_.B.n0 _359_.B.t2 12.7147
R26714 _359_.B.n10 _359_.B.t7 11.9603
R26715 _359_.B.n4 _359_.B.n1 11.3562
R26716 _359_.B.n11 _359_.B 11.1457
R26717 _359_.B.n4 _359_.B.n3 10.5637
R26718 _359_.B.n6 _359_.B 9.86874
R26719 _359_.B _359_.B.t1 8.69622
R26720 _359_.B _359_.B.n5 8.15932
R26721 _359_.B.n1 _359_.B.n0 8.0005
R26722 _359_.B.n3 _359_.B.n2 8.0005
R26723 _359_.B.n8 _359_.B.n7 8.0005
R26724 _359_.B _359_.B.t0 6.72245
R26725 _359_.B.n6 _359_.B.n4 5.5805
R26726 _359_.B _359_.B.n10 4.08607
R26727 _359_.B.n11 _359_.B.n9 3.0605
R26728 _359_.B.n9 _359_.B.n6 2.7005
R26729 _359_.B.n8 _359_.B 0.114184
R26730 _359_.B.n1 _359_.B 0.0820131
R26731 _359_.B.n3 _359_.B 0.00997368
R26732 a_26916_25640.n3 a_26916_25640.t3 121.874
R26733 a_26916_25640.t3 a_26916_25640.t4 61.5152
R26734 a_26916_25640.n0 a_26916_25640.t6 52.378
R26735 a_26916_25640.n0 a_26916_25640.t2 17.7882
R26736 a_26916_25640.n2 a_26916_25640.t1 11.1158
R26737 a_26916_25640.n4 a_26916_25640.n3 9.95623
R26738 a_26916_25640.t0 a_26916_25640.n4 8.02846
R26739 a_26916_25640.n2 a_26916_25640.n1 8.0005
R26740 a_26916_25640.n3 a_26916_25640.t5 6.7165
R26741 a_26916_25640.n1 a_26916_25640.t7 5.96217
R26742 a_26916_25640.n1 a_26916_25640.n0 1.33883
R26743 a_26916_25640.n4 a_26916_25640.n2 0.376152
R26744 _287_.A1.n46 _287_.A1.n45 18.9805
R26745 _287_.A1.n41 _287_.A1.n40 18.9805
R26746 _287_.A1.n22 _287_.A1.n21 18.9805
R26747 _287_.A1.n17 _287_.A1.n16 18.9805
R26748 _287_.A1.n34 _287_.A1.n33 18.9805
R26749 _287_.A1.n28 _287_.A1.n27 18.9805
R26750 _287_.A1.n11 _287_.A1.n10 18.9805
R26751 _287_.A1.n6 _287_.A1.n5 18.9805
R26752 _287_.A1.n21 _287_.A1.t11 15.2088
R26753 _287_.A1.n22 _287_.A1.t15 15.2088
R26754 _287_.A1.n16 _287_.A1.t23 15.2088
R26755 _287_.A1.n17 _287_.A1.t20 15.2088
R26756 _287_.A1.n11 _287_.A1.t24 15.2088
R26757 _287_.A1.n10 _287_.A1.t28 15.2088
R26758 _287_.A1.n5 _287_.A1.t8 15.2088
R26759 _287_.A1.n6 _287_.A1.t33 15.2088
R26760 _287_.A1.n46 _287_.A1.t34 15.148
R26761 _287_.A1.n45 _287_.A1.t31 15.148
R26762 _287_.A1.n40 _287_.A1.t12 15.148
R26763 _287_.A1.n41 _287_.A1.t9 15.148
R26764 _287_.A1.n33 _287_.A1.t22 15.148
R26765 _287_.A1.n34 _287_.A1.t29 15.148
R26766 _287_.A1.n27 _287_.A1.t39 15.148
R26767 _287_.A1.n28 _287_.A1.t37 15.148
R26768 _287_.A1.n47 _287_.A1.t27 14.7222
R26769 _287_.A1.n44 _287_.A1.t36 14.7222
R26770 _287_.A1.n39 _287_.A1.t32 14.7222
R26771 _287_.A1.n42 _287_.A1.t16 14.7222
R26772 _287_.A1.n20 _287_.A1.t18 14.7222
R26773 _287_.A1.n23 _287_.A1.t17 14.7222
R26774 _287_.A1.n15 _287_.A1.t25 14.7222
R26775 _287_.A1.n18 _287_.A1.t26 14.7222
R26776 _287_.A1.n32 _287_.A1.t14 14.7222
R26777 _287_.A1.n35 _287_.A1.t35 14.7222
R26778 _287_.A1.n26 _287_.A1.t30 14.7222
R26779 _287_.A1.n29 _287_.A1.t13 14.7222
R26780 _287_.A1.n12 _287_.A1.t21 14.7222
R26781 _287_.A1.n9 _287_.A1.t10 14.7222
R26782 _287_.A1.n4 _287_.A1.t38 14.7222
R26783 _287_.A1.n7 _287_.A1.t19 14.7222
R26784 _287_.A1.n38 _287_.A1.n14 14.0405
R26785 _287_.A1.n51 _287_.A1.n50 11.3405
R26786 _287_.A1.n50 _287_.A1.n49 9.0005
R26787 _287_.A1.n48 _287_.A1.n44 8.34081
R26788 _287_.A1.n19 _287_.A1.n15 8.34081
R26789 _287_.A1.n13 _287_.A1.n9 8.34081
R26790 _287_.A1.n43 _287_.A1.n39 8.33378
R26791 _287_.A1.n24 _287_.A1.n20 8.33378
R26792 _287_.A1.n30 _287_.A1.n26 8.33378
R26793 _287_.A1.n8 _287_.A1.n4 8.33378
R26794 _287_.A1.n43 _287_.A1.n42 8.0005
R26795 _287_.A1.n48 _287_.A1.n47 8.0005
R26796 _287_.A1.n19 _287_.A1.n18 8.0005
R26797 _287_.A1.n24 _287_.A1.n23 8.0005
R26798 _287_.A1.n30 _287_.A1.n29 8.0005
R26799 _287_.A1.n36 _287_.A1.n35 8.0005
R26800 _287_.A1.n32 _287_.A1.n31 8.0005
R26801 _287_.A1.n8 _287_.A1.n7 8.0005
R26802 _287_.A1.n13 _287_.A1.n12 8.0005
R26803 _287_.A1.n3 _287_.A1.n2 7.33746
R26804 _287_.A1.n3 _287_.A1.n1 6.46093
R26805 _287_.A1 _287_.A1.n0 5.81118
R26806 _287_.A1.n37 _287_.A1.n25 5.7605
R26807 _287_.A1.n53 _287_.A1.n52 5.4118
R26808 _287_.A1.n50 _287_.A1.n38 5.3105
R26809 _287_.A1.n38 _287_.A1.n37 4.6805
R26810 _287_.A1.n37 _287_.A1.n36 4.61862
R26811 _287_.A1.n2 _287_.A1.t4 3.6005
R26812 _287_.A1.n2 _287_.A1.t5 3.6005
R26813 _287_.A1.n1 _287_.A1.t6 3.6005
R26814 _287_.A1.n1 _287_.A1.t7 3.6005
R26815 _287_.A1.n0 _287_.A1.t1 2.06607
R26816 _287_.A1.n52 _287_.A1.t3 2.06607
R26817 _287_.A1.n0 _287_.A1.t2 1.4923
R26818 _287_.A1.n52 _287_.A1.t0 1.4923
R26819 _287_.A1.n47 _287_.A1.n46 1.0955
R26820 _287_.A1.n45 _287_.A1.n44 1.0955
R26821 _287_.A1.n40 _287_.A1.n39 1.0955
R26822 _287_.A1.n42 _287_.A1.n41 1.0955
R26823 _287_.A1.n21 _287_.A1.n20 1.0955
R26824 _287_.A1.n23 _287_.A1.n22 1.0955
R26825 _287_.A1.n16 _287_.A1.n15 1.0955
R26826 _287_.A1.n18 _287_.A1.n17 1.0955
R26827 _287_.A1.n33 _287_.A1.n32 1.0955
R26828 _287_.A1.n35 _287_.A1.n34 1.0955
R26829 _287_.A1.n27 _287_.A1.n26 1.0955
R26830 _287_.A1.n29 _287_.A1.n28 1.0955
R26831 _287_.A1.n12 _287_.A1.n11 1.0955
R26832 _287_.A1.n10 _287_.A1.n9 1.0955
R26833 _287_.A1.n5 _287_.A1.n4 1.0955
R26834 _287_.A1.n7 _287_.A1.n6 1.0955
R26835 _287_.A1.n31 _287_.A1 0.487062
R26836 _287_.A1 _287_.A1.n13 0.487062
R26837 _287_.A1 _287_.A1.n43 0.43925
R26838 _287_.A1 _287_.A1.n24 0.43925
R26839 _287_.A1 _287_.A1.n30 0.43925
R26840 _287_.A1.n36 _287_.A1.n31 0.340813
R26841 _287_.A1.n49 _287_.A1.n48 0.329562
R26842 _287_.A1.n25 _287_.A1.n19 0.329562
R26843 _287_.A1.n14 _287_.A1.n8 0.28175
R26844 _287_.A1.n53 _287_.A1.n51 0.2255
R26845 _287_.A1.n51 _287_.A1.n3 0.214189
R26846 _287_.A1 _287_.A1.n53 0.203
R26847 _287_.A1.n49 _287_.A1 0.158
R26848 _287_.A1.n25 _287_.A1 0.158
R26849 _287_.A1.n14 _287_.A1 0.158
R26850 uo_out[6].n8 uo_out[6] 23.3626
R26851 uo_out[6].n5 uo_out[6].n4 7.21811
R26852 uo_out[6].n5 uo_out[6].n3 6.36507
R26853 uo_out[6].n6 uo_out[6].n2 6.36507
R26854 uo_out[6].n7 uo_out[6].n1 6.36507
R26855 uo_out[6] uo_out[6].n10 3.81667
R26856 uo_out[6].n4 uo_out[6].t9 2.89962
R26857 uo_out[6].n4 uo_out[6].t2 2.89962
R26858 uo_out[6].n3 uo_out[6].t1 2.89962
R26859 uo_out[6].n3 uo_out[6].t10 2.89962
R26860 uo_out[6].n2 uo_out[6].t8 2.89962
R26861 uo_out[6].n2 uo_out[6].t3 2.89962
R26862 uo_out[6].n1 uo_out[6].t0 2.89962
R26863 uo_out[6].n1 uo_out[6].t11 2.89962
R26864 uo_out[6].n9 uo_out[6].n0 2.70811
R26865 uo_out[6].n10 uo_out[6].t6 2.06607
R26866 uo_out[6].n10 uo_out[6].t4 2.06607
R26867 uo_out[6].n0 uo_out[6].t7 2.06607
R26868 uo_out[6].n0 uo_out[6].t5 2.06607
R26869 uo_out[6].n8 uo_out[6].n7 1.34342
R26870 uo_out[6].n7 uo_out[6].n6 0.877022
R26871 uo_out[6].n6 uo_out[6].n5 0.877022
R26872 uo_out[6] uo_out[6].n9 0.267929
R26873 uo_out[6].n9 uo_out[6].n8 0.165071
R26874 _268_.A1.n8 _268_.A1.t2 19.2725
R26875 _268_.A1.n0 _268_.A1.t7 18.6885
R26876 _268_.A1.n2 _268_.A1.t4 16.0118
R26877 _268_.A1.n4 _268_.A1.t3 15.3305
R26878 _268_.A1.n4 _268_.A1.t8 15.148
R26879 _268_.A1.n6 _268_.A1.n5 14.7605
R26880 _268_.A1.n8 _268_.A1.t6 13.8948
R26881 _268_.A1.n2 _268_.A1.t5 13.2622
R26882 _268_.A1.n10 _268_.A1.n9 12.9236
R26883 _268_.A1.n0 _268_.A1.t9 11.8873
R26884 _268_.A1.n10 _268_.A1.t1 9.713
R26885 _268_.A1.n9 _268_.A1 9.0005
R26886 _268_.A1 _268_.A1.n8 8.11085
R26887 _268_.A1.n5 _268_.A1.n4 8.01109
R26888 _268_.A1.n3 _268_.A1.n2 8.0005
R26889 _268_.A1.n9 _268_.A1.n7 6.6605
R26890 _268_.A1.n7 _268_.A1.n1 4.98927
R26891 _268_.A1.n6 _268_.A1.n3 4.71591
R26892 _268_.A1 _268_.A1.t0 4.35156
R26893 _268_.A1.n1 _268_.A1.n0 4.0005
R26894 _268_.A1.n7 _268_.A1.n6 1.0355
R26895 _268_.A1 _268_.A1.n10 0.293336
R26896 _268_.A1.n5 _268_.A1 0.148735
R26897 _268_.A1.n3 _268_.A1 0.130336
R26898 _268_.A1.n1 _268_.A1 0.0860738
R26899 _474_.CLK.n34 _474_.CLK.t32 28.5265
R26900 _474_.CLK.n26 _474_.CLK.t54 18.6885
R26901 _474_.CLK.n39 _474_.CLK.t51 18.6885
R26902 _474_.CLK.n33 _474_.CLK.t44 18.6885
R26903 _474_.CLK.n19 _474_.CLK 18.0005
R26904 _474_.CLK.n28 _474_.CLK.t38 17.5205
R26905 _474_.CLK.n35 _474_.CLK 17.2805
R26906 _474_.CLK.n22 _474_.CLK.n19 15.5255
R26907 _474_.CLK.n30 _474_.CLK.n27 13.9461
R26908 _474_.CLK.n43 _474_.CLK.t50 13.907
R26909 _474_.CLK.n32 _474_.CLK.t34 13.907
R26910 _474_.CLK.n23 _474_.CLK.t43 13.907
R26911 _474_.CLK.n16 _474_.CLK.t39 13.907
R26912 _474_.CLK.n31 _474_.CLK.t49 13.8462
R26913 _474_.CLK.n37 _474_.CLK.t42 13.8462
R26914 _474_.CLK.n18 _474_.CLK.t35 13.8462
R26915 _474_.CLK.n20 _474_.CLK.t37 13.8462
R26916 _474_.CLK.n33 _474_.CLK.t56 12.1672
R26917 _474_.CLK.n31 _474_.CLK.t48 12.1185
R26918 _474_.CLK.n37 _474_.CLK.t41 12.1185
R26919 _474_.CLK.n18 _474_.CLK.t47 12.1185
R26920 _474_.CLK.n20 _474_.CLK.t33 12.1185
R26921 _474_.CLK.n43 _474_.CLK.t46 12.0455
R26922 _474_.CLK.n32 _474_.CLK.t55 12.0455
R26923 _474_.CLK.n23 _474_.CLK.t36 12.0455
R26924 _474_.CLK.n16 _474_.CLK.t53 12.0455
R26925 _474_.CLK.n26 _474_.CLK.t40 11.9603
R26926 _474_.CLK.n39 _474_.CLK.t52 11.8873
R26927 _474_.CLK.n28 _474_.CLK.t45 11.5588
R26928 _474_.CLK.n47 _474_.CLK.n46 10.8005
R26929 _474_.CLK.n36 _474_.CLK 10.4405
R26930 _474_.CLK.n46 _474_.CLK.n25 10.2605
R26931 _474_.CLK.n30 _474_.CLK.n29 9.46296
R26932 _474_.CLK.n36 _474_.CLK.n35 9.4505
R26933 _474_.CLK.n38 _474_.CLK 9.1805
R26934 _474_.CLK.n41 _474_.CLK.n40 9.0005
R26935 _474_.CLK _474_.CLK.n31 8.01471
R26936 _474_.CLK _474_.CLK.n37 8.01471
R26937 _474_.CLK _474_.CLK.n32 8.01471
R26938 _474_.CLK _474_.CLK.n18 8.01471
R26939 _474_.CLK.n44 _474_.CLK.n43 8.0005
R26940 _474_.CLK.n29 _474_.CLK.n28 8.0005
R26941 _474_.CLK.n24 _474_.CLK.n23 8.0005
R26942 _474_.CLK.n17 _474_.CLK.n16 8.0005
R26943 _474_.CLK.n21 _474_.CLK.n20 8.0005
R26944 _474_.CLK.n11 _474_.CLK.n10 7.0655
R26945 _474_.CLK.n4 _474_.CLK.n3 7.0655
R26946 _474_.CLK.n42 _474_.CLK.n41 6.8405
R26947 _474_.CLK.n45 _474_.CLK.n42 6.7505
R26948 _474_.CLK.n22 _474_.CLK.n21 6.55392
R26949 _474_.CLK.n11 _474_.CLK.n9 6.4355
R26950 _474_.CLK.n12 _474_.CLK.n8 6.4355
R26951 _474_.CLK.n13 _474_.CLK.n7 6.4355
R26952 _474_.CLK.n6 _474_.CLK.n0 6.4355
R26953 _474_.CLK.n5 _474_.CLK.n1 6.4355
R26954 _474_.CLK.n4 _474_.CLK.n2 6.4355
R26955 _474_.CLK.n46 _474_.CLK.n45 5.9405
R26956 _474_.CLK.n42 _474_.CLK.n30 5.5805
R26957 _474_.CLK.n38 _474_.CLK.n36 4.6805
R26958 _474_.CLK.n45 _474_.CLK.n44 4.61892
R26959 _474_.CLK.n25 _474_.CLK.n24 4.61892
R26960 _474_.CLK.n19 _474_.CLK.n17 4.61892
R26961 _474_.CLK.n35 _474_.CLK 4.5005
R26962 _474_.CLK.n40 _474_.CLK.n39 4.08017
R26963 _474_.CLK.n27 _474_.CLK.n26 4.0005
R26964 _474_.CLK.n10 _474_.CLK.t17 3.37782
R26965 _474_.CLK.n10 _474_.CLK.t22 3.37782
R26966 _474_.CLK.n9 _474_.CLK.t21 3.37782
R26967 _474_.CLK.n9 _474_.CLK.t12 3.37782
R26968 _474_.CLK.n8 _474_.CLK.t8 3.37782
R26969 _474_.CLK.n8 _474_.CLK.t2 3.37782
R26970 _474_.CLK.n7 _474_.CLK.t7 3.37782
R26971 _474_.CLK.n7 _474_.CLK.t27 3.37782
R26972 _474_.CLK.n0 _474_.CLK.t30 3.37782
R26973 _474_.CLK.n0 _474_.CLK.t25 3.37782
R26974 _474_.CLK.n1 _474_.CLK.t23 3.37782
R26975 _474_.CLK.n1 _474_.CLK.t19 3.37782
R26976 _474_.CLK.n2 _474_.CLK.t14 3.37782
R26977 _474_.CLK.n2 _474_.CLK.t18 3.37782
R26978 _474_.CLK.n3 _474_.CLK.t13 3.37782
R26979 _474_.CLK.n3 _474_.CLK.t10 3.37782
R26980 _474_.CLK.n56 _474_.CLK.n54 2.93257
R26981 _474_.CLK _474_.CLK.n34 2.6957
R26982 _474_.CLK.n47 _474_.CLK.n15 2.62533
R26983 _474_.CLK.n49 _474_.CLK.n48 2.6005
R26984 _474_.CLK.n51 _474_.CLK.n50 2.6005
R26985 _474_.CLK.n53 _474_.CLK.n52 2.6005
R26986 _474_.CLK.n60 _474_.CLK.n59 2.6005
R26987 _474_.CLK.n58 _474_.CLK.n57 2.6005
R26988 _474_.CLK.n56 _474_.CLK.n55 2.6005
R26989 _474_.CLK.n41 _474_.CLK.n38 2.2505
R26990 _474_.CLK.n55 _474_.CLK.t1 2.06607
R26991 _474_.CLK.n57 _474_.CLK.t11 2.06607
R26992 _474_.CLK.n59 _474_.CLK.t20 2.06607
R26993 _474_.CLK.n52 _474_.CLK.t26 2.06607
R26994 _474_.CLK.n50 _474_.CLK.t28 2.06607
R26995 _474_.CLK.n48 _474_.CLK.t6 2.06607
R26996 _474_.CLK.n15 _474_.CLK.t3 2.06607
R26997 _474_.CLK.n54 _474_.CLK.t29 2.06607
R26998 _474_.CLK.n55 _474_.CLK.t4 1.4923
R26999 _474_.CLK.n57 _474_.CLK.t5 1.4923
R27000 _474_.CLK.n59 _474_.CLK.t15 1.4923
R27001 _474_.CLK.n52 _474_.CLK.t16 1.4923
R27002 _474_.CLK.n50 _474_.CLK.t24 1.4923
R27003 _474_.CLK.n48 _474_.CLK.t31 1.4923
R27004 _474_.CLK.n15 _474_.CLK.t9 1.4923
R27005 _474_.CLK.n54 _474_.CLK.t0 1.4923
R27006 _474_.CLK.n25 _474_.CLK.n22 1.0355
R27007 _474_.CLK.n34 _474_.CLK.n33 1.0005
R27008 _474_.CLK.n6 _474_.CLK.n5 0.6305
R27009 _474_.CLK.n5 _474_.CLK.n4 0.6305
R27010 _474_.CLK.n12 _474_.CLK.n11 0.6305
R27011 _474_.CLK.n13 _474_.CLK.n12 0.6305
R27012 _474_.CLK.n51 _474_.CLK.n49 0.348086
R27013 _474_.CLK.n53 _474_.CLK.n51 0.348086
R27014 _474_.CLK.n60 _474_.CLK.n58 0.348086
R27015 _474_.CLK.n58 _474_.CLK.n56 0.348086
R27016 _474_.CLK.n49 _474_.CLK.n47 0.323259
R27017 _474_.CLK.n27 _474_.CLK 0.245418
R27018 _474_.CLK.n14 _474_.CLK.n13 0.195969
R27019 _474_.CLK.n14 _474_.CLK.n6 0.181906
R27020 _474_.CLK.n40 _474_.CLK 0.165746
R27021 _474_.CLK.n61 _474_.CLK.n60 0.116103
R27022 _474_.CLK.n61 _474_.CLK.n53 0.0928276
R27023 _474_.CLK _474_.CLK.n61 0.0755
R27024 _474_.CLK _474_.CLK.n14 0.059
R27025 _474_.CLK.n29 _474_.CLK 0.0531154
R27026 _474_.CLK.n44 _474_.CLK 0.0147105
R27027 _474_.CLK.n24 _474_.CLK 0.0147105
R27028 _474_.CLK.n17 _474_.CLK 0.0147105
R27029 _474_.CLK.n21 _474_.CLK 0.0147105
R27030 _402_.A1.n22 _402_.A1 24.1205
R27031 _402_.A1.n2 _402_.A1.t17 22.1195
R27032 _402_.A1.n7 _402_.A1.t12 20.1161
R27033 _402_.A1.n3 _402_.A1.t7 19.5645
R27034 _402_.A1.n4 _402_.A1.t20 19.5645
R27035 _402_.A1.n12 _402_.A1.t15 18.9805
R27036 _402_.A1.n3 _402_.A1.t5 18.4938
R27037 _402_.A1.n7 _402_.A1.t18 18.2505
R27038 _402_.A1.n14 _402_.A1.t16 17.7395
R27039 _402_.A1.n6 _402_.A1.t14 17.5205
R27040 _402_.A1.n19 _402_.A1.t22 17.484
R27041 _402_.A1.n8 _402_.A1.t9 17.3623
R27042 _402_.A1.n4 _402_.A1.t4 17.1312
R27043 _402_.A1.n17 _402_.A1.t21 16.3282
R27044 _402_.A1.n17 _402_.A1.t19 14.7465
R27045 _402_.A1.n8 _402_.A1.t8 14.6735
R27046 _402_.A1.n13 _402_.A1.n11 14.0405
R27047 _402_.A1.n14 _402_.A1.t11 12.6782
R27048 _402_.A1.n19 _402_.A1.t6 11.863
R27049 _402_.A1.n11 _402_.A1.n5 11.7005
R27050 _402_.A1.n6 _402_.A1.t13 11.5588
R27051 _402_.A1.n12 _402_.A1.t10 11.4372
R27052 _402_.A1.n16 _402_.A1.n15 9.78214
R27053 _402_.A1.n13 _402_.A1 9.7205
R27054 _402_.A1.n2 _402_.A1.t23 9.02817
R27055 _402_.A1.n22 _402_.A1.n21 8.8205
R27056 _402_.A1 _402_.A1.n3 8.51318
R27057 _402_.A1.n21 _402_.A1.n20 8.4605
R27058 _402_.A1 _402_.A1.n2 8.35407
R27059 _402_.A1 _402_.A1.n12 8.11457
R27060 _402_.A1.n9 _402_.A1.n7 8.10471
R27061 _402_.A1 _402_.A1.n19 8.08781
R27062 _402_.A1 _402_.A1.n6 8.05312
R27063 _402_.A1 _402_.A1.n8 8.02171
R27064 _402_.A1.n18 _402_.A1.n17 8.00405
R27065 _402_.A1.n5 _402_.A1.n4 8.0005
R27066 _402_.A1.n20 _402_.A1.n18 7.9655
R27067 _402_.A1.n10 _402_.A1 7.6505
R27068 _402_.A1 _402_.A1.n1 6.75428
R27069 _402_.A1 _402_.A1.n0 5.26469
R27070 _402_.A1 _402_.A1.n22 4.8605
R27071 _402_.A1.n20 _402_.A1 4.65095
R27072 _402_.A1.n10 _402_.A1.n9 4.5005
R27073 _402_.A1.n11 _402_.A1.n10 4.5005
R27074 _402_.A1.n15 _402_.A1.n14 4.0005
R27075 _402_.A1.n1 _402_.A1.t3 1.99806
R27076 _402_.A1.n1 _402_.A1.t2 1.99806
R27077 _402_.A1.n9 _402_.A1 1.68584
R27078 _402_.A1.n0 _402_.A1.t0 1.4923
R27079 _402_.A1.n0 _402_.A1.t1 1.4923
R27080 _402_.A1.n21 _402_.A1.n16 0.9005
R27081 _402_.A1.n16 _402_.A1.n13 0.3605
R27082 _402_.A1.n5 _402_.A1 0.1405
R27083 _402_.A1.n18 _402_.A1 0.133132
R27084 _402_.A1.n15 _402_.A1 0.0769384
R27085 _324_.B.n3 _324_.B.t25 23.5065
R27086 _324_.B.n13 _324_.B 18.8208
R27087 _324_.B.n2 _324_.B.t32 18.6885
R27088 _324_.B.n1 _324_.B.t20 17.5205
R27089 _324_.B.n4 _324_.B.n3 16.5048
R27090 _324_.B.n11 _324_.B.t29 16.4012
R27091 _324_.B.n10 _324_.B.t31 16.3282
R27092 _324_.B.n9 _324_.B.t22 16.3038
R27093 _324_.B.n10 _324_.B.t33 15.1845
R27094 _324_.B.n11 _324_.B.t24 15.1115
R27095 _324_.B.n9 _324_.B.t23 14.7222
R27096 _324_.B.n5 _324_.B.t27 14.6735
R27097 _324_.B.n2 _324_.B.t21 11.9603
R27098 _324_.B.n1 _324_.B.t26 11.5588
R27099 _324_.B.n7 _324_.B 11.1605
R27100 _324_.B.n7 _324_.B.n6 10.7832
R27101 _324_.B.n3 _324_.B.t28 9.69733
R27102 _324_.B.n8 _324_.B 9.27873
R27103 _324_.B.n4 _324_.B.t30 8.88217
R27104 _324_.B.n5 _324_.B.n4 8.55367
R27105 _324_.B _324_.B.n10 8.37737
R27106 _324_.B.n12 _324_.B.n11 8.15519
R27107 _324_.B _324_.B.n1 8.05312
R27108 _324_.B _324_.B.n9 8.02581
R27109 _324_.B.n6 _324_.B.n5 8.0005
R27110 _324_.B.n14 _324_.B.n8 7.5605
R27111 _324_.B.n27 _324_.B.n25 7.17702
R27112 _324_.B.n29 _324_.B.n28 6.3005
R27113 _324_.B.n31 _324_.B.n30 6.3005
R27114 _324_.B.n27 _324_.B.n26 6.3005
R27115 _324_.B.n20 _324_.B.n18 5.73397
R27116 _324_.B.n17 _324_.B.n16 5.2005
R27117 _324_.B.n20 _324_.B.n19 5.2005
R27118 _324_.B.n22 _324_.B.n21 5.2005
R27119 _324_.B.n24 _324_.B.n23 5.2005
R27120 _324_.B.n13 _324_.B.n12 4.5005
R27121 _324_.B.n15 _324_.B.n14 4.5005
R27122 _324_.B _324_.B.n2 4.08607
R27123 _324_.B.n30 _324_.B.t2 3.83001
R27124 _324_.B.n25 _324_.B.t1 3.83001
R27125 _324_.B.n15 _324_.B.n0 2.64381
R27126 _324_.B.n28 _324_.B.t0 1.99806
R27127 _324_.B.n28 _324_.B.t8 1.99806
R27128 _324_.B.n26 _324_.B.t7 1.99806
R27129 _324_.B.n26 _324_.B.t3 1.99806
R27130 _324_.B.n8 _324_.B.n7 1.9805
R27131 _324_.B.n23 _324_.B.t15 1.84822
R27132 _324_.B.n23 _324_.B.t17 1.84822
R27133 _324_.B.n21 _324_.B.t18 1.84822
R27134 _324_.B.n21 _324_.B.t13 1.84822
R27135 _324_.B.n19 _324_.B.t14 1.84822
R27136 _324_.B.n19 _324_.B.t16 1.84822
R27137 _324_.B.n18 _324_.B.t19 1.84822
R27138 _324_.B.n18 _324_.B.t12 1.84822
R27139 _324_.B.n30 _324_.B.t9 1.70267
R27140 _324_.B.n25 _324_.B.t6 1.70267
R27141 _324_.B.n16 _324_.B.t10 1.6626
R27142 _324_.B.n16 _324_.B.t11 1.6626
R27143 _324_.B.n0 _324_.B.t4 1.6626
R27144 _324_.B.n0 _324_.B.t5 1.6626
R27145 _324_.B.n17 _324_.B.n15 1.23977
R27146 _324_.B.n32 _324_.B.n31 0.985548
R27147 _324_.B.n14 _324_.B.n13 0.9005
R27148 _324_.B.n29 _324_.B.n27 0.877022
R27149 _324_.B.n31 _324_.B.n29 0.877022
R27150 _324_.B.n22 _324_.B.n20 0.533966
R27151 _324_.B.n24 _324_.B.n22 0.533966
R27152 _324_.B _324_.B.n17 0.388625
R27153 _324_.B.n12 _324_.B 0.3155
R27154 _324_.B _324_.B.n32 0.283766
R27155 _324_.B.n32 _324_.B.n24 0.227215
R27156 _324_.B.n6 _324_.B 0.127885
R27157 uo_out[2].n10 uo_out[2] 16.7026
R27158 uo_out[2].n5 uo_out[2].n4 7.21811
R27159 uo_out[2].n7 uo_out[2].n1 6.36507
R27160 uo_out[2].n6 uo_out[2].n2 6.36507
R27161 uo_out[2].n5 uo_out[2].n3 6.36507
R27162 uo_out[2].n10 uo_out[2].n9 3.01668
R27163 uo_out[2].n1 uo_out[2].t9 2.89962
R27164 uo_out[2].n1 uo_out[2].t6 2.89962
R27165 uo_out[2].n2 uo_out[2].t7 2.89962
R27166 uo_out[2].n2 uo_out[2].t11 2.89962
R27167 uo_out[2].n3 uo_out[2].t10 2.89962
R27168 uo_out[2].n3 uo_out[2].t4 2.89962
R27169 uo_out[2].n4 uo_out[2].t5 2.89962
R27170 uo_out[2].n4 uo_out[2].t8 2.89962
R27171 uo_out[2].n8 uo_out[2].n0 2.70811
R27172 uo_out[2].n0 uo_out[2].t2 2.06607
R27173 uo_out[2].n0 uo_out[2].t3 2.06607
R27174 uo_out[2].n9 uo_out[2].t0 2.06607
R27175 uo_out[2].n9 uo_out[2].t1 2.06607
R27176 uo_out[2].n8 uo_out[2].n7 1.50949
R27177 uo_out[2].n7 uo_out[2].n6 0.877022
R27178 uo_out[2].n6 uo_out[2].n5 0.877022
R27179 uo_out[2] uo_out[2].n10 0.800488
R27180 uo_out[2] uo_out[2].n8 0.267929
R27181 vgaringosc.workerclkbuff_notouch_.I.n4 vgaringosc.workerclkbuff_notouch_.I.t9 31.6987
R27182 vgaringosc.workerclkbuff_notouch_.I.n4 vgaringosc.workerclkbuff_notouch_.I.t7 18.6885
R27183 vgaringosc.workerclkbuff_notouch_.I.n2 vgaringosc.workerclkbuff_notouch_.I.t8 18.6885
R27184 vgaringosc.workerclkbuff_notouch_.I.n3 vgaringosc.workerclkbuff_notouch_.I.t4 18.6885
R27185 vgaringosc.workerclkbuff_notouch_.I.n4 vgaringosc.workerclkbuff_notouch_.I.t10 11.133
R27186 vgaringosc.workerclkbuff_notouch_.I.n2 vgaringosc.workerclkbuff_notouch_.I.t6 11.133
R27187 vgaringosc.workerclkbuff_notouch_.I.n3 vgaringosc.workerclkbuff_notouch_.I.t5 11.133
R27188 vgaringosc.workerclkbuff_notouch_.I.n3 vgaringosc.workerclkbuff_notouch_.I.n2 10.5449
R27189 vgaringosc.workerclkbuff_notouch_.I vgaringosc.workerclkbuff_notouch_.I.n0 6.62914
R27190 vgaringosc.workerclkbuff_notouch_.I.n5 vgaringosc.workerclkbuff_notouch_.I.n4 6.48939
R27191 vgaringosc.workerclkbuff_notouch_.I vgaringosc.workerclkbuff_notouch_.I.n1 5.57959
R27192 vgaringosc.workerclkbuff_notouch_.I.n5 vgaringosc.workerclkbuff_notouch_.I.n3 4.05606
R27193 vgaringosc.workerclkbuff_notouch_.I.n0 vgaringosc.workerclkbuff_notouch_.I.t0 2.01032
R27194 vgaringosc.workerclkbuff_notouch_.I.n0 vgaringosc.workerclkbuff_notouch_.I.t2 2.01032
R27195 vgaringosc.workerclkbuff_notouch_.I.n1 vgaringosc.workerclkbuff_notouch_.I.t3 1.49844
R27196 vgaringosc.workerclkbuff_notouch_.I.n1 vgaringosc.workerclkbuff_notouch_.I.t1 1.49844
R27197 vgaringosc.workerclkbuff_notouch_.I vgaringosc.workerclkbuff_notouch_.I.n5 1.1478
R27198 a_41048_29816.n5 a_41048_29816.t16 15.7685
R27199 a_41048_29816.n6 a_41048_29816.t9 15.7685
R27200 a_41048_29816.n7 a_41048_29816.t18 15.7685
R27201 a_41048_29816.n8 a_41048_29816.t11 15.7685
R27202 a_41048_29816.n9 a_41048_29816.t8 15.7685
R27203 a_41048_29816.n10 a_41048_29816.t14 15.7685
R27204 a_41048_29816.n3 a_41048_29816.t20 15.7685
R27205 a_41048_29816.n4 a_41048_29816.t22 15.7685
R27206 a_41048_29816.n5 a_41048_29816.t15 11.6197
R27207 a_41048_29816.n6 a_41048_29816.t13 11.6197
R27208 a_41048_29816.n7 a_41048_29816.t17 11.6197
R27209 a_41048_29816.n8 a_41048_29816.t19 11.6197
R27210 a_41048_29816.n9 a_41048_29816.t7 11.6197
R27211 a_41048_29816.n10 a_41048_29816.t10 11.6197
R27212 a_41048_29816.n3 a_41048_29816.t12 11.6197
R27213 a_41048_29816.n4 a_41048_29816.t21 11.6197
R27214 a_41048_29816.n6 a_41048_29816.n5 10.5449
R27215 a_41048_29816.n7 a_41048_29816.n6 10.5449
R27216 a_41048_29816.n8 a_41048_29816.n7 10.5449
R27217 a_41048_29816.n9 a_41048_29816.n8 10.5449
R27218 a_41048_29816.n10 a_41048_29816.n9 10.5449
R27219 a_41048_29816.n4 a_41048_29816.n3 10.5449
R27220 a_41048_29816.n2 a_41048_29816.t4 10.4819
R27221 a_41048_29816.n11 a_41048_29816.n10 8.41578
R27222 a_41048_29816.n2 a_41048_29816.n1 7.31398
R27223 a_41048_29816.n14 a_41048_29816.n13 6.25311
R27224 a_41048_29816.n13 a_41048_29816.n0 5.37659
R27225 a_41048_29816.n1 a_41048_29816.t5 4.04494
R27226 a_41048_29816.n1 a_41048_29816.t6 4.04494
R27227 a_41048_29816.n0 a_41048_29816.t2 3.07367
R27228 a_41048_29816.n0 a_41048_29816.t0 3.07367
R27229 a_41048_29816.n14 a_41048_29816.t1 3.07367
R27230 a_41048_29816.t3 a_41048_29816.n14 3.07367
R27231 a_41048_29816.n11 a_41048_29816.n4 2.12967
R27232 a_41048_29816.n12 a_41048_29816.n11 1.98284
R27233 a_41048_29816.n13 a_41048_29816.n12 0.538543
R27234 a_41048_29816.n12 a_41048_29816.n2 0.415283
R27235 _355_.C.n12 _355_.C.n11 22.1361
R27236 _355_.C.n4 _355_.C.t14 18.6885
R27237 _355_.C.n20 _355_.C.t16 18.6885
R27238 _355_.C.n10 _355_.C.t11 18.6885
R27239 _355_.C.n9 _355_.C.t13 18.6885
R27240 _355_.C.n7 _355_.C.t6 17.703
R27241 _355_.C.n13 _355_.C.t5 17.5205
R27242 _355_.C.n6 _355_.C.t15 15.3305
R27243 _355_.C.n17 _355_.C.t20 15.3305
R27244 _355_.C.n15 _355_.C.t8 15.3305
R27245 _355_.C.n2 _355_.C.t19 15.3305
R27246 _355_.C.n17 _355_.C.t9 15.148
R27247 _355_.C.n2 _355_.C.t21 15.148
R27248 _355_.C.n6 _355_.C.t10 15.0872
R27249 _355_.C.n15 _355_.C.t22 15.0872
R27250 _355_.C.n7 _355_.C.t17 14.8195
R27251 _355_.C.n12 _355_.C 14.2057
R27252 _355_.C.n8 _355_.C 13.1405
R27253 _355_.C.n24 _355_.C.n3 12.9605
R27254 _355_.C.n25 _355_.C.n24 12.6005
R27255 _355_.C.n4 _355_.C.t23 11.9603
R27256 _355_.C.n20 _355_.C.t7 11.9603
R27257 _355_.C.n10 _355_.C.t12 11.9603
R27258 _355_.C.n9 _355_.C.t18 11.9603
R27259 _355_.C.n13 _355_.C.t4 11.5588
R27260 _355_.C.n8 _355_.C 10.2131
R27261 _355_.C.n16 _355_.C.n14 9.9005
R27262 _355_.C.n19 _355_.C.n16 9.1805
R27263 _355_.C.n19 _355_.C.n18 9.0005
R27264 _355_.C.n14 _355_.C 9.0005
R27265 _355_.C.n22 _355_.C.n8 8.9555
R27266 _355_.C _355_.C.n6 8.15932
R27267 _355_.C _355_.C.n15 8.15932
R27268 _355_.C _355_.C.n13 8.05312
R27269 _355_.C.n18 _355_.C.n17 8.01109
R27270 _355_.C.n3 _355_.C.n2 8.01109
R27271 _355_.C _355_.C.n7 8.00997
R27272 _355_.C.n25 _355_.C.n1 6.92347
R27273 _355_.C.n22 _355_.C.n19 6.6605
R27274 _355_.C.n23 _355_.C.n5 5.16795
R27275 _355_.C.n23 _355_.C.n22 4.8155
R27276 _355_.C.n22 _355_.C.n21 4.67295
R27277 _355_.C.n16 _355_.C 4.5005
R27278 _355_.C.n24 _355_.C.n23 4.5005
R27279 _355_.C _355_.C.n9 4.08607
R27280 _355_.C.n5 _355_.C.n4 4.0005
R27281 _355_.C.n21 _355_.C.n20 4.0005
R27282 _355_.C.n11 _355_.C.n10 4.0005
R27283 _355_.C _355_.C.n0 2.74964
R27284 _355_.C.n0 _355_.C.t0 2.06607
R27285 _355_.C.n1 _355_.C.t2 1.99806
R27286 _355_.C.n1 _355_.C.t3 1.99806
R27287 _355_.C.n14 _355_.C.n12 1.5305
R27288 _355_.C.n0 _355_.C.t1 1.4923
R27289 _355_.C.n11 _355_.C 0.245418
R27290 _355_.C.n18 _355_.C 0.148735
R27291 _355_.C.n3 _355_.C 0.148735
R27292 _355_.C _355_.C.n25 0.103357
R27293 _355_.C.n5 _355_.C 0.0860738
R27294 _355_.C.n21 _355_.C 0.0860738
R27295 a_42168_25640.n7 a_42168_25640.t10 9.93567
R27296 a_42168_25640.n1 a_42168_25640.t1 9.26067
R27297 a_42168_25640.n7 a_42168_25640.n6 6.3005
R27298 a_42168_25640.n1 a_42168_25640.n0 6.3005
R27299 a_42168_25640.n3 a_42168_25640.n2 6.3005
R27300 a_42168_25640.n5 a_42168_25640.n4 6.3005
R27301 a_42168_25640.n9 a_42168_25640.n8 6.3005
R27302 a_42168_25640.n4 a_42168_25640.t6 1.99806
R27303 a_42168_25640.n4 a_42168_25640.t7 1.99806
R27304 a_42168_25640.n2 a_42168_25640.t3 1.99806
R27305 a_42168_25640.n2 a_42168_25640.t2 1.99806
R27306 a_42168_25640.n0 a_42168_25640.t4 1.99806
R27307 a_42168_25640.n0 a_42168_25640.t5 1.99806
R27308 a_42168_25640.n6 a_42168_25640.t8 1.99806
R27309 a_42168_25640.n6 a_42168_25640.t9 1.99806
R27310 a_42168_25640.t0 a_42168_25640.n9 1.99806
R27311 a_42168_25640.n9 a_42168_25640.t11 1.99806
R27312 a_42168_25640.n8 a_42168_25640.n7 1.71833
R27313 a_42168_25640.n8 a_42168_25640.n5 0.963109
R27314 a_42168_25640.n3 a_42168_25640.n1 0.877022
R27315 a_42168_25640.n5 a_42168_25640.n3 0.877022
R27316 _230_.I.n12 _230_.I.t9 20.5135
R27317 _230_.I.n8 _230_.I.t6 20.4405
R27318 _230_.I.n1 _230_.I.t10 19.4185
R27319 _230_.I.n11 _230_.I.t3 18.5425
R27320 _230_.I.n7 _230_.I.n6 18.148
R27321 _230_.I.n4 _230_.I.t13 17.7395
R27322 _230_.I.n5 _230_.I.t7 17.5205
R27323 _230_.I.n0 _230_.I.t11 15.659
R27324 _230_.I.n8 _230_.I.t5 15.4035
R27325 _230_.I.n0 _230_.I.t8 14.6735
R27326 _230_.I.n11 _230_.I.t4 14.053
R27327 _230_.I.n4 _230_.I.t2 12.6782
R27328 _230_.I.n1 _230_.I.t12 11.6683
R27329 _230_.I.n5 _230_.I.t15 11.5588
R27330 _230_.I.n12 _230_.I.t14 11.4372
R27331 _230_.I.n9 _230_.I 10.4005
R27332 _230_.I.n3 _230_.I 10.3505
R27333 _230_.I.n3 _230_.I.n2 10.2605
R27334 _230_.I _230_.I.n11 9.08093
R27335 _230_.I.n15 _230_.I.t1 8.30886
R27336 _230_.I.n13 _230_.I.n12 8.26282
R27337 _230_.I _230_.I.n8 8.06925
R27338 _230_.I.n2 _230_.I.n1 8.0005
R27339 _230_.I _230_.I.n0 8.0005
R27340 _230_.I.n6 _230_.I.n5 8.0005
R27341 _230_.I.n9 _230_.I.n7 7.3805
R27342 _230_.I.n15 _230_.I.n14 6.7955
R27343 _230_.I.n7 _230_.I 4.6805
R27344 _230_.I.n14 _230_.I.n10 4.6805
R27345 _230_.I.n14 _230_.I.n13 4.5005
R27346 _230_.I _230_.I.t0 4.3844
R27347 _230_.I _230_.I.n4 4.07694
R27348 _230_.I.n10 _230_.I.n3 2.1605
R27349 _230_.I.n10 _230_.I.n9 0.9905
R27350 _230_.I.n13 _230_.I 0.702167
R27351 _230_.I _230_.I.n15 0.08114
R27352 _230_.I.n2 _230_.I 0.068
R27353 _230_.I.n6 _230_.I 0.0531154
R27354 _350_.A1.n4 _350_.A1 24.7357
R27355 _350_.A1.n6 _350_.A1.t10 20.9944
R27356 _350_.A1.n1 _350_.A1.t15 18.9805
R27357 _350_.A1.n0 _350_.A1.t5 18.6885
R27358 _350_.A1.n3 _350_.A1.t2 18.6885
R27359 _350_.A1.n7 _350_.A1.t14 18.3034
R27360 _350_.A1.n7 _350_.A1.n6 17.457
R27361 _350_.A1.n9 _350_.A1.t13 15.8868
R27362 _350_.A1.n8 _350_.A1.t7 14.8195
R27363 _350_.A1.n5 _350_.A1.t8 14.8195
R27364 _350_.A1.n11 _350_.A1.t6 14.8039
R27365 _350_.A1.n10 _350_.A1.n9 14.6005
R27366 _350_.A1.n10 _350_.A1.t3 13.9965
R27367 _350_.A1.n0 _350_.A1.t9 11.9603
R27368 _350_.A1.n3 _350_.A1.t12 11.9603
R27369 _350_.A1.n1 _350_.A1.t11 11.4372
R27370 _350_.A1.n6 _350_.A1.t4 11.133
R27371 _350_.A1.n2 _350_.A1 9.9905
R27372 _350_.A1.n2 _350_.A1 9.13858
R27373 _350_.A1 _350_.A1.n8 8.71206
R27374 _350_.A1 _350_.A1.t1 8.69622
R27375 _350_.A1.n13 _350_.A1.n5 8.27613
R27376 _350_.A1 _350_.A1.n1 8.11457
R27377 _350_.A1.n12 _350_.A1.n11 8.0005
R27378 _350_.A1.n14 _350_.A1.n13 7.2005
R27379 _350_.A1.n4 _350_.A1.n2 6.8405
R27380 _350_.A1 _350_.A1.t0 6.72245
R27381 _350_.A1 _350_.A1.n14 4.5005
R27382 _350_.A1 _350_.A1.n0 4.08607
R27383 _350_.A1 _350_.A1.n3 4.08607
R27384 _350_.A1.n8 _350_.A1.n7 2.7015
R27385 _350_.A1.n14 _350_.A1.n4 1.6205
R27386 _350_.A1.n9 _350_.A1.n5 1.5335
R27387 _350_.A1.n11 _350_.A1.n10 1.36925
R27388 _350_.A1.n12 _350_.A1 0.148156
R27389 _350_.A1.n13 _350_.A1.n12 0.0103438
R27390 _452_.CLK.n24 _452_.CLK 14.4005
R27391 _452_.CLK.n39 _452_.CLK.n36 14.2655
R27392 _452_.CLK.n50 _452_.CLK.t37 13.907
R27393 _452_.CLK.n40 _452_.CLK.t58 13.907
R27394 _452_.CLK.n28 _452_.CLK.t39 13.907
R27395 _452_.CLK.n25 _452_.CLK.t32 13.907
R27396 _452_.CLK.n42 _452_.CLK.t49 13.907
R27397 _452_.CLK.n31 _452_.CLK.n30 13.8605
R27398 _452_.CLK.n52 _452_.CLK.t44 13.8462
R27399 _452_.CLK.n47 _452_.CLK.t54 13.8462
R27400 _452_.CLK.n35 _452_.CLK.t45 13.8462
R27401 _452_.CLK.n32 _452_.CLK.t47 13.8462
R27402 _452_.CLK.n21 _452_.CLK.t53 13.8462
R27403 _452_.CLK.n22 _452_.CLK.t34 13.8462
R27404 _452_.CLK.n19 _452_.CLK.t59 13.8462
R27405 _452_.CLK.n37 _452_.CLK.t52 13.8462
R27406 _452_.CLK.n44 _452_.CLK.t48 13.8462
R27407 _452_.CLK.n43 _452_.CLK.n41 13.3205
R27408 _452_.CLK.n41 _452_.CLK.n39 12.9605
R27409 _452_.CLK.n52 _452_.CLK.t57 12.1185
R27410 _452_.CLK.n47 _452_.CLK.t40 12.1185
R27411 _452_.CLK.n35 _452_.CLK.t46 12.1185
R27412 _452_.CLK.n32 _452_.CLK.t56 12.1185
R27413 _452_.CLK.n21 _452_.CLK.t42 12.1185
R27414 _452_.CLK.n22 _452_.CLK.t41 12.1185
R27415 _452_.CLK.n19 _452_.CLK.t50 12.1185
R27416 _452_.CLK.n37 _452_.CLK.t36 12.1185
R27417 _452_.CLK.n44 _452_.CLK.t35 12.1185
R27418 _452_.CLK.n50 _452_.CLK.t33 12.0455
R27419 _452_.CLK.n40 _452_.CLK.t43 12.0455
R27420 _452_.CLK.n28 _452_.CLK.t55 12.0455
R27421 _452_.CLK.n25 _452_.CLK.t38 12.0455
R27422 _452_.CLK.n42 _452_.CLK.t51 12.0455
R27423 _452_.CLK.n30 _452_.CLK.n27 10.4405
R27424 _452_.CLK.n27 _452_.CLK.n26 10.3789
R27425 _452_.CLK.n46 _452_.CLK.n45 10.3789
R27426 _452_.CLK.n49 _452_.CLK.n46 9.5405
R27427 _452_.CLK.n24 _452_.CLK.n23 9.11892
R27428 _452_.CLK.n43 _452_.CLK 9.0005
R27429 _452_.CLK.n54 _452_.CLK.n53 8.2355
R27430 _452_.CLK _452_.CLK.n52 8.01471
R27431 _452_.CLK _452_.CLK.n50 8.01471
R27432 _452_.CLK _452_.CLK.n40 8.01471
R27433 _452_.CLK _452_.CLK.n35 8.01471
R27434 _452_.CLK _452_.CLK.n21 8.01471
R27435 _452_.CLK _452_.CLK.n42 8.01471
R27436 _452_.CLK.n48 _452_.CLK.n47 8.0005
R27437 _452_.CLK.n33 _452_.CLK.n32 8.0005
R27438 _452_.CLK.n29 _452_.CLK.n28 8.0005
R27439 _452_.CLK.n23 _452_.CLK.n22 8.0005
R27440 _452_.CLK.n26 _452_.CLK.n25 8.0005
R27441 _452_.CLK.n20 _452_.CLK.n19 8.0005
R27442 _452_.CLK.n38 _452_.CLK.n37 8.0005
R27443 _452_.CLK.n45 _452_.CLK.n44 8.0005
R27444 _452_.CLK.n61 _452_.CLK.n60 7.0655
R27445 _452_.CLK.n54 _452_.CLK.n18 6.67738
R27446 _452_.CLK.n57 _452_.CLK.n15 6.4355
R27447 _452_.CLK.n56 _452_.CLK.n16 6.4355
R27448 _452_.CLK.n55 _452_.CLK.n17 6.4355
R27449 _452_.CLK.n61 _452_.CLK.n59 6.4355
R27450 _452_.CLK.n62 _452_.CLK.n58 6.4355
R27451 _452_.CLK.n64 _452_.CLK.n63 6.4355
R27452 _452_.CLK.n39 _452_.CLK.n38 4.79892
R27453 _452_.CLK.n49 _452_.CLK.n48 4.61892
R27454 _452_.CLK.n34 _452_.CLK.n33 4.61892
R27455 _452_.CLK.n30 _452_.CLK.n29 4.61892
R27456 _452_.CLK.n31 _452_.CLK.n20 4.61892
R27457 _452_.CLK.n36 _452_.CLK 4.5005
R27458 _452_.CLK.n41 _452_.CLK 4.5005
R27459 _452_.CLK.n51 _452_.CLK 4.5005
R27460 _452_.CLK.n53 _452_.CLK 4.5005
R27461 _452_.CLK.n27 _452_.CLK.n24 4.1405
R27462 _452_.CLK.n36 _452_.CLK.n34 3.8255
R27463 _452_.CLK.n15 _452_.CLK.t12 3.37782
R27464 _452_.CLK.n15 _452_.CLK.t31 3.37782
R27465 _452_.CLK.n16 _452_.CLK.t13 3.37782
R27466 _452_.CLK.n16 _452_.CLK.t7 3.37782
R27467 _452_.CLK.n17 _452_.CLK.t22 3.37782
R27468 _452_.CLK.n17 _452_.CLK.t4 3.37782
R27469 _452_.CLK.n18 _452_.CLK.t23 3.37782
R27470 _452_.CLK.n18 _452_.CLK.t26 3.37782
R27471 _452_.CLK.n60 _452_.CLK.t19 3.37782
R27472 _452_.CLK.n60 _452_.CLK.t3 3.37782
R27473 _452_.CLK.n59 _452_.CLK.t17 3.37782
R27474 _452_.CLK.n59 _452_.CLK.t15 3.37782
R27475 _452_.CLK.n58 _452_.CLK.t29 3.37782
R27476 _452_.CLK.n58 _452_.CLK.t21 3.37782
R27477 _452_.CLK.n63 _452_.CLK.t30 3.37782
R27478 _452_.CLK.n63 _452_.CLK.t0 3.37782
R27479 _452_.CLK.n2 _452_.CLK.n0 2.94809
R27480 _452_.CLK.n9 _452_.CLK.n7 2.93257
R27481 _452_.CLK.n34 _452_.CLK.n31 2.7905
R27482 _452_.CLK.n6 _452_.CLK.n5 2.6005
R27483 _452_.CLK.n4 _452_.CLK.n3 2.6005
R27484 _452_.CLK.n2 _452_.CLK.n1 2.6005
R27485 _452_.CLK.n9 _452_.CLK.n8 2.6005
R27486 _452_.CLK.n11 _452_.CLK.n10 2.6005
R27487 _452_.CLK.n13 _452_.CLK.n12 2.6005
R27488 _452_.CLK.n12 _452_.CLK.t1 2.06607
R27489 _452_.CLK.n10 _452_.CLK.t2 2.06607
R27490 _452_.CLK.n8 _452_.CLK.t11 2.06607
R27491 _452_.CLK.n7 _452_.CLK.t18 2.06607
R27492 _452_.CLK.n0 _452_.CLK.t8 2.06607
R27493 _452_.CLK.n1 _452_.CLK.t9 2.06607
R27494 _452_.CLK.n3 _452_.CLK.t27 2.06607
R27495 _452_.CLK.n5 _452_.CLK.t28 2.06607
R27496 _452_.CLK.n53 _452_.CLK.n51 1.5305
R27497 _452_.CLK.n12 _452_.CLK.t5 1.4923
R27498 _452_.CLK.n10 _452_.CLK.t6 1.4923
R27499 _452_.CLK.n8 _452_.CLK.t16 1.4923
R27500 _452_.CLK.n7 _452_.CLK.t20 1.4923
R27501 _452_.CLK.n0 _452_.CLK.t14 1.4923
R27502 _452_.CLK.n1 _452_.CLK.t10 1.4923
R27503 _452_.CLK.n3 _452_.CLK.t24 1.4923
R27504 _452_.CLK.n5 _452_.CLK.t25 1.4923
R27505 _452_.CLK.n51 _452_.CLK.n49 1.2155
R27506 _452_.CLK.n46 _452_.CLK.n43 0.7205
R27507 _452_.CLK.n56 _452_.CLK.n55 0.6305
R27508 _452_.CLK.n57 _452_.CLK.n56 0.6305
R27509 _452_.CLK.n64 _452_.CLK.n62 0.6305
R27510 _452_.CLK.n62 _452_.CLK.n61 0.6305
R27511 _452_.CLK.n55 _452_.CLK.n54 0.388625
R27512 _452_.CLK.n6 _452_.CLK.n4 0.348086
R27513 _452_.CLK.n4 _452_.CLK.n2 0.348086
R27514 _452_.CLK.n11 _452_.CLK.n9 0.348086
R27515 _452_.CLK.n13 _452_.CLK.n11 0.348086
R27516 _452_.CLK.n65 _452_.CLK.n64 0.195969
R27517 _452_.CLK.n65 _452_.CLK.n57 0.181906
R27518 _452_.CLK.n14 _452_.CLK.n13 0.116103
R27519 _452_.CLK.n14 _452_.CLK.n6 0.0928276
R27520 _452_.CLK _452_.CLK.n14 0.0755
R27521 _452_.CLK _452_.CLK.n65 0.059
R27522 _452_.CLK.n48 _452_.CLK 0.0147105
R27523 _452_.CLK.n33 _452_.CLK 0.0147105
R27524 _452_.CLK.n29 _452_.CLK 0.0147105
R27525 _452_.CLK.n23 _452_.CLK 0.0147105
R27526 _452_.CLK.n26 _452_.CLK 0.0147105
R27527 _452_.CLK.n20 _452_.CLK 0.0147105
R27528 _452_.CLK.n38 _452_.CLK 0.0147105
R27529 _452_.CLK.n45 _452_.CLK 0.0147105
R27530 a_36548_27591.n0 a_36548_27591.t2 121.874
R27531 a_36548_27591.t2 a_36548_27591.t6 61.5152
R27532 a_36548_27591.n1 a_36548_27591.t4 52.378
R27533 a_36548_27591.n1 a_36548_27591.t3 17.7152
R27534 a_36548_27591.n3 a_36548_27591.t1 11.1158
R27535 a_36548_27591.n4 a_36548_27591.n0 9.95623
R27536 a_36548_27591.t0 a_36548_27591.n4 8.02846
R27537 a_36548_27591.n3 a_36548_27591.n2 8.0005
R27538 a_36548_27591.n0 a_36548_27591.t5 6.7165
R27539 a_36548_27591.n2 a_36548_27591.t7 6.023
R27540 a_36548_27591.n2 a_36548_27591.n1 1.33883
R27541 a_36548_27591.n4 a_36548_27591.n3 0.376152
R27542 _424_.B1.n3 _424_.B1.t8 19.4185
R27543 _424_.B1.n11 _424_.B1 19.0805
R27544 _424_.B1.n12 _424_.B1.n8 16.7405
R27545 _424_.B1.n3 _424_.B1.t10 16.535
R27546 _424_.B1.n8 _424_.B1.n7 16.1105
R27547 _424_.B1.n11 _424_.B1 15.9456
R27548 _424_.B1.n5 _424_.B1.t14 15.9023
R27549 _424_.B1.n6 _424_.B1.t15 15.9023
R27550 _424_.B1.n9 _424_.B1.t11 15.9023
R27551 _424_.B1.n10 _424_.B1.t9 15.9023
R27552 _424_.B1.n7 _424_.B1 14.0405
R27553 _424_.B1.n5 _424_.B1.t13 13.4447
R27554 _424_.B1.n6 _424_.B1.t7 13.4447
R27555 _424_.B1.n9 _424_.B1.t6 13.4447
R27556 _424_.B1.n10 _424_.B1.t12 13.4447
R27557 _424_.B1.n7 _424_.B1 11.2505
R27558 _424_.B1.n14 _424_.B1.n12 9.0005
R27559 _424_.B1 _424_.B1.n5 8.01083
R27560 _424_.B1 _424_.B1.n6 8.01083
R27561 _424_.B1 _424_.B1.n9 8.01083
R27562 _424_.B1 _424_.B1.n10 8.01083
R27563 _424_.B1.n4 _424_.B1.n3 8.0005
R27564 _424_.B1.n2 _424_.B1.n0 7.51504
R27565 _424_.B1.n12 _424_.B1.n11 6.6605
R27566 _424_.B1.n8 _424_.B1.n4 4.68238
R27567 _424_.B1.n2 _424_.B1.n1 2.71593
R27568 _424_.B1.n14 _424_.B1.n13 2.71425
R27569 _424_.B1.n0 _424_.B1.t4 1.99806
R27570 _424_.B1.n0 _424_.B1.t5 1.99806
R27571 _424_.B1.n13 _424_.B1.t3 1.61112
R27572 _424_.B1.n13 _424_.B1.t0 1.61112
R27573 _424_.B1.n1 _424_.B1.t1 1.61112
R27574 _424_.B1.n1 _424_.B1.t2 1.61112
R27575 _424_.B1 _424_.B1.n14 0.422375
R27576 _424_.B1.n4 _424_.B1 0.103625
R27577 _424_.B1 _424_.B1.n2 0.096125
R27578 _304_.A1.n12 _304_.A1.t9 24.9665
R27579 _304_.A1.n15 _304_.A1.t16 19.7835
R27580 _304_.A1.n8 _304_.A1.t7 19.2725
R27581 _304_.A1.n1 _304_.A1.t15 19.1995
R27582 _304_.A1.n10 _304_.A1.t5 18.6885
R27583 _304_.A1.n0 _304_.A1.t6 18.6885
R27584 _304_.A1.n4 _304_.A1.t10 16.8513
R27585 _304_.A1.n5 _304_.A1.t17 16.8513
R27586 _304_.A1.n5 _304_.A1.n4 16.5048
R27587 _304_.A1.n9 _304_.A1 14.3277
R27588 _304_.A1.n15 _304_.A1.t8 14.3085
R27589 _304_.A1.n8 _304_.A1.t3 13.8948
R27590 _304_.A1.n1 _304_.A1.t14 13.6637
R27591 _304_.A1.n10 _304_.A1.t13 11.9603
R27592 _304_.A1.n0 _304_.A1.t4 11.9603
R27593 _304_.A1.n3 _304_.A1.t12 11.5588
R27594 _304_.A1.n6 _304_.A1.t11 11.5588
R27595 _304_.A1.n16 _304_.A1 10.508
R27596 _304_.A1.n2 _304_.A1 9.9005
R27597 _304_.A1.n9 _304_.A1 9.5405
R27598 _304_.A1.n14 _304_.A1.n13 9.31815
R27599 _304_.A1.n2 _304_.A1 9.1805
R27600 _304_.A1.n11 _304_.A1 9.0005
R27601 _304_.A1.n12 _304_.A1.t2 8.73617
R27602 _304_.A1 _304_.A1.t1 8.69622
R27603 _304_.A1.n7 _304_.A1.n3 8.28737
R27604 _304_.A1 _304_.A1.n8 8.11085
R27605 _304_.A1.n7 _304_.A1.n6 8.0005
R27606 _304_.A1 _304_.A1.n15 8.0005
R27607 _304_.A1.n13 _304_.A1.n12 8.0005
R27608 _304_.A1 _304_.A1.n1 8.0005
R27609 _304_.A1 _304_.A1.t0 6.72245
R27610 _304_.A1.n17 _304_.A1.n2 6.4805
R27611 _304_.A1.n17 _304_.A1.n16 5.5805
R27612 _304_.A1 _304_.A1.n17 5.5355
R27613 _304_.A1 _304_.A1.n10 4.24542
R27614 _304_.A1 _304_.A1.n0 4.08607
R27615 _304_.A1.n11 _304_.A1.n9 3.8705
R27616 _304_.A1.n16 _304_.A1.n14 2.7005
R27617 _304_.A1.n14 _304_.A1.n11 1.4405
R27618 _304_.A1 _304_.A1.n7 0.950062
R27619 _304_.A1.n4 _304_.A1.n3 0.3655
R27620 _304_.A1.n6 _304_.A1.n5 0.3655
R27621 _304_.A1.n13 _304_.A1 0.0110882
R27622 a_54864_22461.n3 a_54864_22461.t2 121.874
R27623 a_54864_22461.t2 a_54864_22461.t5 61.5152
R27624 a_54864_22461.n0 a_54864_22461.t6 52.378
R27625 a_54864_22461.n0 a_54864_22461.t4 17.7882
R27626 a_54864_22461.n2 a_54864_22461.t1 11.1158
R27627 a_54864_22461.n4 a_54864_22461.n3 9.95623
R27628 a_54864_22461.t0 a_54864_22461.n4 8.02846
R27629 a_54864_22461.n2 a_54864_22461.n1 8.0005
R27630 a_54864_22461.n3 a_54864_22461.t7 6.7165
R27631 a_54864_22461.n1 a_54864_22461.t3 5.96217
R27632 a_54864_22461.n1 a_54864_22461.n0 1.33883
R27633 a_54864_22461.n4 a_54864_22461.n2 0.376152
R27634 _447_.Q.n11 _447_.Q.t17 24.9665
R27635 _447_.Q.n6 _447_.Q.t10 19.2725
R27636 _447_.Q.n16 _447_.Q.t15 19.1995
R27637 _447_.Q.n2 _447_.Q 19.0386
R27638 _447_.Q.n0 _447_.Q.t14 18.9805
R27639 _447_.Q.n1 _447_.Q.t5 18.9805
R27640 _447_.Q.n14 _447_.Q.t8 18.6885
R27641 _447_.Q.n9 _447_.Q.t13 18.6885
R27642 _447_.Q.n3 _447_.Q.t11 17.484
R27643 _447_.Q.n12 _447_.Q.n10 15.2061
R27644 _447_.Q.n6 _447_.Q.t16 13.8948
R27645 _447_.Q.n16 _447_.Q.t3 13.6637
R27646 _447_.Q.n2 _447_.Q 12.3305
R27647 _447_.Q.n9 _447_.Q.t6 11.9603
R27648 _447_.Q.n14 _447_.Q.t7 11.8873
R27649 _447_.Q.n3 _447_.Q.t4 11.863
R27650 _447_.Q.n0 _447_.Q.t12 11.4372
R27651 _447_.Q.n1 _447_.Q.t2 11.4372
R27652 _447_.Q.n17 _447_.Q 10.6205
R27653 _447_.Q _447_.Q.n17 9.5405
R27654 _447_.Q.n8 _447_.Q.n7 9.10336
R27655 _447_.Q.n5 _447_.Q.n4 9.0722
R27656 _447_.Q.n11 _447_.Q.t9 8.73617
R27657 _447_.Q _447_.Q.t1 8.69622
R27658 _447_.Q _447_.Q.n1 8.11576
R27659 _447_.Q _447_.Q.n0 8.11457
R27660 _447_.Q _447_.Q.n11 8.01109
R27661 _447_.Q.n4 _447_.Q.n3 8.0005
R27662 _447_.Q.n7 _447_.Q.n6 8.0005
R27663 _447_.Q _447_.Q.n16 8.0005
R27664 _447_.Q.n15 _447_.Q.n13 6.8405
R27665 _447_.Q _447_.Q.t0 6.72245
R27666 _447_.Q.n17 _447_.Q.n15 6.3005
R27667 _447_.Q.n13 _447_.Q.n12 5.7605
R27668 _447_.Q.n15 _447_.Q 4.66575
R27669 _447_.Q.n12 _447_.Q 4.64874
R27670 _447_.Q _447_.Q.n14 4.08607
R27671 _447_.Q.n10 _447_.Q.n9 4.0005
R27672 _447_.Q.n8 _447_.Q.n5 1.8005
R27673 _447_.Q.n13 _447_.Q.n8 1.1705
R27674 _447_.Q.n10 _447_.Q 0.245418
R27675 _447_.Q.n7 _447_.Q 0.107139
R27676 _447_.Q.n4 _447_.Q 0.0996525
R27677 _447_.Q.n5 _447_.Q.n2 0.0905
R27678 _350_.A2.n17 _350_.A2.t21 20.9576
R27679 _350_.A2.n21 _350_.A2.t22 19.5418
R27680 _350_.A2.n20 _350_.A2.t25 19.1995
R27681 _350_.A2.n16 _350_.A2.t26 17.7395
R27682 _350_.A2.n24 _350_.A2.t24 16.5472
R27683 _350_.A2.n27 _350_.A2.n26 15.6605
R27684 _350_.A2.n24 _350_.A2.t23 14.8925
R27685 _350_.A2.n16 _350_.A2.t28 12.6782
R27686 _350_.A2.n21 _350_.A2.n20 12.0614
R27687 _350_.A2.n19 _350_.A2.t29 9.673
R27688 _350_.A2.n26 _350_.A2 8.5955
R27689 _350_.A2 _350_.A2.n17 8.48925
R27690 _350_.A2.n22 _350_.A2.t27 8.45633
R27691 _350_.A2.n17 _350_.A2.t20 8.45633
R27692 _350_.A2.n25 _350_.A2.n24 8.00621
R27693 _350_.A2.n23 _350_.A2.n22 8.0005
R27694 _350_.A2.n19 _350_.A2.n18 8.0005
R27695 _350_.A2.n2 _350_.A2.n0 7.17702
R27696 _350_.A2.n4 _350_.A2.n3 6.3005
R27697 _350_.A2.n2 _350_.A2.n1 6.3005
R27698 _350_.A2.n6 _350_.A2.n5 6.3005
R27699 _350_.A2.n9 _350_.A2.n7 5.73397
R27700 _350_.A2.n26 _350_.A2.n25 5.4005
R27701 _350_.A2.n29 _350_.A2.n28 5.2005
R27702 _350_.A2.n9 _350_.A2.n8 5.2005
R27703 _350_.A2.n11 _350_.A2.n10 5.2005
R27704 _350_.A2.n13 _350_.A2.n12 5.2005
R27705 _350_.A2 _350_.A2.n16 4.07694
R27706 _350_.A2.n0 _350_.A2.t7 3.83001
R27707 _350_.A2.n5 _350_.A2.t5 3.83001
R27708 _350_.A2.n20 _350_.A2.n19 3.80867
R27709 _350_.A2.n22 _350_.A2.n21 2.67717
R27710 _350_.A2.n27 _350_.A2.n15 2.64381
R27711 _350_.A2.n1 _350_.A2.t4 1.99806
R27712 _350_.A2.n1 _350_.A2.t9 1.99806
R27713 _350_.A2.n3 _350_.A2.t11 1.99806
R27714 _350_.A2.n3 _350_.A2.t6 1.99806
R27715 _350_.A2.n10 _350_.A2.t16 1.84822
R27716 _350_.A2.n10 _350_.A2.t1 1.84822
R27717 _350_.A2.n8 _350_.A2.t2 1.84822
R27718 _350_.A2.n8 _350_.A2.t18 1.84822
R27719 _350_.A2.n7 _350_.A2.t17 1.84822
R27720 _350_.A2.n7 _350_.A2.t0 1.84822
R27721 _350_.A2.n12 _350_.A2.t3 1.84822
R27722 _350_.A2.n12 _350_.A2.t19 1.84822
R27723 _350_.A2.n0 _350_.A2.t15 1.70267
R27724 _350_.A2.n5 _350_.A2.t12 1.70267
R27725 _350_.A2.n28 _350_.A2.t8 1.6626
R27726 _350_.A2.n28 _350_.A2.t13 1.6626
R27727 _350_.A2.n15 _350_.A2.t14 1.6626
R27728 _350_.A2.n15 _350_.A2.t10 1.6626
R27729 _350_.A2.n29 _350_.A2.n27 1.23977
R27730 _350_.A2.n25 _350_.A2.n23 1.11368
R27731 _350_.A2.n14 _350_.A2.n6 0.985548
R27732 _350_.A2.n6 _350_.A2.n4 0.877022
R27733 _350_.A2.n4 _350_.A2.n2 0.877022
R27734 _350_.A2.n11 _350_.A2.n9 0.533966
R27735 _350_.A2.n13 _350_.A2.n11 0.533966
R27736 _350_.A2 _350_.A2.n29 0.388625
R27737 _350_.A2.n23 _350_.A2.n18 0.375194
R27738 _350_.A2.n18 _350_.A2 0.315321
R27739 _350_.A2 _350_.A2.n14 0.283766
R27740 _350_.A2.n14 _350_.A2.n13 0.227215
R27741 a_48272_25156.n22 a_48272_25156.t43 15.4765
R27742 a_48272_25156.n23 a_48272_25156.t14 15.4765
R27743 a_48272_25156.n24 a_48272_25156.t18 15.4765
R27744 a_48272_25156.n8 a_48272_25156.t17 15.4765
R27745 a_48272_25156.n9 a_48272_25156.t23 15.4765
R27746 a_48272_25156.n10 a_48272_25156.t20 15.4765
R27747 a_48272_25156.n11 a_48272_25156.t45 15.4765
R27748 a_48272_25156.n12 a_48272_25156.t42 15.4765
R27749 a_48272_25156.n13 a_48272_25156.t38 15.4765
R27750 a_48272_25156.n14 a_48272_25156.t40 15.4765
R27751 a_48272_25156.n15 a_48272_25156.t30 15.4765
R27752 a_48272_25156.n16 a_48272_25156.t34 15.4765
R27753 a_48272_25156.n17 a_48272_25156.t29 15.4765
R27754 a_48272_25156.n18 a_48272_25156.t25 15.4765
R27755 a_48272_25156.n21 a_48272_25156.t19 15.4765
R27756 a_48272_25156.n25 a_48272_25156.t15 15.4765
R27757 a_48272_25156.n22 a_48272_25156.t24 11.8022
R27758 a_48272_25156.n23 a_48272_25156.t27 11.8022
R27759 a_48272_25156.n24 a_48272_25156.t32 11.8022
R27760 a_48272_25156.n8 a_48272_25156.t31 11.8022
R27761 a_48272_25156.n9 a_48272_25156.t36 11.8022
R27762 a_48272_25156.n10 a_48272_25156.t35 11.8022
R27763 a_48272_25156.n11 a_48272_25156.t26 11.8022
R27764 a_48272_25156.n12 a_48272_25156.t22 11.8022
R27765 a_48272_25156.n13 a_48272_25156.t16 11.8022
R27766 a_48272_25156.n14 a_48272_25156.t21 11.8022
R27767 a_48272_25156.n15 a_48272_25156.t41 11.8022
R27768 a_48272_25156.n16 a_48272_25156.t44 11.8022
R27769 a_48272_25156.n17 a_48272_25156.t39 11.8022
R27770 a_48272_25156.n25 a_48272_25156.t28 11.8022
R27771 a_48272_25156.n19 a_48272_25156.t37 11.7413
R27772 a_48272_25156.n20 a_48272_25156.t33 11.7413
R27773 a_48272_25156.n5 a_48272_25156.t8 11.3584
R27774 a_48272_25156.n23 a_48272_25156.n22 10.5449
R27775 a_48272_25156.n24 a_48272_25156.n23 10.5449
R27776 a_48272_25156.n9 a_48272_25156.n8 10.5449
R27777 a_48272_25156.n10 a_48272_25156.n9 10.5449
R27778 a_48272_25156.n11 a_48272_25156.n10 10.5449
R27779 a_48272_25156.n12 a_48272_25156.n11 10.5449
R27780 a_48272_25156.n13 a_48272_25156.n12 10.5449
R27781 a_48272_25156.n14 a_48272_25156.n13 10.5449
R27782 a_48272_25156.n15 a_48272_25156.n14 10.5449
R27783 a_48272_25156.n16 a_48272_25156.n15 10.5449
R27784 a_48272_25156.n17 a_48272_25156.n16 10.5449
R27785 a_48272_25156.n18 a_48272_25156.n17 10.5449
R27786 a_48272_25156.n25 a_48272_25156.n21 10.5449
R27787 a_48272_25156.n25 a_48272_25156.n24 10.5449
R27788 a_48272_25156.n7 a_48272_25156.t9 10.4819
R27789 a_48272_25156.n20 a_48272_25156.n19 10.26
R27790 a_48272_25156.n6 a_48272_25156.n3 6.43746
R27791 a_48272_25156.n5 a_48272_25156.n4 6.43746
R27792 a_48272_25156.n30 a_48272_25156.n29 6.25311
R27793 a_48272_25156.n29 a_48272_25156.n0 5.37659
R27794 a_48272_25156.n28 a_48272_25156.n1 5.37659
R27795 a_48272_25156.n27 a_48272_25156.n2 5.37659
R27796 a_48272_25156.n3 a_48272_25156.t12 4.04494
R27797 a_48272_25156.n3 a_48272_25156.t10 4.04494
R27798 a_48272_25156.n4 a_48272_25156.t11 4.04494
R27799 a_48272_25156.n4 a_48272_25156.t13 4.04494
R27800 a_48272_25156.n0 a_48272_25156.t3 3.07367
R27801 a_48272_25156.n1 a_48272_25156.t4 3.07367
R27802 a_48272_25156.n2 a_48272_25156.t1 3.07367
R27803 a_48272_25156.n30 a_48272_25156.t6 3.07367
R27804 a_48272_25156.n0 a_48272_25156.t5 2.22001
R27805 a_48272_25156.n1 a_48272_25156.t2 2.22001
R27806 a_48272_25156.n2 a_48272_25156.t0 2.22001
R27807 a_48272_25156.t7 a_48272_25156.n30 2.22001
R27808 a_48272_25156.n26 a_48272_25156.n25 1.9195
R27809 a_48272_25156.n7 a_48272_25156.n6 0.877022
R27810 a_48272_25156.n6 a_48272_25156.n5 0.877022
R27811 a_48272_25156.n28 a_48272_25156.n27 0.877022
R27812 a_48272_25156.n29 a_48272_25156.n28 0.877022
R27813 a_48272_25156.n27 a_48272_25156.n26 0.430935
R27814 a_48272_25156.n26 a_48272_25156.n7 0.313543
R27815 a_48272_25156.n19 a_48272_25156.n18 0.0613333
R27816 a_48272_25156.n21 a_48272_25156.n20 0.0613333
R27817 _362_.B.n15 _362_.B.t17 22.3385
R27818 _362_.B.n10 _362_.B.t4 19.7835
R27819 _362_.B.n18 _362_.B.t14 18.6885
R27820 _362_.B.n12 _362_.B.t11 17.8003
R27821 _362_.B.n8 _362_.B.t18 17.2772
R27822 _362_.B.n14 _362_.B.t9 16.6445
R27823 _362_.B.n8 _362_.B.t12 16.5715
R27824 _362_.B.n3 _362_.B.t10 16.5715
R27825 _362_.B.n6 _362_.B.t15 16.5715
R27826 _362_.B.n1 _362_.B.t13 16.5715
R27827 _362_.B.n5 _362_.B.n4 16.5048
R27828 _362_.B.n1 _362_.B.t5 15.6468
R27829 _362_.B.n14 _362_.B.t21 15.4522
R27830 _362_.B.n12 _362_.B.t6 14.8195
R27831 _362_.B.n4 _362_.B.t16 14.7952
R27832 _362_.B.n5 _362_.B.t8 14.7952
R27833 _362_.B.n10 _362_.B.t19 14.3085
R27834 _362_.B.n18 _362_.B.t7 11.9603
R27835 _362_.B.n13 _362_.B 11.2596
R27836 _362_.B.n15 _362_.B.t20 9.75817
R27837 _362_.B _362_.B.n14 9.01391
R27838 _362_.B _362_.B.n1 8.11638
R27839 _362_.B _362_.B.n12 8.11418
R27840 _362_.B.n9 _362_.B.n8 8.05865
R27841 _362_.B _362_.B.n10 8.00997
R27842 _362_.B.n16 _362_.B.n15 8.0005
R27843 _362_.B.n7 _362_.B.n6 8.0005
R27844 _362_.B.n3 _362_.B.n2 8.0005
R27845 _362_.B.n20 _362_.B.n19 6.9755
R27846 _362_.B.n11 _362_.B.n9 6.9305
R27847 _362_.B.n13 _362_.B.n11 6.6605
R27848 _362_.B.n20 _362_.B.n0 6.35795
R27849 _362_.B _362_.B.n21 5.26469
R27850 _362_.B.n19 _362_.B 4.84575
R27851 _362_.B.n11 _362_.B 4.8155
R27852 _362_.B.n17 _362_.B.n16 4.7899
R27853 _362_.B.n17 _362_.B.n13 4.5005
R27854 _362_.B _362_.B.n18 4.08607
R27855 _362_.B.n4 _362_.B.n3 2.4825
R27856 _362_.B.n6 _362_.B.n5 2.4825
R27857 _362_.B.n0 _362_.B.t2 1.99806
R27858 _362_.B.n0 _362_.B.t3 1.99806
R27859 _362_.B.n21 _362_.B.t1 1.4923
R27860 _362_.B.n21 _362_.B.t0 1.4923
R27861 _362_.B.n9 _362_.B.n7 1.20982
R27862 _362_.B.n2 _362_.B 1.08463
R27863 _362_.B.n19 _362_.B.n17 0.6755
R27864 _362_.B _362_.B.n20 0.396829
R27865 _362_.B.n7 _362_.B.n2 0.39425
R27866 _362_.B.n16 _362_.B 0.0170789
R27867 a_42820_29159.n0 a_42820_29159.t7 121.874
R27868 a_42820_29159.t7 a_42820_29159.t4 61.5152
R27869 a_42820_29159.n2 a_42820_29159.t2 52.378
R27870 a_42820_29159.n2 a_42820_29159.t6 17.7152
R27871 a_42820_29159.t0 a_42820_29159.n4 11.1158
R27872 a_42820_29159.n1 a_42820_29159.n0 9.95623
R27873 a_42820_29159.n1 a_42820_29159.t1 8.02846
R27874 a_42820_29159.n4 a_42820_29159.n3 8.0005
R27875 a_42820_29159.n0 a_42820_29159.t5 6.7165
R27876 a_42820_29159.n3 a_42820_29159.t3 6.023
R27877 a_42820_29159.n3 a_42820_29159.n2 1.33883
R27878 a_42820_29159.n4 a_42820_29159.n1 0.376152
R27879 _371_.A1.n8 _371_.A1.t13 18.6885
R27880 _371_.A1.n9 _371_.A1.n7 16.9205
R27881 _371_.A1.n12 _371_.A1.t11 16.7418
R27882 _371_.A1.n13 _371_.A1.t18 16.7418
R27883 _371_.A1.n10 _371_.A1.t9 15.7077
R27884 _371_.A1.n18 _371_.A1.t16 15.7077
R27885 _371_.A1.n6 _371_.A1.t17 15.3305
R27886 _371_.A1.n6 _371_.A1.t8 15.148
R27887 _371_.A1.n21 _371_.A1.n20 14.4005
R27888 _371_.A1.n17 _371_.A1.n16 13.3198
R27889 _371_.A1.n13 _371_.A1.n12 13.3198
R27890 _371_.A1.n16 _371_.A1.t15 12.0455
R27891 _371_.A1.n17 _371_.A1.t12 12.0455
R27892 _371_.A1.n8 _371_.A1.t14 11.8873
R27893 _371_.A1.n20 _371_.A1 10.7105
R27894 _371_.A1.n20 _371_.A1.n9 8.6405
R27895 _371_.A1.n15 _371_.A1.n11 8.43876
R27896 _371_.A1.n11 _371_.A1.t19 8.3955
R27897 _371_.A1.n14 _371_.A1.t10 8.3955
R27898 _371_.A1 _371_.A1.n10 8.20879
R27899 _371_.A1.n7 _371_.A1.n6 8.01109
R27900 _371_.A1.n15 _371_.A1.n14 8.0005
R27901 _371_.A1.n19 _371_.A1.n18 8.0005
R27902 _371_.A1 _371_.A1.n0 6.79383
R27903 _371_.A1.n3 _371_.A1.n1 5.98178
R27904 _371_.A1.n5 _371_.A1.n4 5.2005
R27905 _371_.A1.n3 _371_.A1.n2 5.2005
R27906 _371_.A1.n9 _371_.A1 4.66575
R27907 _371_.A1 _371_.A1.n8 4.08607
R27908 _371_.A1.n12 _371_.A1.n11 3.6505
R27909 _371_.A1.n14 _371_.A1.n13 3.6505
R27910 _371_.A1.n0 _371_.A1.t2 1.99806
R27911 _371_.A1.n0 _371_.A1.t3 1.99806
R27912 _371_.A1.n4 _371_.A1.t7 1.84822
R27913 _371_.A1.n4 _371_.A1.t4 1.84822
R27914 _371_.A1.n1 _371_.A1.t5 1.84822
R27915 _371_.A1.n1 _371_.A1.t6 1.84822
R27916 _371_.A1.n2 _371_.A1.t1 1.84822
R27917 _371_.A1.n2 _371_.A1.t0 1.84822
R27918 _371_.A1.n19 _371_.A1.n15 1.34296
R27919 _371_.A1.n21 _371_.A1.n5 1.2458
R27920 _371_.A1.n16 _371_.A1.n10 1.03467
R27921 _371_.A1.n18 _371_.A1.n17 1.03467
R27922 _371_.A1.n5 _371_.A1.n3 0.781777
R27923 _371_.A1 _371_.A1.n21 0.187167
R27924 _371_.A1.n7 _371_.A1 0.148735
R27925 _371_.A1 _371_.A1.n19 0.0545
R27926 _397_.A2.n9 _397_.A2.t15 20.2215
R27927 _397_.A2.n10 _397_.A2.t6 20.2215
R27928 _397_.A2.n12 _397_.A2.t21 19.4185
R27929 _397_.A2.n17 _397_.A2.n13 19.0374
R27930 _397_.A2.n6 _397_.A2.t11 18.9805
R27931 _397_.A2.n10 _397_.A2.n9 18.9805
R27932 _397_.A2.n4 _397_.A2.t19 17.5205
R27933 _397_.A2.n12 _397_.A2.t5 16.535
R27934 _397_.A2.n20 _397_.A2.t17 16.2795
R27935 _397_.A2.n2 _397_.A2.t12 16.2795
R27936 _397_.A2.n15 _397_.A2.t16 15.5008
R27937 _397_.A2.n20 _397_.A2.t8 15.2818
R27938 _397_.A2.n2 _397_.A2.t10 15.2818
R27939 _397_.A2.n14 _397_.A2.t9 14.8317
R27940 _397_.A2.n14 _397_.A2.t13 13.8705
R27941 _397_.A2.n15 _397_.A2.t4 13.2013
R27942 _397_.A2.n4 _397_.A2.t7 11.5588
R27943 _397_.A2.n6 _397_.A2.t20 11.4372
R27944 _397_.A2.n7 _397_.A2.n5 10.723
R27945 _397_.A2.n21 _397_.A2 10.5437
R27946 _397_.A2 _397_.A2.n14 9.04897
R27947 _397_.A2.n7 _397_.A2 9.0005
R27948 _397_.A2.n8 _397_.A2.t18 8.74833
R27949 _397_.A2.n11 _397_.A2.t14 8.74833
R27950 _397_.A2 _397_.A2.n11 8.27205
R27951 _397_.A2 _397_.A2.n20 8.17653
R27952 _397_.A2 _397_.A2.n6 8.11576
R27953 _397_.A2 _397_.A2.n8 8.04395
R27954 _397_.A2.n3 _397_.A2.n2 8.02829
R27955 _397_.A2.n5 _397_.A2.n4 8.0005
R27956 _397_.A2.n16 _397_.A2.n15 8.0005
R27957 _397_.A2.n13 _397_.A2.n12 8.0005
R27958 _397_.A2.n23 _397_.A2.n22 7.4705
R27959 _397_.A2.n23 _397_.A2.n1 6.35795
R27960 _397_.A2.n22 _397_.A2.n3 6.2555
R27961 _397_.A2.n19 _397_.A2.n18 6.0755
R27962 _397_.A2 _397_.A2.n0 5.26469
R27963 _397_.A2.n17 _397_.A2.n16 4.5815
R27964 _397_.A2.n18 _397_.A2 4.5005
R27965 _397_.A2.n22 _397_.A2.n21 4.5005
R27966 _397_.A2.n9 _397_.A2.n8 3.0665
R27967 _397_.A2.n11 _397_.A2.n10 3.0665
R27968 _397_.A2.n18 _397_.A2.n17 2.9705
R27969 _397_.A2.n1 _397_.A2.t2 1.99806
R27970 _397_.A2.n1 _397_.A2.t3 1.99806
R27971 _397_.A2.n0 _397_.A2.t1 1.4923
R27972 _397_.A2.n0 _397_.A2.t0 1.4923
R27973 _397_.A2.n21 _397_.A2.n19 1.3505
R27974 _397_.A2.n19 _397_.A2.n7 1.2605
R27975 _397_.A2 _397_.A2.n23 0.396829
R27976 _397_.A2.n3 _397_.A2 0.148735
R27977 _397_.A2.n13 _397_.A2 0.103625
R27978 _397_.A2.n5 _397_.A2 0.0531154
R27979 _397_.A2.n16 _397_.A2 0.0199245
R27980 _284_.ZN.n39 _284_.ZN.t31 28.7301
R27981 _284_.ZN.n37 _284_.ZN.n25 25.7405
R27982 _284_.ZN.n33 _284_.ZN.n32 18.9805
R27983 _284_.ZN.n28 _284_.ZN.n27 18.9805
R27984 _284_.ZN.n44 _284_.ZN.n43 18.9805
R27985 _284_.ZN.n2 _284_.ZN.n1 18.9805
R27986 _284_.ZN.n38 _284_.ZN.t34 18.7615
R27987 _284_.ZN.n33 _284_.ZN.t29 15.2088
R27988 _284_.ZN.n32 _284_.ZN.t24 15.2088
R27989 _284_.ZN.n27 _284_.ZN.t22 15.2088
R27990 _284_.ZN.n28 _284_.ZN.t36 15.2088
R27991 _284_.ZN.n43 _284_.ZN.t23 15.2088
R27992 _284_.ZN.n44 _284_.ZN.t26 15.2088
R27993 _284_.ZN.n1 _284_.ZN.t37 15.2088
R27994 _284_.ZN.n2 _284_.ZN.t35 15.2088
R27995 _284_.ZN.n34 _284_.ZN.t28 14.7222
R27996 _284_.ZN.n31 _284_.ZN.t33 14.7222
R27997 _284_.ZN.n26 _284_.ZN.t21 14.7222
R27998 _284_.ZN.n29 _284_.ZN.t30 14.7222
R27999 _284_.ZN.n42 _284_.ZN.t27 14.7222
R28000 _284_.ZN.n45 _284_.ZN.t38 14.7222
R28001 _284_.ZN.n0 _284_.ZN.t32 14.7222
R28002 _284_.ZN.n3 _284_.ZN.t20 14.7222
R28003 _284_.ZN.n38 _284_.ZN.t25 13.4447
R28004 _284_.ZN.n40 _284_.ZN.n37 11.5205
R28005 _284_.ZN.n35 _284_.ZN.n31 8.34081
R28006 _284_.ZN.n30 _284_.ZN.n26 8.33378
R28007 _284_.ZN.n4 _284_.ZN.n0 8.33378
R28008 _284_.ZN.n42 _284_.ZN.n41 8.03988
R28009 _284_.ZN.n30 _284_.ZN.n29 8.0005
R28010 _284_.ZN.n35 _284_.ZN.n34 8.0005
R28011 _284_.ZN.n4 _284_.ZN.n3 8.0005
R28012 _284_.ZN.n46 _284_.ZN.n45 8.0005
R28013 _284_.ZN.n10 _284_.ZN.n8 7.17702
R28014 _284_.ZN.n10 _284_.ZN.n9 6.3005
R28015 _284_.ZN.n12 _284_.ZN.n11 6.3005
R28016 _284_.ZN.n16 _284_.ZN.n15 6.3005
R28017 _284_.ZN.n41 _284_.ZN.n40 5.7605
R28018 _284_.ZN.n20 _284_.ZN.n18 5.73397
R28019 _284_.ZN.n7 _284_.ZN.n6 5.2005
R28020 _284_.ZN.n20 _284_.ZN.n19 5.2005
R28021 _284_.ZN.n22 _284_.ZN.n21 5.2005
R28022 _284_.ZN.n24 _284_.ZN.n23 5.2005
R28023 _284_.ZN.n40 _284_.ZN 4.63313
R28024 _284_.ZN.n37 _284_.ZN.n36 4.5005
R28025 _284_.ZN.n7 _284_.ZN.n5 3.88308
R28026 _284_.ZN.n8 _284_.ZN.t1 3.83001
R28027 _284_.ZN _284_.ZN.n39 2.69796
R28028 _284_.ZN.n15 _284_.ZN.n14 2.53863
R28029 _284_.ZN.n11 _284_.ZN.t2 1.99806
R28030 _284_.ZN.n11 _284_.ZN.t10 1.99806
R28031 _284_.ZN.n9 _284_.ZN.t9 1.99806
R28032 _284_.ZN.n9 _284_.ZN.t3 1.99806
R28033 _284_.ZN.n23 _284_.ZN.t16 1.84822
R28034 _284_.ZN.n23 _284_.ZN.t7 1.84822
R28035 _284_.ZN.n21 _284_.ZN.t4 1.84822
R28036 _284_.ZN.n21 _284_.ZN.t18 1.84822
R28037 _284_.ZN.n19 _284_.ZN.t19 1.84822
R28038 _284_.ZN.n19 _284_.ZN.t6 1.84822
R28039 _284_.ZN.n18 _284_.ZN.t5 1.84822
R28040 _284_.ZN.n18 _284_.ZN.t17 1.84822
R28041 _284_.ZN.n8 _284_.ZN.t8 1.70267
R28042 _284_.ZN.n15 _284_.ZN.t11 1.70267
R28043 _284_.ZN.n6 _284_.ZN.t12 1.6626
R28044 _284_.ZN.n6 _284_.ZN.t15 1.6626
R28045 _284_.ZN.n5 _284_.ZN.t13 1.6626
R28046 _284_.ZN.n5 _284_.ZN.t14 1.6626
R28047 _284_.ZN.n14 _284_.ZN.t0 1.29188
R28048 _284_.ZN.n34 _284_.ZN.n33 1.0955
R28049 _284_.ZN.n32 _284_.ZN.n31 1.0955
R28050 _284_.ZN.n27 _284_.ZN.n26 1.0955
R28051 _284_.ZN.n29 _284_.ZN.n28 1.0955
R28052 _284_.ZN.n43 _284_.ZN.n42 1.0955
R28053 _284_.ZN.n45 _284_.ZN.n44 1.0955
R28054 _284_.ZN.n1 _284_.ZN.n0 1.0955
R28055 _284_.ZN.n3 _284_.ZN.n2 1.0955
R28056 _284_.ZN.n39 _284_.ZN.n38 1.01439
R28057 _284_.ZN.n17 _284_.ZN.n16 0.985548
R28058 _284_.ZN.n14 _284_.ZN.n13 0.9455
R28059 _284_.ZN.n12 _284_.ZN.n10 0.877022
R28060 _284_.ZN.n16 _284_.ZN.n12 0.877022
R28061 _284_.ZN.n22 _284_.ZN.n20 0.533966
R28062 _284_.ZN.n24 _284_.ZN.n22 0.533966
R28063 _284_.ZN _284_.ZN.n35 0.487062
R28064 _284_.ZN _284_.ZN.n46 0.487062
R28065 _284_.ZN _284_.ZN.n4 0.43925
R28066 _284_.ZN _284_.ZN.n7 0.388625
R28067 _284_.ZN.n36 _284_.ZN 0.3155
R28068 _284_.ZN.n46 _284_.ZN.n41 0.301438
R28069 _284_.ZN.n17 _284_.ZN 0.283766
R28070 _284_.ZN.n36 _284_.ZN.n30 0.12425
R28071 _284_.ZN.n25 _284_.ZN.n17 0.122046
R28072 _284_.ZN.n25 _284_.ZN.n24 0.105669
R28073 uo_out[0].n10 uo_out[0] 15.2626
R28074 uo_out[0].n5 uo_out[0].n4 7.21811
R28075 uo_out[0].n5 uo_out[0].n3 6.36507
R28076 uo_out[0].n6 uo_out[0].n2 6.36507
R28077 uo_out[0].n7 uo_out[0].n1 6.36507
R28078 uo_out[0].n10 uo_out[0].n9 3.01668
R28079 uo_out[0].n4 uo_out[0].t11 2.89962
R28080 uo_out[0].n4 uo_out[0].t0 2.89962
R28081 uo_out[0].n3 uo_out[0].t2 2.89962
R28082 uo_out[0].n3 uo_out[0].t10 2.89962
R28083 uo_out[0].n2 uo_out[0].t9 2.89962
R28084 uo_out[0].n2 uo_out[0].t1 2.89962
R28085 uo_out[0].n1 uo_out[0].t3 2.89962
R28086 uo_out[0].n1 uo_out[0].t8 2.89962
R28087 uo_out[0].n8 uo_out[0].n0 2.70811
R28088 uo_out[0].n0 uo_out[0].t7 2.06607
R28089 uo_out[0].n0 uo_out[0].t4 2.06607
R28090 uo_out[0].n9 uo_out[0].t5 2.06607
R28091 uo_out[0].n9 uo_out[0].t6 2.06607
R28092 uo_out[0].n8 uo_out[0].n7 1.50799
R28093 uo_out[0].n7 uo_out[0].n6 0.877022
R28094 uo_out[0].n6 uo_out[0].n5 0.877022
R28095 uo_out[0] uo_out[0].n10 0.800488
R28096 uo_out[0] uo_out[0].n8 0.267929
R28097 a_43440_19325.n3 a_43440_19325.t4 121.874
R28098 a_43440_19325.t4 a_43440_19325.t2 61.5152
R28099 a_43440_19325.n0 a_43440_19325.t3 52.378
R28100 a_43440_19325.n0 a_43440_19325.t7 17.7882
R28101 a_43440_19325.n2 a_43440_19325.t1 11.1158
R28102 a_43440_19325.n4 a_43440_19325.n3 9.95623
R28103 a_43440_19325.t0 a_43440_19325.n4 8.02846
R28104 a_43440_19325.n2 a_43440_19325.n1 8.0005
R28105 a_43440_19325.n3 a_43440_19325.t5 6.7165
R28106 a_43440_19325.n1 a_43440_19325.t6 5.96217
R28107 a_43440_19325.n1 a_43440_19325.n0 1.33883
R28108 a_43440_19325.n4 a_43440_19325.n2 0.376152
R28109 _459_.CLK.n11 _459_.CLK.t50 20.2337
R28110 _459_.CLK.n40 _459_.CLK.n37 19.0189
R28111 _459_.CLK.n28 _459_.CLK 17.9605
R28112 _459_.CLK.n15 _459_.CLK.n12 16.3897
R28113 _459_.CLK.n52 _459_.CLK 15.5255
R28114 _459_.CLK.n33 _459_.CLK.n32 13.9505
R28115 _459_.CLK.n53 _459_.CLK.t35 13.907
R28116 _459_.CLK.n10 _459_.CLK.t25 13.907
R28117 _459_.CLK.n21 _459_.CLK.t29 13.907
R28118 _459_.CLK.n30 _459_.CLK.t17 13.907
R28119 _459_.CLK.n42 _459_.CLK.t46 13.907
R28120 _459_.CLK.n48 _459_.CLK.t41 13.907
R28121 _459_.CLK.n36 _459_.CLK.t48 13.907
R28122 _459_.CLK.n9 _459_.CLK.t47 13.8462
R28123 _459_.CLK.n13 _459_.CLK.t19 13.8462
R28124 _459_.CLK.n26 _459_.CLK.t39 13.8462
R28125 _459_.CLK.n25 _459_.CLK.t18 13.8462
R28126 _459_.CLK.n23 _459_.CLK.t43 13.8462
R28127 _459_.CLK.n16 _459_.CLK.t23 13.8462
R28128 _459_.CLK.n18 _459_.CLK.t24 13.8462
R28129 _459_.CLK.n45 _459_.CLK.t22 13.8462
R28130 _459_.CLK.n38 _459_.CLK.t34 13.8462
R28131 _459_.CLK.n51 _459_.CLK.t20 13.8462
R28132 _459_.CLK.n34 _459_.CLK.n33 12.6005
R28133 _459_.CLK.n35 _459_.CLK.n34 12.4205
R28134 _459_.CLK.n9 _459_.CLK.t51 12.1185
R28135 _459_.CLK.n13 _459_.CLK.t33 12.1185
R28136 _459_.CLK.n26 _459_.CLK.t45 12.1185
R28137 _459_.CLK.n25 _459_.CLK.t42 12.1185
R28138 _459_.CLK.n23 _459_.CLK.t21 12.1185
R28139 _459_.CLK.n16 _459_.CLK.t37 12.1185
R28140 _459_.CLK.n18 _459_.CLK.t16 12.1185
R28141 _459_.CLK.n45 _459_.CLK.t36 12.1185
R28142 _459_.CLK.n38 _459_.CLK.t30 12.1185
R28143 _459_.CLK.n51 _459_.CLK.t40 12.1185
R28144 _459_.CLK.n53 _459_.CLK.t26 12.0455
R28145 _459_.CLK.n10 _459_.CLK.t44 12.0455
R28146 _459_.CLK.n21 _459_.CLK.t31 12.0455
R28147 _459_.CLK.n30 _459_.CLK.t28 12.0455
R28148 _459_.CLK.n42 _459_.CLK.t32 12.0455
R28149 _459_.CLK.n48 _459_.CLK.t38 12.0455
R28150 _459_.CLK.n36 _459_.CLK.t27 12.0455
R28151 _459_.CLK.n55 _459_.CLK 11.8805
R28152 _459_.CLK.n29 _459_.CLK.n24 11.2855
R28153 _459_.CLK.n11 _459_.CLK.t49 10.8288
R28154 _459_.CLK.n41 _459_.CLK.n40 10.7555
R28155 _459_.CLK.n47 _459_.CLK.n46 10.3789
R28156 _459_.CLK.n32 _459_.CLK.n29 10.3505
R28157 _459_.CLK.n55 _459_.CLK.n54 9.1805
R28158 _459_.CLK.n44 _459_.CLK.n43 9.11892
R28159 _459_.CLK.n50 _459_.CLK.n49 9.11892
R28160 _459_.CLK.n54 _459_.CLK 9.0005
R28161 _459_.CLK.n41 _459_.CLK.n35 9.0005
R28162 _459_.CLK _459_.CLK.n25 8.0155
R28163 _459_.CLK _459_.CLK.n9 8.01471
R28164 _459_.CLK _459_.CLK.n53 8.01471
R28165 _459_.CLK _459_.CLK.n10 8.01471
R28166 _459_.CLK _459_.CLK.n51 8.01471
R28167 _459_.CLK.n14 _459_.CLK.n13 8.0005
R28168 _459_.CLK.n12 _459_.CLK.n11 8.0005
R28169 _459_.CLK.n22 _459_.CLK.n21 8.0005
R28170 _459_.CLK.n31 _459_.CLK.n30 8.0005
R28171 _459_.CLK.n27 _459_.CLK.n26 8.0005
R28172 _459_.CLK.n24 _459_.CLK.n23 8.0005
R28173 _459_.CLK.n17 _459_.CLK.n16 8.0005
R28174 _459_.CLK.n19 _459_.CLK.n18 8.0005
R28175 _459_.CLK.n43 _459_.CLK.n42 8.0005
R28176 _459_.CLK.n49 _459_.CLK.n48 8.0005
R28177 _459_.CLK.n46 _459_.CLK.n45 8.0005
R28178 _459_.CLK.n39 _459_.CLK.n38 8.0005
R28179 _459_.CLK.n37 _459_.CLK.n36 8.0005
R28180 _459_.CLK.n20 _459_.CLK.n19 7.45392
R28181 _459_.CLK.n29 _459_.CLK.n28 7.2005
R28182 _459_.CLK.n5 _459_.CLK.n4 7.13263
R28183 _459_.CLK.n2 _459_.CLK.n1 7.13263
R28184 _459_.CLK.n5 _459_.CLK.n3 6.43746
R28185 _459_.CLK.n2 _459_.CLK.n0 6.43746
R28186 _459_.CLK.n56 _459_.CLK 5.7605
R28187 _459_.CLK.n57 _459_.CLK.n56 5.7155
R28188 _459_.CLK.n54 _459_.CLK.n52 5.4005
R28189 _459_.CLK.n40 _459_.CLK.n39 5.15892
R28190 _459_.CLK.n28 _459_.CLK.n27 4.6255
R28191 _459_.CLK.n15 _459_.CLK.n14 4.61892
R28192 _459_.CLK.n33 _459_.CLK.n22 4.61892
R28193 _459_.CLK.n32 _459_.CLK.n31 4.61892
R28194 _459_.CLK.n20 _459_.CLK.n17 4.61892
R28195 _459_.CLK.n56 _459_.CLK.n55 4.5005
R28196 _459_.CLK.n50 _459_.CLK.n47 4.3205
R28197 _459_.CLK.n4 _459_.CLK.t13 3.8098
R28198 _459_.CLK.n4 _459_.CLK.t8 3.8098
R28199 _459_.CLK.n3 _459_.CLK.t14 3.8098
R28200 _459_.CLK.n3 _459_.CLK.t15 3.8098
R28201 _459_.CLK.n0 _459_.CLK.t9 3.8098
R28202 _459_.CLK.n0 _459_.CLK.t10 3.8098
R28203 _459_.CLK.n1 _459_.CLK.t12 3.8098
R28204 _459_.CLK.n1 _459_.CLK.t11 3.8098
R28205 _459_.CLK.n61 _459_.CLK.n59 3.34593
R28206 _459_.CLK.n57 _459_.CLK.n8 2.78906
R28207 _459_.CLK.n58 _459_.CLK.n7 2.71593
R28208 _459_.CLK.n61 _459_.CLK.n60 2.71593
R28209 _459_.CLK.n8 _459_.CLK.t6 2.06607
R28210 _459_.CLK.n8 _459_.CLK.t3 2.06607
R28211 _459_.CLK.n7 _459_.CLK.t5 2.06607
R28212 _459_.CLK.n7 _459_.CLK.t2 2.06607
R28213 _459_.CLK.n59 _459_.CLK.t1 2.06607
R28214 _459_.CLK.n59 _459_.CLK.t0 2.06607
R28215 _459_.CLK.n60 _459_.CLK.t4 2.06607
R28216 _459_.CLK.n60 _459_.CLK.t7 2.06607
R28217 _459_.CLK.n47 _459_.CLK.n44 1.9805
R28218 _459_.CLK.n35 _459_.CLK.n15 1.2605
R28219 _459_.CLK.n34 _459_.CLK.n20 1.2155
R28220 _459_.CLK.n58 _459_.CLK.n57 0.557375
R28221 _459_.CLK.n52 _459_.CLK.n50 0.5405
R28222 _459_.CLK.n44 _459_.CLK.n41 0.5405
R28223 _459_.CLK.n6 _459_.CLK.n5 0.382224
R28224 _459_.CLK.n62 _459_.CLK.n61 0.346437
R28225 _459_.CLK.n6 _459_.CLK.n2 0.196017
R28226 _459_.CLK.n62 _459_.CLK.n58 0.177688
R28227 _459_.CLK _459_.CLK.n6 0.141421
R28228 _459_.CLK _459_.CLK.n62 0.133132
R28229 _459_.CLK.n12 _459_.CLK 0.065101
R28230 _459_.CLK.n27 _459_.CLK 0.0155
R28231 _459_.CLK.n24 _459_.CLK 0.0155
R28232 _459_.CLK.n14 _459_.CLK 0.0147105
R28233 _459_.CLK.n22 _459_.CLK 0.0147105
R28234 _459_.CLK.n31 _459_.CLK 0.0147105
R28235 _459_.CLK.n17 _459_.CLK 0.0147105
R28236 _459_.CLK.n19 _459_.CLK 0.0147105
R28237 _459_.CLK.n43 _459_.CLK 0.0147105
R28238 _459_.CLK.n49 _459_.CLK 0.0147105
R28239 _459_.CLK.n46 _459_.CLK 0.0147105
R28240 _459_.CLK.n39 _459_.CLK 0.0147105
R28241 _459_.CLK.n37 _459_.CLK 0.0147105
R28242 a_45284_19751.n0 a_45284_19751.t7 121.874
R28243 a_45284_19751.t7 a_45284_19751.t6 61.5152
R28244 a_45284_19751.n1 a_45284_19751.t5 52.378
R28245 a_45284_19751.n1 a_45284_19751.t4 17.7152
R28246 a_45284_19751.n3 a_45284_19751.t1 11.1158
R28247 a_45284_19751.n4 a_45284_19751.n0 9.95623
R28248 a_45284_19751.t0 a_45284_19751.n4 8.02846
R28249 a_45284_19751.n3 a_45284_19751.n2 8.0005
R28250 a_45284_19751.n0 a_45284_19751.t3 6.7165
R28251 a_45284_19751.n2 a_45284_19751.t2 6.023
R28252 a_45284_19751.n2 a_45284_19751.n1 1.33883
R28253 a_45284_19751.n4 a_45284_19751.n3 0.376152
R28254 a_23668_25640.n3 a_23668_25640.t7 121.874
R28255 a_23668_25640.t7 a_23668_25640.t6 61.5152
R28256 a_23668_25640.n0 a_23668_25640.t5 52.378
R28257 a_23668_25640.n0 a_23668_25640.t3 17.7882
R28258 a_23668_25640.n2 a_23668_25640.t1 11.1158
R28259 a_23668_25640.n4 a_23668_25640.n3 9.95623
R28260 a_23668_25640.t0 a_23668_25640.n4 8.02846
R28261 a_23668_25640.n2 a_23668_25640.n1 8.0005
R28262 a_23668_25640.n3 a_23668_25640.t4 6.7165
R28263 a_23668_25640.n1 a_23668_25640.t2 5.96217
R28264 a_23668_25640.n1 a_23668_25640.n0 1.33883
R28265 a_23668_25640.n4 a_23668_25640.n2 0.376152
R28266 _251_.A1.n26 _251_.A1.t31 20.9945
R28267 _251_.A1.n22 _251_.A1.t10 20.9945
R28268 _251_.A1.n12 _251_.A1.t29 20.9945
R28269 _251_.A1.n9 _251_.A1.t15 20.9945
R28270 _251_.A1.n29 _251_.A1.t12 19.4185
R28271 _251_.A1.n18 _251_.A1.t22 19.3455
R28272 _251_.A1.n17 _251_.A1.t14 18.6885
R28273 _251_.A1.n7 _251_.A1.t30 18.6885
R28274 _251_.A1.n6 _251_.A1.t18 17.5205
R28275 _251_.A1.n27 _251_.A1.t26 17.0442
R28276 _251_.A1.n23 _251_.A1.t11 17.0442
R28277 _251_.A1.n13 _251_.A1.t20 17.0442
R28278 _251_.A1.n10 _251_.A1.t23 16.9182
R28279 _251_.A1.n25 _251_.A1.t28 16.1822
R28280 _251_.A1.n21 _251_.A1.t32 16.1822
R28281 _251_.A1.n11 _251_.A1.t19 16.1822
R28282 _251_.A1.n8 _251_.A1.t16 16.1822
R28283 _251_.A1.n33 _251_.A1.t17 16.097
R28284 _251_.A1.n33 _251_.A1.t21 14.6735
R28285 _251_.A1.n25 _251_.A1.t35 14.0165
R28286 _251_.A1.n21 _251_.A1.t27 14.0165
R28287 _251_.A1.n11 _251_.A1.t33 14.0165
R28288 _251_.A1.n8 _251_.A1.t9 14.0165
R28289 _251_.A1.n7 _251_.A1.t25 11.9603
R28290 _251_.A1.n17 _251_.A1.t13 11.8873
R28291 _251_.A1.n16 _251_.A1.n15 11.7005
R28292 _251_.A1.n29 _251_.A1.t8 11.5884
R28293 _251_.A1.n18 _251_.A1.t34 11.5884
R28294 _251_.A1.n6 _251_.A1.t24 11.5588
R28295 _251_.A1.n32 _251_.A1.n16 10.8905
R28296 _251_.A1.n20 _251_.A1.n19 9.95734
R28297 _251_.A1.n20 _251_.A1 9.9005
R28298 _251_.A1.n24 _251_.A1.n23 9.0005
R28299 _251_.A1.n26 _251_.A1.n25 8.39556
R28300 _251_.A1.n22 _251_.A1.n21 8.39556
R28301 _251_.A1.n12 _251_.A1.n11 8.39556
R28302 _251_.A1.n9 _251_.A1.n8 8.39556
R28303 _251_.A1.n28 _251_.A1.n24 8.2805
R28304 _251_.A1 _251_.A1.n33 8.158
R28305 _251_.A1 _251_.A1.n6 8.05312
R28306 _251_.A1.n30 _251_.A1.n29 8.0005
R28307 _251_.A1.n19 _251_.A1.n18 8.0005
R28308 _251_.A1.n3 _251_.A1.n2 7.33746
R28309 _251_.A1.n35 _251_.A1.n34 7.3355
R28310 _251_.A1.n14 _251_.A1.n10 6.5705
R28311 _251_.A1.n34 _251_.A1.n32 6.4805
R28312 _251_.A1.n3 _251_.A1.n1 6.46093
R28313 _251_.A1.n32 _251_.A1.n31 5.9405
R28314 _251_.A1.n15 _251_.A1 5.88075
R28315 _251_.A1.n35 _251_.A1.n5 5.49618
R28316 _251_.A1.n4 _251_.A1.n0 5.4118
R28317 _251_.A1.n31 _251_.A1.n28 5.0405
R28318 _251_.A1.n16 _251_.A1 4.83558
R28319 _251_.A1.n15 _251_.A1.n14 4.7255
R28320 _251_.A1.n34 _251_.A1 4.658
R28321 _251_.A1.n31 _251_.A1.n30 4.55734
R28322 _251_.A1.n28 _251_.A1.n27 4.5005
R28323 _251_.A1.n14 _251_.A1.n13 4.5005
R28324 _251_.A1 _251_.A1.n17 4.08607
R28325 _251_.A1 _251_.A1.n7 4.08607
R28326 _251_.A1.n2 _251_.A1.t6 3.6005
R28327 _251_.A1.n2 _251_.A1.t7 3.6005
R28328 _251_.A1.n1 _251_.A1.t5 3.6005
R28329 _251_.A1.n1 _251_.A1.t4 3.6005
R28330 _251_.A1.n0 _251_.A1.t1 2.06607
R28331 _251_.A1.n5 _251_.A1.t3 2.06607
R28332 _251_.A1.n0 _251_.A1.t0 1.4923
R28333 _251_.A1.n5 _251_.A1.t2 1.4923
R28334 _251_.A1.n24 _251_.A1.n20 0.9005
R28335 _251_.A1.n4 _251_.A1.n3 0.439189
R28336 _251_.A1 _251_.A1.n35 0.3155
R28337 _251_.A1.n10 _251_.A1 0.301187
R28338 _251_.A1 _251_.A1.n4 0.203
R28339 _251_.A1.n27 _251_.A1 0.175187
R28340 _251_.A1.n23 _251_.A1 0.175187
R28341 _251_.A1.n13 _251_.A1 0.175187
R28342 _251_.A1.n30 _251_.A1 0.0498764
R28343 _251_.A1.n19 _251_.A1 0.0498764
R28344 _251_.A1 _251_.A1.n26 0.0449156
R28345 _251_.A1 _251_.A1.n22 0.0449156
R28346 _251_.A1 _251_.A1.n12 0.0449156
R28347 _251_.A1 _251_.A1.n9 0.0449156
R28348 a_20084_26023.n0 a_20084_26023.t6 121.874
R28349 a_20084_26023.t6 a_20084_26023.t3 61.5152
R28350 a_20084_26023.n1 a_20084_26023.t2 52.378
R28351 a_20084_26023.n1 a_20084_26023.t7 17.7152
R28352 a_20084_26023.n3 a_20084_26023.t1 11.1158
R28353 a_20084_26023.n4 a_20084_26023.n0 9.95623
R28354 a_20084_26023.t0 a_20084_26023.n4 8.02846
R28355 a_20084_26023.n3 a_20084_26023.n2 8.0005
R28356 a_20084_26023.n0 a_20084_26023.t5 6.7165
R28357 a_20084_26023.n2 a_20084_26023.t4 6.023
R28358 a_20084_26023.n2 a_20084_26023.n1 1.33883
R28359 a_20084_26023.n4 a_20084_26023.n3 0.376152
R28360 uo_out[1].n10 uo_out[1] 18.8871
R28361 uo_out[1].n5 uo_out[1].n4 7.21811
R28362 uo_out[1].n5 uo_out[1].n3 6.36507
R28363 uo_out[1].n6 uo_out[1].n2 6.36507
R28364 uo_out[1].n7 uo_out[1].n1 6.36507
R28365 uo_out[1].n4 uo_out[1].t4 2.89962
R28366 uo_out[1].n4 uo_out[1].t8 2.89962
R28367 uo_out[1].n3 uo_out[1].t10 2.89962
R28368 uo_out[1].n3 uo_out[1].t3 2.89962
R28369 uo_out[1].n2 uo_out[1].t2 2.89962
R28370 uo_out[1].n2 uo_out[1].t9 2.89962
R28371 uo_out[1].n1 uo_out[1].t11 2.89962
R28372 uo_out[1].n1 uo_out[1].t5 2.89962
R28373 uo_out[1].n8 uo_out[1].n0 2.70811
R28374 uo_out[1].n10 uo_out[1].n9 2.6005
R28375 uo_out[1].n9 uo_out[1].t6 2.06607
R28376 uo_out[1].n9 uo_out[1].t7 2.06607
R28377 uo_out[1].n0 uo_out[1].t1 2.06607
R28378 uo_out[1].n0 uo_out[1].t0 2.06607
R28379 uo_out[1].n8 uo_out[1].n7 1.50799
R28380 uo_out[1] uo_out[1].n10 1.21273
R28381 uo_out[1].n7 uo_out[1].n6 0.877022
R28382 uo_out[1].n6 uo_out[1].n5 0.877022
R28383 uo_out[1] uo_out[1].n8 0.267929
R28384 _335_.ZN.n14 _335_.ZN.t23 22.7157
R28385 _335_.ZN.n23 _335_.ZN.n22 19.9805
R28386 _335_.ZN.n19 _335_.ZN.t24 17.5448
R28387 _335_.ZN.n18 _335_.ZN.t22 17.5448
R28388 _335_.ZN.n15 _335_.ZN.t26 16.5107
R28389 _335_.ZN.n15 _335_.ZN.t25 14.6005
R28390 _335_.ZN.n19 _335_.ZN.n18 13.3198
R28391 _335_.ZN _335_.ZN.n15 9.14877
R28392 _335_.ZN.n22 _335_.ZN.n14 8.98846
R28393 _335_.ZN.n20 _335_.ZN.t27 8.3955
R28394 _335_.ZN.n17 _335_.ZN.t21 8.3955
R28395 _335_.ZN.n14 _335_.ZN.t20 8.3955
R28396 _335_.ZN.n4 _335_.ZN.n2 8.0692
R28397 _335_.ZN.n17 _335_.ZN.n16 8.0005
R28398 _335_.ZN.n21 _335_.ZN.n20 8.0005
R28399 _335_.ZN.n4 _335_.ZN.n3 6.3005
R28400 _335_.ZN.n23 _335_.ZN.n13 5.37335
R28401 _335_.ZN.n24 _335_.ZN.n12 5.3668
R28402 _335_.ZN.n25 _335_.ZN.n11 5.3668
R28403 _335_.ZN.n26 _335_.ZN.n10 5.3668
R28404 _335_.ZN.n27 _335_.ZN.n9 5.3668
R28405 _335_.ZN.n6 _335_.ZN.n0 5.3668
R28406 _335_.ZN.n5 _335_.ZN.n1 5.3668
R28407 _335_.ZN.n8 _335_.ZN.n7 5.3668
R28408 _335_.ZN.n20 _335_.ZN.n19 5.17133
R28409 _335_.ZN.n18 _335_.ZN.n17 5.17133
R28410 _335_.ZN.n2 _335_.ZN.t4 3.6883
R28411 _335_.ZN.n2 _335_.ZN.t7 3.6883
R28412 _335_.ZN.n3 _335_.ZN.t6 3.6883
R28413 _335_.ZN.n3 _335_.ZN.t5 3.6883
R28414 _335_.ZN.n13 _335_.ZN.t18 2.15435
R28415 _335_.ZN.n13 _335_.ZN.t8 2.15435
R28416 _335_.ZN.n12 _335_.ZN.t10 2.15435
R28417 _335_.ZN.n12 _335_.ZN.t19 2.15435
R28418 _335_.ZN.n11 _335_.ZN.t17 2.15435
R28419 _335_.ZN.n11 _335_.ZN.t11 2.15435
R28420 _335_.ZN.n10 _335_.ZN.t9 2.15435
R28421 _335_.ZN.n10 _335_.ZN.t16 2.15435
R28422 _335_.ZN.n9 _335_.ZN.t0 2.15435
R28423 _335_.ZN.n9 _335_.ZN.t14 2.15435
R28424 _335_.ZN.n0 _335_.ZN.t2 2.15435
R28425 _335_.ZN.n0 _335_.ZN.t15 2.15435
R28426 _335_.ZN.n1 _335_.ZN.t13 2.15435
R28427 _335_.ZN.n1 _335_.ZN.t1 2.15435
R28428 _335_.ZN.n7 _335_.ZN.t12 2.15435
R28429 _335_.ZN.n7 _335_.ZN.t3 2.15435
R28430 _335_.ZN.n5 _335_.ZN.n4 1.64833
R28431 _335_.ZN.n6 _335_.ZN.n5 0.812136
R28432 _335_.ZN _335_.ZN.n8 0.727045
R28433 _335_.ZN.n8 _335_.ZN.n6 0.668136
R28434 _335_.ZN.n27 _335_.ZN.n26 0.668136
R28435 _335_.ZN.n26 _335_.ZN.n25 0.668136
R28436 _335_.ZN.n25 _335_.ZN.n24 0.668136
R28437 _335_.ZN.n24 _335_.ZN.n23 0.661591
R28438 _335_.ZN.n21 _335_.ZN.n16 0.301396
R28439 _335_.ZN.n22 _335_.ZN.n21 0.0918433
R28440 _335_.ZN _335_.ZN.n27 0.0855909
R28441 _335_.ZN.n16 _335_.ZN 0.0596045
R28442 _381_.A2.n4 _381_.A2 23.6755
R28443 _381_.A2.n0 _381_.A2.t4 19.5645
R28444 _381_.A2.n0 _381_.A2.t7 17.1312
R28445 _381_.A2.n1 _381_.A2.t2 16.3525
R28446 _381_.A2.n2 _381_.A2.t5 15.5008
R28447 _381_.A2.n2 _381_.A2.t6 14.7222
R28448 _381_.A2.n1 _381_.A2.t3 13.8705
R28449 _381_.A2.n5 _381_.A2.n4 13.7035
R28450 _381_.A2 _381_.A2.n2 9.51081
R28451 _381_.A2.n4 _381_.A2.n3 9.0005
R28452 _381_.A2.n3 _381_.A2.n1 8.59522
R28453 _381_.A2.n5 _381_.A2.t1 8.30853
R28454 _381_.A2 _381_.A2.n0 8.1405
R28455 _381_.A2 _381_.A2.t0 4.1573
R28456 _381_.A2 _381_.A2.n5 0.374266
R28457 _381_.A2.n3 _381_.A2 0.296971
R28458 _352_.A2.n18 _352_.A2.t20 27.8865
R28459 _352_.A2.n14 _352_.A2.t22 20.5135
R28460 _352_.A2.n21 _352_.A2.t30 19.4185
R28461 _352_.A2.n13 _352_.A2.t28 18.5425
R28462 _352_.A2.n25 _352_.A2.t21 16.3282
R28463 _352_.A2.n19 _352_.A2.t31 16.3282
R28464 _352_.A2.n9 _352_.A2.t24 15.7685
R28465 _352_.A2.n11 _352_.A2.t26 15.3305
R28466 _352_.A2.n11 _352_.A2.t29 15.148
R28467 _352_.A2.n25 _352_.A2.t18 14.7465
R28468 _352_.A2.n19 _352_.A2.t19 14.6735
R28469 _352_.A2.n9 _352_.A2.t27 14.637
R28470 _352_.A2.n13 _352_.A2.t16 14.053
R28471 _352_.A2.n16 _352_.A2.n12 13.5131
R28472 _352_.A2.n21 _352_.A2.t17 11.5884
R28473 _352_.A2.n14 _352_.A2.t25 11.4372
R28474 _352_.A2.n23 _352_.A2 11.4305
R28475 _352_.A2.n17 _352_.A2.n10 10.7298
R28476 _352_.A2.n16 _352_.A2.n15 9.8105
R28477 _352_.A2 _352_.A2.n14 8.96449
R28478 _352_.A2.n15 _352_.A2.n13 8.7076
R28479 _352_.A2.n22 _352_.A2 8.4155
R28480 _352_.A2 _352_.A2.n18 8.09214
R28481 _352_.A2 _352_.A2.n21 8.04988
R28482 _352_.A2 _352_.A2.n25 8.0005
R28483 _352_.A2.n20 _352_.A2.n19 8.0005
R28484 _352_.A2.n12 _352_.A2.n11 8.0005
R28485 _352_.A2.n10 _352_.A2.n9 8.0005
R28486 _352_.A2.n7 _352_.A2.n5 7.85007
R28487 _352_.A2.n29 _352_.A2.n8 6.40811
R28488 _352_.A2.n7 _352_.A2.n6 6.3005
R28489 _352_.A2.n24 _352_.A2.n23 6.3005
R28490 _352_.A2.n28 _352_.A2.n27 6.3005
R28491 _352_.A2.n24 _352_.A2.n17 6.1205
R28492 _352_.A2.n18 _352_.A2.t23 5.8405
R28493 _352_.A2.n2 _352_.A2.n0 5.67738
R28494 _352_.A2.n28 _352_.A2.n26 5.5715
R28495 _352_.A2.n4 _352_.A2.n3 5.2005
R28496 _352_.A2.n32 _352_.A2.n31 5.2005
R28497 _352_.A2.n2 _352_.A2.n1 5.2005
R28498 _352_.A2.n22 _352_.A2.n20 4.62366
R28499 _352_.A2.n23 _352_.A2.n22 4.5005
R28500 _352_.A2.n26 _352_.A2 4.5005
R28501 _352_.A2.n27 _352_.A2.t4 3.21226
R28502 _352_.A2.n27 _352_.A2.t7 3.21226
R28503 _352_.A2.n8 _352_.A2.t5 3.21226
R28504 _352_.A2.n8 _352_.A2.t6 3.21226
R28505 _352_.A2.n6 _352_.A2.t12 1.99806
R28506 _352_.A2.n6 _352_.A2.t15 1.99806
R28507 _352_.A2.n5 _352_.A2.t14 1.99806
R28508 _352_.A2.n5 _352_.A2.t13 1.99806
R28509 _352_.A2.n17 _352_.A2.n16 1.9805
R28510 _352_.A2.n31 _352_.A2.t8 1.51717
R28511 _352_.A2.n31 _352_.A2.t1 1.51717
R28512 _352_.A2.n3 _352_.A2.t2 1.51717
R28513 _352_.A2.n3 _352_.A2.t10 1.51717
R28514 _352_.A2.n0 _352_.A2.t3 1.51717
R28515 _352_.A2.n0 _352_.A2.t9 1.51717
R28516 _352_.A2.n1 _352_.A2.t11 1.51717
R28517 _352_.A2.n1 _352_.A2.t0 1.51717
R28518 _352_.A2.n26 _352_.A2.n24 1.2605
R28519 _352_.A2.n30 _352_.A2.n7 0.930189
R28520 _352_.A2.n29 _352_.A2.n28 0.741246
R28521 _352_.A2.n32 _352_.A2.n30 0.494593
R28522 _352_.A2.n4 _352_.A2.n2 0.477383
R28523 _352_.A2 _352_.A2.n4 0.444656
R28524 _352_.A2.n15 _352_.A2 0.373833
R28525 _352_.A2.n30 _352_.A2.n29 0.284786
R28526 _352_.A2.n12 _352_.A2 0.190411
R28527 _352_.A2.n10 _352_.A2 0.125214
R28528 _352_.A2 _352_.A2.n32 0.0332273
R28529 _352_.A2.n20 _352_.A2 0.00997368
R28530 _459_.Q.n17 _459_.Q.n10 22.6805
R28531 _459_.Q.n15 _459_.Q.t7 19.7105
R28532 _459_.Q.n7 _459_.Q.t17 19.0535
R28533 _459_.Q.n6 _459_.Q.t15 19.0535
R28534 _459_.Q.n1 _459_.Q.t3 19.0535
R28535 _459_.Q.n2 _459_.Q.t12 19.0535
R28536 _459_.Q.n11 _459_.Q.t10 18.6885
R28537 _459_.Q.n12 _459_.Q.t11 18.6885
R28538 _459_.Q.n14 _459_.Q.t4 17.8003
R28539 _459_.Q.n7 _459_.Q.n6 16.5048
R28540 _459_.Q.n2 _459_.Q.n1 16.5048
R28541 _459_.Q.n14 _459_.Q.t6 14.7465
R28542 _459_.Q.n15 _459_.Q.t2 14.3085
R28543 _459_.Q.n16 _459_.Q 14.2205
R28544 _459_.Q.n17 _459_.Q.n16 13.3205
R28545 _459_.Q.n12 _459_.Q.t5 11.9603
R28546 _459_.Q.n11 _459_.Q.t16 11.8752
R28547 _459_.Q.n13 _459_.Q 10.5607
R28548 _459_.Q.n8 _459_.Q.t9 8.73617
R28549 _459_.Q.n5 _459_.Q.t13 8.73617
R28550 _459_.Q.n0 _459_.Q.t14 8.73617
R28551 _459_.Q.n3 _459_.Q.t8 8.73617
R28552 _459_.Q _459_.Q.t1 8.69622
R28553 _459_.Q.n4 _459_.Q.n0 8.39376
R28554 _459_.Q.n9 _459_.Q.n5 8.3918
R28555 _459_.Q _459_.Q.n14 8.11418
R28556 _459_.Q _459_.Q.n11 8.06425
R28557 _459_.Q _459_.Q.n15 8.00997
R28558 _459_.Q.n9 _459_.Q.n8 8.0005
R28559 _459_.Q.n4 _459_.Q.n3 8.0005
R28560 _459_.Q _459_.Q.t0 6.72245
R28561 _459_.Q.n8 _459_.Q.n7 6.0595
R28562 _459_.Q.n6 _459_.Q.n5 6.0595
R28563 _459_.Q.n1 _459_.Q.n0 6.0595
R28564 _459_.Q.n3 _459_.Q.n2 6.0595
R28565 _459_.Q _459_.Q.n17 5.5805
R28566 _459_.Q.n13 _459_.Q 4.6405
R28567 _459_.Q.n16 _459_.Q 4.63313
R28568 _459_.Q _459_.Q.n12 4.08607
R28569 _459_.Q.n16 _459_.Q.n13 1.5755
R28570 _459_.Q _459_.Q.n4 0.520283
R28571 _459_.Q.n10 _459_.Q.n9 0.251587
R28572 _459_.Q.n10 _459_.Q 0.146587
R28573 _452_.Q.n1 _452_.Q.t14 29.2005
R28574 _452_.Q.n13 _452_.Q 26.6405
R28575 _452_.Q.n10 _452_.Q.t6 20.3675
R28576 _452_.Q.n17 _452_.Q.t11 19.7105
R28577 _452_.Q.n0 _452_.Q.t18 19.4915
R28578 _452_.Q.n15 _452_.Q.t19 17.8003
R28579 _452_.Q.n11 _452_.Q.t12 16.2795
R28580 _452_.Q.n3 _452_.Q.t10 15.5738
R28581 _452_.Q.n8 _452_.Q.t9 15.3305
R28582 _452_.Q.n11 _452_.Q.t17 15.2818
R28583 _452_.Q.n8 _452_.Q.t13 15.0872
R28584 _452_.Q.n4 _452_.Q.t20 14.8317
R28585 _452_.Q.n15 _452_.Q.t15 14.8195
R28586 _452_.Q.n17 _452_.Q.t21 14.3085
R28587 _452_.Q.n4 _452_.Q.t5 13.9435
R28588 _452_.Q.n0 _452_.Q.t4 13.6758
R28589 _452_.Q.n10 _452_.Q.t8 13.3352
R28590 _452_.Q.n3 _452_.Q.t16 13.2013
R28591 _452_.Q.n1 _452_.Q.t7 12.1428
R28592 _452_.Q.n16 _452_.Q.n14 10.2605
R28593 _452_.Q.n9 _452_.Q 9.50873
R28594 _452_.Q _452_.Q.n8 8.19041
R28595 _452_.Q _452_.Q.n15 8.11418
R28596 _452_.Q.n2 _452_.Q.n1 8.07925
R28597 _452_.Q _452_.Q.n10 8.05321
R28598 _452_.Q _452_.Q.n0 8.03988
R28599 _452_.Q.n12 _452_.Q.n11 8.02829
R28600 _452_.Q _452_.Q.n3 8.01992
R28601 _452_.Q.n5 _452_.Q.n4 8.0005
R28602 _452_.Q _452_.Q.n17 8.0005
R28603 _452_.Q.n7 _452_.Q 7.898
R28604 _452_.Q _452_.Q.n21 6.75428
R28605 _452_.Q.n6 _452_.Q.n5 6.65127
R28606 _452_.Q.n14 _452_.Q.n13 6.4805
R28607 _452_.Q.n18 _452_.Q 6.413
R28608 _452_.Q.n9 _452_.Q.n7 5.9405
R28609 _452_.Q.n20 _452_.Q.n19 5.2005
R28610 _452_.Q.n6 _452_.Q.n2 4.9955
R28611 _452_.Q.n20 _452_.Q.n18 4.51445
R28612 _452_.Q.n13 _452_.Q.n12 4.5005
R28613 _452_.Q.n16 _452_.Q 4.5005
R28614 _452_.Q.n18 _452_.Q.n16 2.6555
R28615 _452_.Q.n21 _452_.Q.t2 1.99806
R28616 _452_.Q.n21 _452_.Q.t3 1.99806
R28617 _452_.Q.n19 _452_.Q.t0 1.4923
R28618 _452_.Q.n19 _452_.Q.t1 1.4923
R28619 _452_.Q.n5 _452_.Q 1.01483
R28620 _452_.Q.n14 _452_.Q.n9 0.5405
R28621 _452_.Q.n12 _452_.Q 0.148735
R28622 _452_.Q.n7 _452_.Q.n6 0.1355
R28623 _452_.Q.n2 _452_.Q 0.1265
R28624 _452_.Q _452_.Q.n20 0.064686
R28625 a_49152_30301.n3 a_49152_30301.t2 121.874
R28626 a_49152_30301.t2 a_49152_30301.t3 61.5152
R28627 a_49152_30301.n0 a_49152_30301.t6 52.378
R28628 a_49152_30301.n0 a_49152_30301.t7 17.7882
R28629 a_49152_30301.n2 a_49152_30301.t1 11.1158
R28630 a_49152_30301.n4 a_49152_30301.n3 9.95623
R28631 a_49152_30301.t0 a_49152_30301.n4 8.02846
R28632 a_49152_30301.n2 a_49152_30301.n1 8.0005
R28633 a_49152_30301.n3 a_49152_30301.t5 6.7165
R28634 a_49152_30301.n1 a_49152_30301.t4 5.96217
R28635 a_49152_30301.n1 a_49152_30301.n0 1.33883
R28636 a_49152_30301.n4 a_49152_30301.n2 0.376152
R28637 a_36996_18183.n0 a_36996_18183.t4 121.874
R28638 a_36996_18183.t4 a_36996_18183.t3 61.5152
R28639 a_36996_18183.n1 a_36996_18183.t2 52.378
R28640 a_36996_18183.n1 a_36996_18183.t7 17.7152
R28641 a_36996_18183.n3 a_36996_18183.t1 11.1158
R28642 a_36996_18183.n4 a_36996_18183.n0 9.95623
R28643 a_36996_18183.t0 a_36996_18183.n4 8.02846
R28644 a_36996_18183.n3 a_36996_18183.n2 8.0005
R28645 a_36996_18183.n0 a_36996_18183.t5 6.7165
R28646 a_36996_18183.n2 a_36996_18183.t6 6.023
R28647 a_36996_18183.n2 a_36996_18183.n1 1.33883
R28648 a_36996_18183.n4 a_36996_18183.n3 0.376152
R28649 a_42392_22825.n11 a_42392_22825.t22 15.4765
R28650 a_42392_22825.n12 a_42392_22825.t28 15.4765
R28651 a_42392_22825.n13 a_42392_22825.t23 15.4765
R28652 a_42392_22825.n14 a_42392_22825.t24 15.4765
R28653 a_42392_22825.n15 a_42392_22825.t41 15.4765
R28654 a_42392_22825.n16 a_42392_22825.t38 15.4765
R28655 a_42392_22825.n17 a_42392_22825.t42 15.4765
R28656 a_42392_22825.n18 a_42392_22825.t39 15.4765
R28657 a_42392_22825.n19 a_42392_22825.t15 15.4765
R28658 a_42392_22825.n20 a_42392_22825.t19 15.4765
R28659 a_42392_22825.n21 a_42392_22825.t16 15.4765
R28660 a_42392_22825.n24 a_42392_22825.t20 15.4765
R28661 a_42392_22825.n8 a_42392_22825.t32 15.4765
R28662 a_42392_22825.n9 a_42392_22825.t34 15.4765
R28663 a_42392_22825.n10 a_42392_22825.t30 15.4765
R28664 a_42392_22825.n25 a_42392_22825.t25 15.4765
R28665 a_42392_22825.n11 a_42392_22825.t17 11.863
R28666 a_42392_22825.n12 a_42392_22825.t33 11.863
R28667 a_42392_22825.n13 a_42392_22825.t29 11.863
R28668 a_42392_22825.n14 a_42392_22825.t31 11.863
R28669 a_42392_22825.n15 a_42392_22825.t35 11.863
R28670 a_42392_22825.n16 a_42392_22825.t43 11.863
R28671 a_42392_22825.n17 a_42392_22825.t14 11.863
R28672 a_42392_22825.n18 a_42392_22825.t44 11.863
R28673 a_42392_22825.n19 a_42392_22825.t45 11.863
R28674 a_42392_22825.n20 a_42392_22825.t26 11.863
R28675 a_42392_22825.n8 a_42392_22825.t37 11.863
R28676 a_42392_22825.n9 a_42392_22825.t40 11.863
R28677 a_42392_22825.n10 a_42392_22825.t36 11.863
R28678 a_42392_22825.n25 a_42392_22825.t18 11.863
R28679 a_42392_22825.n22 a_42392_22825.t21 11.8022
R28680 a_42392_22825.n23 a_42392_22825.t27 11.8022
R28681 a_42392_22825.n5 a_42392_22825.t9 11.3584
R28682 a_42392_22825.n12 a_42392_22825.n11 10.5449
R28683 a_42392_22825.n13 a_42392_22825.n12 10.5449
R28684 a_42392_22825.n14 a_42392_22825.n13 10.5449
R28685 a_42392_22825.n15 a_42392_22825.n14 10.5449
R28686 a_42392_22825.n16 a_42392_22825.n15 10.5449
R28687 a_42392_22825.n17 a_42392_22825.n16 10.5449
R28688 a_42392_22825.n18 a_42392_22825.n17 10.5449
R28689 a_42392_22825.n19 a_42392_22825.n18 10.5449
R28690 a_42392_22825.n20 a_42392_22825.n19 10.5449
R28691 a_42392_22825.n21 a_42392_22825.n20 10.5449
R28692 a_42392_22825.n9 a_42392_22825.n8 10.5449
R28693 a_42392_22825.n10 a_42392_22825.n9 10.5449
R28694 a_42392_22825.n25 a_42392_22825.n10 10.5449
R28695 a_42392_22825.n25 a_42392_22825.n24 10.5449
R28696 a_42392_22825.n7 a_42392_22825.t12 10.4819
R28697 a_42392_22825.n23 a_42392_22825.n22 10.26
R28698 a_42392_22825.n6 a_42392_22825.n3 6.43746
R28699 a_42392_22825.n5 a_42392_22825.n4 6.43746
R28700 a_42392_22825.n29 a_42392_22825.n0 6.25311
R28701 a_42392_22825.n28 a_42392_22825.n1 5.37659
R28702 a_42392_22825.n27 a_42392_22825.n2 5.37659
R28703 a_42392_22825.n30 a_42392_22825.n29 5.37659
R28704 a_42392_22825.n3 a_42392_22825.t11 4.04494
R28705 a_42392_22825.n3 a_42392_22825.t13 4.04494
R28706 a_42392_22825.n4 a_42392_22825.t10 4.04494
R28707 a_42392_22825.n4 a_42392_22825.t8 4.04494
R28708 a_42392_22825.n0 a_42392_22825.t5 3.07367
R28709 a_42392_22825.n1 a_42392_22825.t1 3.07367
R28710 a_42392_22825.n2 a_42392_22825.t2 3.07367
R28711 a_42392_22825.n30 a_42392_22825.t4 3.07367
R28712 a_42392_22825.n0 a_42392_22825.t3 2.22001
R28713 a_42392_22825.n1 a_42392_22825.t6 2.22001
R28714 a_42392_22825.n2 a_42392_22825.t0 2.22001
R28715 a_42392_22825.t7 a_42392_22825.n30 2.22001
R28716 a_42392_22825.n26 a_42392_22825.n25 1.9195
R28717 a_42392_22825.n6 a_42392_22825.n5 0.877022
R28718 a_42392_22825.n7 a_42392_22825.n6 0.877022
R28719 a_42392_22825.n29 a_42392_22825.n28 0.877022
R28720 a_42392_22825.n28 a_42392_22825.n27 0.877022
R28721 a_42392_22825.n27 a_42392_22825.n26 0.430935
R28722 a_42392_22825.n26 a_42392_22825.n7 0.313543
R28723 a_42392_22825.n22 a_42392_22825.n21 0.0613333
R28724 a_42392_22825.n24 a_42392_22825.n23 0.0613333
R28725 a_17060_28776.n3 a_17060_28776.t5 121.874
R28726 a_17060_28776.t5 a_17060_28776.t3 61.5152
R28727 a_17060_28776.n0 a_17060_28776.t2 52.378
R28728 a_17060_28776.n0 a_17060_28776.t4 17.7882
R28729 a_17060_28776.n2 a_17060_28776.t1 11.1158
R28730 a_17060_28776.n4 a_17060_28776.n3 9.99927
R28731 a_17060_28776.n2 a_17060_28776.n1 8.0005
R28732 a_17060_28776.n3 a_17060_28776.t7 6.7165
R28733 a_17060_28776.n1 a_17060_28776.t6 5.96217
R28734 a_17060_28776.t0 a_17060_28776.n4 5.40498
R28735 a_17060_28776.n1 a_17060_28776.n0 1.33883
R28736 a_17060_28776.n4 a_17060_28776.n2 0.333109
R28737 uio_out[6].n2 uio_out[6].t8 20.4405
R28738 uio_out[6].n3 uio_out[6].t11 17.7395
R28739 uio_out[6].n2 uio_out[6].t9 15.3305
R28740 uio_out[6].n3 uio_out[6].t10 12.6782
R28741 uio_out[6].n5 uio_out[6] 12.3826
R28742 uio_out[6].n6 uio_out[6].n5 11.8237
R28743 uio_out[6] uio_out[6].n2 8.06925
R28744 uio_out[6].n9 uio_out[6].n1 7.02935
R28745 uio_out[6].n8 uio_out[6].n7 6.3005
R28746 uio_out[6].n8 uio_out[6].n6 6.1853
R28747 uio_out[6] uio_out[6].n11 5.3505
R28748 uio_out[6].n10 uio_out[6].n0 5.2005
R28749 uio_out[6].n6 uio_out[6] 4.6405
R28750 uio_out[6].n5 uio_out[6].n4 4.56214
R28751 uio_out[6].n4 uio_out[6].n3 4.0005
R28752 uio_out[6].n11 uio_out[6].t3 2.06607
R28753 uio_out[6].n11 uio_out[6].t1 2.06607
R28754 uio_out[6].n0 uio_out[6].t2 2.06607
R28755 uio_out[6].n0 uio_out[6].t0 2.06607
R28756 uio_out[6].n7 uio_out[6].t5 2.01032
R28757 uio_out[6].n7 uio_out[6].t4 2.01032
R28758 uio_out[6].n1 uio_out[6].t7 2.01032
R28759 uio_out[6].n1 uio_out[6].t6 2.01032
R28760 uio_out[6].n10 uio_out[6].n9 0.304937
R28761 uio_out[6] uio_out[6].n10 0.1865
R28762 uio_out[6].n4 uio_out[6] 0.0769384
R28763 uio_out[6].n9 uio_out[6].n8 0.0104
R28764 uio_out[7].n6 uio_out[7].t10 22.1195
R28765 uio_out[7].n5 uio_out[7].t9 19.5645
R28766 uio_out[7].n5 uio_out[7].t8 18.4938
R28767 uio_out[7].n7 uio_out[7] 13.9576
R28768 uio_out[7].n6 uio_out[7].t11 9.02817
R28769 uio_out[7].n9 uio_out[7].n7 8.7935
R28770 uio_out[7] uio_out[7].n5 8.51318
R28771 uio_out[7] uio_out[7].n6 8.35407
R28772 uio_out[7].n2 uio_out[7].n0 7.06159
R28773 uio_out[7].n2 uio_out[7].n1 6.31353
R28774 uio_out[7].n4 uio_out[7].n3 5.2005
R28775 uio_out[7].n9 uio_out[7].n8 5.2005
R28776 uio_out[7].n7 uio_out[7] 4.5005
R28777 uio_out[7].n8 uio_out[7].t3 2.06607
R28778 uio_out[7].n8 uio_out[7].t0 2.06607
R28779 uio_out[7].n3 uio_out[7].t2 2.06607
R28780 uio_out[7].n3 uio_out[7].t1 2.06607
R28781 uio_out[7].n1 uio_out[7].t7 2.01032
R28782 uio_out[7].n1 uio_out[7].t5 2.01032
R28783 uio_out[7].n0 uio_out[7].t6 2.01032
R28784 uio_out[7].n0 uio_out[7].t4 2.01032
R28785 uio_out[7].n4 uio_out[7].n2 0.314316
R28786 uio_out[7] uio_out[7].n4 0.1865
R28787 uio_out[7] uio_out[7].n9 0.1505
R28788 uio_out[5].n5 uio_out[5].t13 19.8565
R28789 uio_out[5].n9 uio_out[5].t8 18.9805
R28790 uio_out[5].n7 uio_out[5].t11 18.6885
R28791 uio_out[5].n5 uio_out[5].t12 15.9145
R28792 uio_out[5].n7 uio_out[5].t9 11.9603
R28793 uio_out[5].n8 uio_out[5].n6 11.903
R28794 uio_out[5].n9 uio_out[5].t10 11.4372
R28795 uio_out[5].n13 uio_out[5].n11 10.8185
R28796 uio_out[5].n8 uio_out[5] 9.16575
R28797 uio_out[5].n10 uio_out[5] 9.13858
R28798 uio_out[5] uio_out[5].n9 8.11576
R28799 uio_out[5].n6 uio_out[5].n5 8.0005
R28800 uio_out[5].n2 uio_out[5].n0 7.06159
R28801 uio_out[5].n11 uio_out[5] 6.44257
R28802 uio_out[5].n2 uio_out[5].n1 6.31353
R28803 uio_out[5].n4 uio_out[5].n3 5.2005
R28804 uio_out[5].n13 uio_out[5].n12 5.2005
R28805 uio_out[5] uio_out[5].n7 4.08607
R28806 uio_out[5].n12 uio_out[5].t3 2.06607
R28807 uio_out[5].n12 uio_out[5].t1 2.06607
R28808 uio_out[5].n3 uio_out[5].t2 2.06607
R28809 uio_out[5].n3 uio_out[5].t0 2.06607
R28810 uio_out[5].n1 uio_out[5].t5 2.01032
R28811 uio_out[5].n1 uio_out[5].t6 2.01032
R28812 uio_out[5].n0 uio_out[5].t4 2.01032
R28813 uio_out[5].n0 uio_out[5].t7 2.01032
R28814 uio_out[5].n10 uio_out[5].n8 1.0805
R28815 uio_out[5].n11 uio_out[5].n10 0.3605
R28816 uio_out[5].n4 uio_out[5].n2 0.314316
R28817 uio_out[5] uio_out[5].n4 0.1865
R28818 uio_out[5] uio_out[5].n13 0.1505
R28819 uio_out[5].n6 uio_out[5] 0.053
R28820 _448_.Q.n5 _448_.Q.t11 24.9665
R28821 _448_.Q.n4 _448_.Q 23.1755
R28822 _448_.Q.n11 _448_.Q.t3 19.1995
R28823 _448_.Q.n0 _448_.Q.t5 18.6885
R28824 _448_.Q.n2 _448_.Q.t8 17.7395
R28825 _448_.Q.n1 _448_.Q.t9 17.5692
R28826 _448_.Q.n9 _448_.Q.t6 17.5205
R28827 _448_.Q.n3 _448_.Q.t14 16.3768
R28828 _448_.Q.n1 _448_.Q.t4 16.1335
R28829 _448_.Q.n3 _448_.Q.t12 14.7222
R28830 _448_.Q.n11 _448_.Q.t13 13.6637
R28831 _448_.Q.n2 _448_.Q.t7 12.6782
R28832 _448_.Q.n0 _448_.Q.t2 11.9603
R28833 _448_.Q.n9 _448_.Q.t15 11.5588
R28834 _448_.Q.n7 _448_.Q.n6 9.85815
R28835 _448_.Q.n5 _448_.Q.t10 8.73617
R28836 _448_.Q _448_.Q.t1 8.69622
R28837 _448_.Q _448_.Q.n9 8.05312
R28838 _448_.Q _448_.Q.n1 8.0265
R28839 _448_.Q _448_.Q.n3 8.02581
R28840 _448_.Q _448_.Q.n11 8.0005
R28841 _448_.Q.n6 _448_.Q.n5 8.0005
R28842 _448_.Q.n8 _448_.Q.n7 7.1105
R28843 _448_.Q _448_.Q.t0 6.72245
R28844 _448_.Q.n8 _448_.Q 6.4405
R28845 _448_.Q.n7 _448_.Q.n4 6.3005
R28846 _448_.Q _448_.Q.n13 6.1655
R28847 _448_.Q.n13 _448_.Q 5.4455
R28848 _448_.Q.n12 _448_.Q 4.8205
R28849 _448_.Q.n10 _448_.Q 4.65558
R28850 _448_.Q.n4 _448_.Q 4.5005
R28851 _448_.Q _448_.Q.n0 4.08607
R28852 _448_.Q _448_.Q.n2 4.07694
R28853 _448_.Q.n12 _448_.Q.n10 2.3855
R28854 _448_.Q.n10 _448_.Q.n8 0.3605
R28855 _448_.Q.n13 _448_.Q.n12 0.1805
R28856 _448_.Q.n6 _448_.Q 0.0110882
R28857 _229_.I.n1 _229_.I.t10 20.2945
R28858 _229_.I.n9 _229_.I.t6 19.8565
R28859 _229_.I.n7 _229_.I.t13 18.9805
R28860 _229_.I.n6 _229_.I.t3 17.5205
R28861 _229_.I.n4 _229_.I.t5 16.3403
R28862 _229_.I.n2 _229_.I.t8 16.3282
R28863 _229_.I.n9 _229_.I.t11 15.9875
R28864 _229_.I.n0 _229_.I.t2 15.659
R28865 _229_.I.n2 _229_.I.t9 15.6225
R28866 _229_.I.n4 _229_.I.t4 14.7465
R28867 _229_.I.n0 _229_.I.t14 14.6735
R28868 _229_.I.n1 _229_.I.t7 12.301
R28869 _229_.I.n6 _229_.I.t15 11.5588
R28870 _229_.I.n7 _229_.I.t12 11.4372
R28871 _229_.I.n11 _229_.I.n10 11.408
R28872 _229_.I.n15 _229_.I.n14 11.1605
R28873 _229_.I.n8 _229_.I 10.4405
R28874 _229_.I.n12 _229_.I.n5 9.7205
R28875 _229_.I.n14 _229_.I 9.64978
R28876 _229_.I.n8 _229_.I 9.1805
R28877 _229_.I _229_.I.n2 8.4405
R28878 _229_.I.n15 _229_.I.t1 8.30886
R28879 _229_.I.n3 _229_.I.n1 8.17606
R28880 _229_.I _229_.I.n7 8.11457
R28881 _229_.I _229_.I.n6 8.05312
R28882 _229_.I _229_.I.n0 8.00596
R28883 _229_.I.n5 _229_.I.n4 8.0005
R28884 _229_.I.n10 _229_.I.n9 8.0005
R28885 _229_.I.n13 _229_.I.n12 5.7605
R28886 _229_.I.n14 _229_.I.n13 4.8605
R28887 _229_.I.n13 _229_.I.n3 4.5005
R28888 _229_.I _229_.I.t0 4.3844
R28889 _229_.I.n11 _229_.I.n8 2.8805
R28890 _229_.I.n12 _229_.I.n11 1.4405
R28891 _229_.I.n3 _229_.I 0.187167
R28892 _229_.I.n5 _229_.I 0.128095
R28893 _229_.I _229_.I.n15 0.08114
R28894 _229_.I.n10 _229_.I 0.053
R28895 a_27588_29159.n0 a_27588_29159.t4 121.874
R28896 a_27588_29159.t4 a_27588_29159.t2 61.5152
R28897 a_27588_29159.n1 a_27588_29159.t7 52.378
R28898 a_27588_29159.n1 a_27588_29159.t6 17.7152
R28899 a_27588_29159.n3 a_27588_29159.t1 11.1158
R28900 a_27588_29159.n4 a_27588_29159.n0 9.95623
R28901 a_27588_29159.t0 a_27588_29159.n4 8.02846
R28902 a_27588_29159.n3 a_27588_29159.n2 8.0005
R28903 a_27588_29159.n0 a_27588_29159.t5 6.7165
R28904 a_27588_29159.n2 a_27588_29159.t3 6.023
R28905 a_27588_29159.n2 a_27588_29159.n1 1.33883
R28906 a_27588_29159.n4 a_27588_29159.n3 0.376152
R28907 _437_.A1.n1 _437_.A1.t10 19.5645
R28908 _437_.A1.n5 _437_.A1.t4 19.1995
R28909 _437_.A1.n14 _437_.A1.t11 18.6885
R28910 _437_.A1.n3 _437_.A1.t14 18.6885
R28911 _437_.A1.n10 _437_.A1.t9 18.6885
R28912 _437_.A1.n1 _437_.A1.t15 18.4938
R28913 _437_.A1.n0 _437_.A1.t2 16.7662
R28914 _437_.A1.n7 _437_.A1.t12 16.2795
R28915 _437_.A1.n7 _437_.A1.t13 15.2818
R28916 _437_.A1.n0 _437_.A1.t5 14.3815
R28917 _437_.A1.n5 _437_.A1.t7 13.6637
R28918 _437_.A1.n16 _437_.A1.n15 12.0605
R28919 _437_.A1.n3 _437_.A1.t6 11.9603
R28920 _437_.A1.n10 _437_.A1.t3 11.9603
R28921 _437_.A1.n14 _437_.A1.t8 11.8873
R28922 _437_.A1.n12 _437_.A1.n11 11.6493
R28923 _437_.A1 _437_.A1.t1 8.69622
R28924 _437_.A1 _437_.A1.n1 8.16594
R28925 _437_.A1.n8 _437_.A1.n7 8.02829
R28926 _437_.A1.n2 _437_.A1.n0 8.01064
R28927 _437_.A1.n6 _437_.A1.n5 8.0005
R28928 _437_.A1.n13 _437_.A1.n12 7.6955
R28929 _437_.A1.n9 _437_.A1.n6 7.1555
R28930 _437_.A1 _437_.A1.t0 6.72245
R28931 _437_.A1.n12 _437_.A1.n9 6.4805
R28932 _437_.A1.n16 _437_.A1.n2 5.5805
R28933 _437_.A1.n13 _437_.A1.n4 5.26107
R28934 _437_.A1.n9 _437_.A1.n8 4.8155
R28935 _437_.A1.n15 _437_.A1 4.5005
R28936 _437_.A1 _437_.A1.n16 4.5005
R28937 _437_.A1 _437_.A1.n14 4.08607
R28938 _437_.A1.n4 _437_.A1.n3 4.0005
R28939 _437_.A1.n11 _437_.A1.n10 4.0005
R28940 _437_.A1.n15 _437_.A1.n13 1.9355
R28941 _437_.A1.n2 _437_.A1 1.18617
R28942 _437_.A1.n4 _437_.A1 0.245418
R28943 _437_.A1.n8 _437_.A1 0.148735
R28944 _437_.A1.n6 _437_.A1 0.1405
R28945 _437_.A1.n11 _437_.A1 0.0860738
R28946 _455_.Q.n11 _455_.Q.t11 17.484
R28947 _455_.Q.n7 _455_.Q.t14 17.2772
R28948 _455_.Q.n7 _455_.Q.t4 16.5715
R28949 _455_.Q.n2 _455_.Q.t3 16.5715
R28950 _455_.Q.n5 _455_.Q.t8 16.5715
R28951 _455_.Q.n0 _455_.Q.t6 16.5715
R28952 _455_.Q.n4 _455_.Q.n3 16.5048
R28953 _455_.Q.n9 _455_.Q.t12 16.3282
R28954 _455_.Q.n12 _455_.Q.t2 16.3282
R28955 _455_.Q.n0 _455_.Q.t5 15.6468
R28956 _455_.Q.n3 _455_.Q.t9 14.7952
R28957 _455_.Q.n4 _455_.Q.t7 14.7952
R28958 _455_.Q.n12 _455_.Q.t15 14.7465
R28959 _455_.Q.n9 _455_.Q.t10 14.6735
R28960 _455_.Q.n10 _455_.Q.n8 12.6905
R28961 _455_.Q.n11 _455_.Q.t13 11.863
R28962 _455_.Q.n14 _455_.Q 10.5909
R28963 _455_.Q.n14 _455_.Q.n13 9.09844
R28964 _455_.Q.n15 _455_.Q.n10 9.0905
R28965 _455_.Q.n10 _455_.Q 9.0005
R28966 _455_.Q _455_.Q.t1 8.69622
R28967 _455_.Q _455_.Q.n9 8.13668
R28968 _455_.Q.n13 _455_.Q.n12 8.13432
R28969 _455_.Q _455_.Q.n0 8.11638
R28970 _455_.Q _455_.Q.n11 8.08781
R28971 _455_.Q.n8 _455_.Q.n7 8.05865
R28972 _455_.Q.n6 _455_.Q.n5 8.0005
R28973 _455_.Q.n2 _455_.Q.n1 8.0005
R28974 _455_.Q.n15 _455_.Q.n14 6.8405
R28975 _455_.Q _455_.Q.t0 6.72245
R28976 _455_.Q _455_.Q.n15 5.7605
R28977 _455_.Q.n3 _455_.Q.n2 2.4825
R28978 _455_.Q.n5 _455_.Q.n4 2.4825
R28979 _455_.Q.n8 _455_.Q.n6 1.20982
R28980 _455_.Q.n1 _455_.Q 1.08463
R28981 _455_.Q.n6 _455_.Q.n1 0.39425
R28982 _455_.Q.n13 _455_.Q 0.00286842
R28983 uo_out[5].n9 uo_out[5] 15.2626
R28984 uo_out[5].n6 uo_out[5].n5 7.21811
R28985 uo_out[5].n8 uo_out[5].n2 6.36507
R28986 uo_out[5].n7 uo_out[5].n3 6.36507
R28987 uo_out[5].n6 uo_out[5].n4 6.36507
R28988 uo_out[5] uo_out[5].n0 3.81667
R28989 uo_out[5].n2 uo_out[5].t9 2.89962
R28990 uo_out[5].n2 uo_out[5].t3 2.89962
R28991 uo_out[5].n3 uo_out[5].t2 2.89962
R28992 uo_out[5].n3 uo_out[5].t8 2.89962
R28993 uo_out[5].n4 uo_out[5].t7 2.89962
R28994 uo_out[5].n4 uo_out[5].t1 2.89962
R28995 uo_out[5].n5 uo_out[5].t0 2.89962
R28996 uo_out[5].n5 uo_out[5].t6 2.89962
R28997 uo_out[5].n10 uo_out[5].n1 2.70811
R28998 uo_out[5].n0 uo_out[5].t4 2.06607
R28999 uo_out[5].n0 uo_out[5].t10 2.06607
R29000 uo_out[5].n1 uo_out[5].t5 2.06607
R29001 uo_out[5].n1 uo_out[5].t11 2.06607
R29002 uo_out[5].n7 uo_out[5].n6 0.877022
R29003 uo_out[5].n8 uo_out[5].n7 0.877022
R29004 uo_out[5].n10 uo_out[5].n9 0.803119
R29005 uo_out[5].n9 uo_out[5].n8 0.70537
R29006 uo_out[5] uo_out[5].n10 0.267929
R29007 clk.n0 clk.t11 31.7717
R29008 clk.n2 clk.t0 29.7439
R29009 clk.n2 clk.t12 18.7615
R29010 clk.n3 clk.t13 18.7615
R29011 clk.n4 clk.t7 18.7615
R29012 clk.n0 clk.t2 18.7615
R29013 clk.n1 clk.t5 18.7615
R29014 clk.n5 clk.t4 18.7615
R29015 clk.n2 clk.t1 11.133
R29016 clk.n3 clk.t3 11.133
R29017 clk.n4 clk.t6 11.133
R29018 clk.n0 clk.t8 11.133
R29019 clk.n1 clk.t10 11.133
R29020 clk.n5 clk.t9 11.133
R29021 clk.n3 clk.n2 10.5449
R29022 clk.n4 clk.n3 10.5449
R29023 clk.n1 clk.n0 10.5449
R29024 clk.n5 clk.n1 10.5449
R29025 clk.n5 clk.n4 10.5449
R29026 clk clk.n5 0.552085
R29027 _325_.A1.n21 _325_.A1.t16 19.7835
R29028 _325_.A1.n9 _325_.A1.t8 18.9805
R29029 _325_.A1.n18 _325_.A1.t12 17.5205
R29030 _325_.A1.n4 _325_.A1.t17 17.484
R29031 _325_.A1.n11 _325_.A1.t14 16.3768
R29032 _325_.A1.n2 _325_.A1.t10 16.3282
R29033 _325_.A1.n5 _325_.A1.t7 16.3282
R29034 _325_.A1.n13 _325_.A1.t4 16.2795
R29035 _325_.A1.n15 _325_.A1.t15 16.2795
R29036 _325_.A1.n13 _325_.A1.t5 15.2818
R29037 _325_.A1.n15 _325_.A1.t18 15.2818
R29038 _325_.A1.n5 _325_.A1.t19 14.7465
R29039 _325_.A1.n11 _325_.A1.t21 14.7222
R29040 _325_.A1.n2 _325_.A1.t20 14.6735
R29041 _325_.A1.n21 _325_.A1.t13 14.3085
R29042 _325_.A1.n4 _325_.A1.t9 11.863
R29043 _325_.A1.n18 _325_.A1.t11 11.5588
R29044 _325_.A1.n8 _325_.A1.n3 11.5205
R29045 _325_.A1.n9 _325_.A1.t6 11.4372
R29046 _325_.A1.n14 _325_.A1.n12 10.5446
R29047 _325_.A1.n14 _325_.A1 10.4087
R29048 _325_.A1.n10 _325_.A1 9.85858
R29049 _325_.A1.n17 _325_.A1.n16 9.3605
R29050 _325_.A1.n24 _325_.A1.n23 9.1805
R29051 _325_.A1.n20 _325_.A1.n17 8.5505
R29052 _325_.A1 _325_.A1.n13 8.17653
R29053 _325_.A1.n6 _325_.A1.n5 8.13432
R29054 _325_.A1 _325_.A1.n9 8.11457
R29055 _325_.A1 _325_.A1.n4 8.09965
R29056 _325_.A1.n16 _325_.A1.n15 8.02829
R29057 _325_.A1 _325_.A1.n21 8.00997
R29058 _325_.A1.n3 _325_.A1.n2 8.00405
R29059 _325_.A1.n19 _325_.A1.n18 8.0005
R29060 _325_.A1.n12 _325_.A1.n11 8.0005
R29061 _325_.A1.n7 _325_.A1.n6 7.11844
R29062 _325_.A1.n24 _325_.A1.n1 6.35795
R29063 _325_.A1.n23 _325_.A1.n22 5.5805
R29064 _325_.A1.n7 _325_.A1 5.48135
R29065 _325_.A1 _325_.A1.n0 5.26469
R29066 _325_.A1.n22 _325_.A1 4.73956
R29067 _325_.A1.n20 _325_.A1.n19 4.60296
R29068 _325_.A1.n8 _325_.A1.n7 4.5005
R29069 _325_.A1.n22 _325_.A1.n20 2.6105
R29070 _325_.A1.n1 _325_.A1.t3 1.99806
R29071 _325_.A1.n1 _325_.A1.t2 1.99806
R29072 _325_.A1.n0 _325_.A1.t0 1.4923
R29073 _325_.A1.n0 _325_.A1.t1 1.4923
R29074 _325_.A1.n10 _325_.A1.n8 1.4405
R29075 _325_.A1.n17 _325_.A1.n14 0.9005
R29076 _325_.A1.n23 _325_.A1.n10 0.5405
R29077 _325_.A1 _325_.A1.n24 0.396829
R29078 _325_.A1.n12 _325_.A1 0.211041
R29079 _325_.A1.n16 _325_.A1 0.148735
R29080 _325_.A1.n3 _325_.A1 0.133132
R29081 _325_.A1.n19 _325_.A1 0.0531154
R29082 _325_.A1.n6 _325_.A1 0.00286842
R29083 a_39124_27208.n3 a_39124_27208.t4 121.874
R29084 a_39124_27208.t4 a_39124_27208.t7 61.5152
R29085 a_39124_27208.n0 a_39124_27208.t5 52.378
R29086 a_39124_27208.n0 a_39124_27208.t6 17.7882
R29087 a_39124_27208.n2 a_39124_27208.t1 11.1158
R29088 a_39124_27208.n4 a_39124_27208.n3 9.95623
R29089 a_39124_27208.t0 a_39124_27208.n4 8.02846
R29090 a_39124_27208.n2 a_39124_27208.n1 8.0005
R29091 a_39124_27208.n3 a_39124_27208.t3 6.7165
R29092 a_39124_27208.n1 a_39124_27208.t2 5.96217
R29093 a_39124_27208.n1 a_39124_27208.n0 1.33883
R29094 a_39124_27208.n4 a_39124_27208.n2 0.376152
R29095 _330_.A1.n20 _330_.A1.n17 19.1705
R29096 _330_.A1.n18 _330_.A1.t7 18.6885
R29097 _330_.A1.n9 _330_.A1.t15 18.6885
R29098 _330_.A1.n21 _330_.A1.t6 16.4012
R29099 _330_.A1.n24 _330_.A1 16.3605
R29100 _330_.A1.n23 _330_.A1.t18 15.9023
R29101 _330_.A1.n16 _330_.A1.t5 15.3305
R29102 _330_.A1.n2 _330_.A1.t11 15.3305
R29103 _330_.A1.n12 _330_.A1.t22 15.3305
R29104 _330_.A1.n3 _330_.A1.t17 15.3305
R29105 _330_.A1.n5 _330_.A1.t12 15.3305
R29106 _330_.A1.n7 _330_.A1.t8 15.3305
R29107 _330_.A1.n16 _330_.A1.t20 15.148
R29108 _330_.A1.n2 _330_.A1.t4 15.148
R29109 _330_.A1.n12 _330_.A1.t21 15.148
R29110 _330_.A1.n3 _330_.A1.t9 15.148
R29111 _330_.A1.n5 _330_.A1.t23 15.148
R29112 _330_.A1.n7 _330_.A1.t16 15.148
R29113 _330_.A1.n22 _330_.A1.n20 14.9405
R29114 _330_.A1.n21 _330_.A1.t10 14.6735
R29115 _330_.A1.n23 _330_.A1.t19 13.4447
R29116 _330_.A1.n18 _330_.A1.t13 11.8873
R29117 _330_.A1.n9 _330_.A1.t14 11.8873
R29118 _330_.A1.n14 _330_.A1.n11 10.8005
R29119 _330_.A1.n10 _330_.A1 10.4257
R29120 _330_.A1.n11 _330_.A1.n10 10.2605
R29121 _330_.A1.n15 _330_.A1 9.86874
R29122 _330_.A1.n22 _330_.A1 9.7205
R29123 _330_.A1.n10 _330_.A1.n8 9.5405
R29124 _330_.A1.n25 _330_.A1.n24 9.0005
R29125 _330_.A1.n17 _330_.A1.n15 8.6405
R29126 _330_.A1 _330_.A1.n16 8.15932
R29127 _330_.A1 _330_.A1.n2 8.15932
R29128 _330_.A1 _330_.A1.n7 8.15932
R29129 _330_.A1 _330_.A1.n23 8.1305
R29130 _330_.A1 _330_.A1.n21 8.12809
R29131 _330_.A1.n13 _330_.A1.n12 8.01109
R29132 _330_.A1.n4 _330_.A1.n3 8.01109
R29133 _330_.A1.n6 _330_.A1.n5 8.01109
R29134 _330_.A1.n15 _330_.A1.n14 7.3805
R29135 _330_.A1.n25 _330_.A1.n1 6.69566
R29136 _330_.A1.n8 _330_.A1.n6 6.6605
R29137 _330_.A1.n17 _330_.A1 4.64874
R29138 _330_.A1.n8 _330_.A1 4.64874
R29139 _330_.A1.n20 _330_.A1.n19 4.58607
R29140 _330_.A1.n11 _330_.A1.n4 4.5005
R29141 _330_.A1.n14 _330_.A1.n13 4.5005
R29142 _330_.A1 _330_.A1.n9 4.08607
R29143 _330_.A1.n19 _330_.A1.n18 4.0005
R29144 _330_.A1 _330_.A1.n0 2.74964
R29145 _330_.A1.n0 _330_.A1.t0 2.06607
R29146 _330_.A1.n1 _330_.A1.t2 1.99806
R29147 _330_.A1.n1 _330_.A1.t3 1.99806
R29148 _330_.A1.n24 _330_.A1.n22 1.8905
R29149 _330_.A1.n0 _330_.A1.t1 1.4923
R29150 _330_.A1 _330_.A1.n25 0.33117
R29151 _330_.A1.n19 _330_.A1 0.245418
R29152 _330_.A1.n13 _330_.A1 0.148735
R29153 _330_.A1.n4 _330_.A1 0.148735
R29154 _330_.A1.n6 _330_.A1 0.148735
R29155 _416_.A1.n14 _416_.A1.n4 19.9355
R29156 _416_.A1.n1 _416_.A1.t10 19.4185
R29157 _416_.A1.n3 _416_.A1.t14 18.6885
R29158 _416_.A1.n9 _416_.A1.t11 17.703
R29159 _416_.A1.n4 _416_.A1.n2 16.6505
R29160 _416_.A1.n8 _416_.A1.n6 16.6505
R29161 _416_.A1.n7 _416_.A1.t5 15.3305
R29162 _416_.A1.n5 _416_.A1.t15 15.3305
R29163 _416_.A1.n10 _416_.A1.t12 15.3305
R29164 _416_.A1.n7 _416_.A1.t13 15.0872
R29165 _416_.A1.n5 _416_.A1.t9 15.0872
R29166 _416_.A1.n10 _416_.A1.t6 15.0872
R29167 _416_.A1.n9 _416_.A1.t8 14.8195
R29168 _416_.A1.n13 _416_.A1.n12 14.1755
R29169 _416_.A1.n13 _416_.A1.n8 12.5105
R29170 _416_.A1.n3 _416_.A1.t4 11.9603
R29171 _416_.A1.n1 _416_.A1.t7 11.6683
R29172 _416_.A1.n14 _416_.A1.n13 10.0805
R29173 _416_.A1 _416_.A1.n7 8.15932
R29174 _416_.A1.n6 _416_.A1.n5 8.01109
R29175 _416_.A1.n11 _416_.A1.n10 8.01109
R29176 _416_.A1 _416_.A1.n9 8.00997
R29177 _416_.A1.n2 _416_.A1.n1 8.0005
R29178 _416_.A1.n12 _416_.A1.n11 7.9655
R29179 _416_.A1.n15 _416_.A1.n0 6.78492
R29180 _416_.A1.n12 _416_.A1 5.26313
R29181 _416_.A1.n4 _416_.A1 4.5005
R29182 _416_.A1.n8 _416_.A1 4.5005
R29183 _416_.A1.n15 _416_.A1.n14 4.5005
R29184 _416_.A1 _416_.A1.n3 4.08607
R29185 _416_.A1.n0 _416_.A1.t2 3.413
R29186 _416_.A1.n0 _416_.A1.t3 3.413
R29187 _416_.A1 _416_.A1.n16 2.83361
R29188 _416_.A1.n16 _416_.A1.t0 2.06607
R29189 _416_.A1.n16 _416_.A1.t1 1.4923
R29190 _416_.A1 _416_.A1.n15 0.361668
R29191 _416_.A1.n6 _416_.A1 0.148735
R29192 _416_.A1.n11 _416_.A1 0.148735
R29193 _416_.A1.n2 _416_.A1 0.068
R29194 a_45508_20936.n3 a_45508_20936.t2 121.874
R29195 a_45508_20936.t2 a_45508_20936.t5 61.5152
R29196 a_45508_20936.n0 a_45508_20936.t7 52.378
R29197 a_45508_20936.n0 a_45508_20936.t4 17.7882
R29198 a_45508_20936.n2 a_45508_20936.t1 11.1158
R29199 a_45508_20936.n4 a_45508_20936.n3 9.95623
R29200 a_45508_20936.t0 a_45508_20936.n4 8.02846
R29201 a_45508_20936.n2 a_45508_20936.n1 8.0005
R29202 a_45508_20936.n3 a_45508_20936.t3 6.7165
R29203 a_45508_20936.n1 a_45508_20936.t6 5.96217
R29204 a_45508_20936.n1 a_45508_20936.n0 1.33883
R29205 a_45508_20936.n4 a_45508_20936.n2 0.376152
R29206 _424_.A2.n12 _424_.A2.n3 24.1362
R29207 _424_.A2.n7 _424_.A2.t9 19.1995
R29208 _424_.A2.n2 _424_.A2.t6 17.119
R29209 _424_.A2.n10 _424_.A2.t14 15.9023
R29210 _424_.A2.n6 _424_.A2.t11 15.9023
R29211 _424_.A2.n4 _424_.A2.t12 15.9023
R29212 _424_.A2.n9 _424_.A2.n5 13.6655
R29213 _424_.A2.n7 _424_.A2.t15 13.6028
R29214 _424_.A2.n10 _424_.A2.t8 13.4447
R29215 _424_.A2.n6 _424_.A2.t10 13.4447
R29216 _424_.A2.n4 _424_.A2.t7 13.4447
R29217 _424_.A2.n12 _424_.A2.n11 13.0505
R29218 _424_.A2.n2 _424_.A2.t13 12.7147
R29219 _424_.A2.n11 _424_.A2 9.1605
R29220 _424_.A2 _424_.A2.n10 8.1305
R29221 _424_.A2 _424_.A2.n6 8.1305
R29222 _424_.A2.n3 _424_.A2.n2 8.0005
R29223 _424_.A2 _424_.A2.n7 8.0005
R29224 _424_.A2.n5 _424_.A2.n4 8.0005
R29225 _424_.A2.n8 _424_.A2 7.7655
R29226 _424_.A2.n8 _424_.A2 7.1155
R29227 _424_.A2.n13 _424_.A2.n1 6.86529
R29228 _424_.A2.n9 _424_.A2.n8 6.4355
R29229 _424_.A2.n13 _424_.A2.n12 4.5005
R29230 _424_.A2 _424_.A2.n15 3.13612
R29231 _424_.A2.n14 _424_.A2.n0 2.71593
R29232 _424_.A2.n11 _424_.A2.n9 2.3405
R29233 _424_.A2.n1 _424_.A2.t4 1.99806
R29234 _424_.A2.n1 _424_.A2.t5 1.99806
R29235 _424_.A2.n0 _424_.A2.t0 1.61112
R29236 _424_.A2.n0 _424_.A2.t3 1.61112
R29237 _424_.A2.n15 _424_.A2.t2 1.61112
R29238 _424_.A2.n15 _424_.A2.t1 1.61112
R29239 _424_.A2.n14 _424_.A2.n13 0.650253
R29240 _424_.A2.n5 _424_.A2 0.1305
R29241 _424_.A2 _424_.A2.n14 0.096125
R29242 _424_.A2.n3 _424_.A2 0.0820131
R29243 _384_.A3.n11 _384_.A3.t11 19.4185
R29244 _384_.A3.n8 _384_.A3.t10 19.1995
R29245 _384_.A3.n9 _384_.A3.t17 17.484
R29246 _384_.A3.n11 _384_.A3.t13 16.535
R29247 _384_.A3.n15 _384_.A3.n14 16.2131
R29248 _384_.A3.n13 _384_.A3.t16 15.3305
R29249 _384_.A3.n13 _384_.A3.t14 15.0872
R29250 _384_.A3.n8 _384_.A3.t12 13.6028
R29251 _384_.A3.n9 _384_.A3.t15 11.863
R29252 _384_.A3.n12 _384_.A3.n10 10.5187
R29253 _384_.A3.n10 _384_.A3 9.5905
R29254 _384_.A3.n5 _384_.A3.n4 8.32963
R29255 _384_.A3 _384_.A3.n8 8.1405
R29256 _384_.A3 _384_.A3.n11 8.10362
R29257 _384_.A3 _384_.A3.n9 8.09965
R29258 _384_.A3.n14 _384_.A3.n13 8.0005
R29259 _384_.A3.n1 _384_.A3.t6 7.90366
R29260 _384_.A3.n5 _384_.A3.t7 7.44983
R29261 _384_.A3.n16 _384_.A3.n15 5.2205
R29262 _384_.A3.n7 _384_.A3.n6 5.2005
R29263 _384_.A3.n1 _384_.A3.n0 5.2005
R29264 _384_.A3.n3 _384_.A3.n2 5.2005
R29265 _384_.A3.n10 _384_.A3 4.85135
R29266 _384_.A3.n12 _384_.A3 4.6055
R29267 _384_.A3.n6 _384_.A3.t5 2.15435
R29268 _384_.A3.n6 _384_.A3.t8 2.15435
R29269 _384_.A3.n0 _384_.A3.t9 2.15435
R29270 _384_.A3.n0 _384_.A3.t4 2.15435
R29271 _384_.A3.n2 _384_.A3.t1 2.15435
R29272 _384_.A3.n2 _384_.A3.t0 2.15435
R29273 _384_.A3.n4 _384_.A3.t2 1.99806
R29274 _384_.A3.n4 _384_.A3.t3 1.99806
R29275 _384_.A3.n15 _384_.A3.n12 1.3955
R29276 _384_.A3.n7 _384_.A3.n5 0.655579
R29277 _384_.A3.n3 _384_.A3.n1 0.567306
R29278 _384_.A3 _384_.A3.n16 0.549879
R29279 _384_.A3.n14 _384_.A3 0.190411
R29280 _384_.A3 _384_.A3.n3 0.0598814
R29281 _384_.A3.n16 _384_.A3.n7 0.00792268
R29282 uo_out[7].n2 uo_out[7] 34.8896
R29283 uo_out[7].n2 uo_out[7].t4 8.29806
R29284 uo_out[7].n3 uo_out[7].n1 7.05647
R29285 uo_out[7].n4 uo_out[7].t2 4.17144
R29286 uo_out[7] uo_out[7].n0 2.88202
R29287 uo_out[7].n0 uo_out[7].t1 2.06607
R29288 uo_out[7].n1 uo_out[7].t3 1.99806
R29289 uo_out[7].n1 uo_out[7].t5 1.99806
R29290 uo_out[7].n0 uo_out[7].t0 1.4923
R29291 uo_out[7].n4 uo_out[7].n3 0.194466
R29292 uo_out[7] uo_out[7].n4 0.1885
R29293 uo_out[7].n3 uo_out[7].n2 0.0470517
R29294 uo_out[3].n6 uo_out[3] 26.6026
R29295 uo_out[3].n4 uo_out[3].n3 7.33746
R29296 uo_out[3].n4 uo_out[3].n2 6.46093
R29297 uo_out[3] uo_out[3].n0 5.81118
R29298 uo_out[3].n5 uo_out[3].n1 5.4118
R29299 uo_out[3].n2 uo_out[3].t6 3.6005
R29300 uo_out[3].n2 uo_out[3].t7 3.6005
R29301 uo_out[3].n3 uo_out[3].t5 3.6005
R29302 uo_out[3].n3 uo_out[3].t4 3.6005
R29303 uo_out[3].n0 uo_out[3].t2 2.06607
R29304 uo_out[3].n1 uo_out[3].t0 2.06607
R29305 uo_out[3].n0 uo_out[3].t1 1.4923
R29306 uo_out[3].n1 uo_out[3].t3 1.4923
R29307 uo_out[3].n5 uo_out[3].n4 0.439189
R29308 uo_out[3] uo_out[3].n6 0.158
R29309 uo_out[3].n6 uo_out[3].n5 0.0455
R29310 uio_in[0].n0 uio_in[0].t1 29.2005
R29311 uio_in[0].n0 uio_in[0].t0 12.1428
R29312 uio_in[0] uio_in[0].n0 8.19963
R29313 a_44784_25987.n0 a_44784_25987.t5 121.874
R29314 a_44784_25987.t5 a_44784_25987.t7 61.5152
R29315 a_44784_25987.n1 a_44784_25987.t3 52.378
R29316 a_44784_25987.n1 a_44784_25987.t2 17.7152
R29317 a_44784_25987.n3 a_44784_25987.t1 11.1158
R29318 a_44784_25987.n4 a_44784_25987.n0 9.95623
R29319 a_44784_25987.t0 a_44784_25987.n4 8.02846
R29320 a_44784_25987.n3 a_44784_25987.n2 8.0005
R29321 a_44784_25987.n0 a_44784_25987.t4 6.7165
R29322 a_44784_25987.n2 a_44784_25987.t6 6.023
R29323 a_44784_25987.n2 a_44784_25987.n1 1.33883
R29324 a_44784_25987.n4 a_44784_25987.n3 0.376152
R29325 _336_.A2.n5 _336_.A2.t10 22.2655
R29326 _336_.A2.n10 _336_.A2.t4 20.2945
R29327 _336_.A2.n0 _336_.A2.t2 19.1995
R29328 _336_.A2.n4 _336_.A2.t3 16.5715
R29329 _336_.A2.n9 _336_.A2.t6 16.3282
R29330 _336_.A2.n2 _336_.A2.t5 16.3282
R29331 _336_.A2.n9 _336_.A2.t7 15.6225
R29332 _336_.A2.n7 _336_.A2.n3 15.4805
R29333 _336_.A2.n4 _336_.A2.t11 15.4643
R29334 _336_.A2.n2 _336_.A2.t9 14.7465
R29335 _336_.A2.n0 _336_.A2.t8 13.6028
R29336 _336_.A2.n10 _336_.A2.t13 12.301
R29337 _336_.A2 _336_.A2.n12 11.3405
R29338 _336_.A2.n8 _336_.A2.n1 11.1605
R29339 _336_.A2.n5 _336_.A2.t12 9.77033
R29340 _336_.A2 _336_.A2.n4 9.01391
R29341 _336_.A2.n12 _336_.A2.n11 9.01236
R29342 _336_.A2 _336_.A2.t1 8.69622
R29343 _336_.A2 _336_.A2.n9 8.4405
R29344 _336_.A2.n3 _336_.A2.n2 8.00405
R29345 _336_.A2.n11 _336_.A2.n10 8.0005
R29346 _336_.A2.n6 _336_.A2.n5 8.0005
R29347 _336_.A2.n1 _336_.A2.n0 8.0005
R29348 _336_.A2.n8 _336_.A2.n7 6.8405
R29349 _336_.A2 _336_.A2.t0 6.72245
R29350 _336_.A2.n7 _336_.A2.n6 4.60663
R29351 _336_.A2.n12 _336_.A2.n8 1.8005
R29352 _336_.A2.n11 _336_.A2 0.311585
R29353 _336_.A2.n1 _336_.A2 0.1405
R29354 _336_.A2.n3 _336_.A2 0.133132
R29355 _336_.A2.n6 _336_.A2 0.0170789
R29356 a_41088_17757.n3 a_41088_17757.t2 121.874
R29357 a_41088_17757.t2 a_41088_17757.t7 61.5152
R29358 a_41088_17757.n0 a_41088_17757.t3 52.378
R29359 a_41088_17757.n0 a_41088_17757.t6 17.7882
R29360 a_41088_17757.n2 a_41088_17757.t1 11.1158
R29361 a_41088_17757.n4 a_41088_17757.n3 9.95623
R29362 a_41088_17757.t0 a_41088_17757.n4 8.02846
R29363 a_41088_17757.n2 a_41088_17757.n1 8.0005
R29364 a_41088_17757.n3 a_41088_17757.t4 6.7165
R29365 a_41088_17757.n1 a_41088_17757.t5 5.96217
R29366 a_41088_17757.n1 a_41088_17757.n0 1.33883
R29367 a_41088_17757.n4 a_41088_17757.n2 0.376152
R29368 a_24452_30344.n3 a_24452_30344.t5 121.874
R29369 a_24452_30344.t5 a_24452_30344.t7 61.5152
R29370 a_24452_30344.n0 a_24452_30344.t6 52.378
R29371 a_24452_30344.n0 a_24452_30344.t3 17.7882
R29372 a_24452_30344.n2 a_24452_30344.t1 11.1158
R29373 a_24452_30344.n4 a_24452_30344.n3 9.95623
R29374 a_24452_30344.t0 a_24452_30344.n4 8.02846
R29375 a_24452_30344.n2 a_24452_30344.n1 8.0005
R29376 a_24452_30344.n3 a_24452_30344.t2 6.7165
R29377 a_24452_30344.n1 a_24452_30344.t4 5.96217
R29378 a_24452_30344.n1 a_24452_30344.n0 1.33883
R29379 a_24452_30344.n4 a_24452_30344.n2 0.376152
R29380 a_32964_24072.n3 a_32964_24072.t7 121.874
R29381 a_32964_24072.t7 a_32964_24072.t6 61.5152
R29382 a_32964_24072.n0 a_32964_24072.t5 52.378
R29383 a_32964_24072.n0 a_32964_24072.t4 17.7882
R29384 a_32964_24072.n2 a_32964_24072.t1 11.1158
R29385 a_32964_24072.n4 a_32964_24072.n3 9.95623
R29386 a_32964_24072.t0 a_32964_24072.n4 8.02846
R29387 a_32964_24072.n2 a_32964_24072.n1 8.0005
R29388 a_32964_24072.n3 a_32964_24072.t3 6.7165
R29389 a_32964_24072.n1 a_32964_24072.t2 5.96217
R29390 a_32964_24072.n1 a_32964_24072.n0 1.33883
R29391 a_32964_24072.n4 a_32964_24072.n2 0.376152
R29392 _294_.ZN.n9 _294_.ZN.n8 25.4264
R29393 _294_.ZN.n7 _294_.ZN.t5 21.5355
R29394 _294_.ZN.n0 _294_.ZN.t3 21.5355
R29395 _294_.ZN.n4 _294_.ZN.n3 18.9805
R29396 _294_.ZN.n3 _294_.ZN.t8 15.8172
R29397 _294_.ZN.n4 _294_.ZN.t9 15.8172
R29398 _294_.ZN.n7 _294_.ZN.t4 9.91633
R29399 _294_.ZN.n2 _294_.ZN.t7 9.91633
R29400 _294_.ZN.n5 _294_.ZN.t6 9.91633
R29401 _294_.ZN.n0 _294_.ZN.t10 9.91633
R29402 _294_.ZN.n1 _294_.ZN.n0 9.26624
R29403 _294_.ZN.n6 _294_.ZN.n5 8.0005
R29404 _294_.ZN.n2 _294_.ZN.n1 8.0005
R29405 _294_.ZN.n8 _294_.ZN.n7 8.0005
R29406 _294_.ZN _294_.ZN.n10 6.8278
R29407 _294_.ZN.n3 _294_.ZN.n2 5.23217
R29408 _294_.ZN.n5 _294_.ZN.n4 5.23217
R29409 _294_.ZN.n9 _294_.ZN.t1 4.18853
R29410 _294_.ZN.n10 _294_.ZN.t2 2.89962
R29411 _294_.ZN.n10 _294_.ZN.t0 2.89962
R29412 _294_.ZN _294_.ZN.n6 1.17906
R29413 _294_.ZN.n6 _294_.ZN.n1 0.425606
R29414 _294_.ZN _294_.ZN.n9 0.158
R29415 _294_.ZN.n8 _294_.ZN 0.0177059
R29416 a_42596_27208.n3 a_42596_27208.t5 121.874
R29417 a_42596_27208.t5 a_42596_27208.t3 61.5152
R29418 a_42596_27208.n0 a_42596_27208.t2 52.378
R29419 a_42596_27208.n0 a_42596_27208.t7 17.7882
R29420 a_42596_27208.n2 a_42596_27208.t1 11.1158
R29421 a_42596_27208.n4 a_42596_27208.n3 9.95623
R29422 a_42596_27208.t0 a_42596_27208.n4 8.02846
R29423 a_42596_27208.n2 a_42596_27208.n1 8.0005
R29424 a_42596_27208.n3 a_42596_27208.t6 6.7165
R29425 a_42596_27208.n1 a_42596_27208.t4 5.96217
R29426 a_42596_27208.n1 a_42596_27208.n0 1.33883
R29427 a_42596_27208.n4 a_42596_27208.n2 0.376152
R29428 a_18404_30344.n3 a_18404_30344.t7 121.874
R29429 a_18404_30344.t7 a_18404_30344.t2 61.5152
R29430 a_18404_30344.n0 a_18404_30344.t4 52.378
R29431 a_18404_30344.n0 a_18404_30344.t5 17.7882
R29432 a_18404_30344.n2 a_18404_30344.t1 11.1158
R29433 a_18404_30344.n4 a_18404_30344.n3 9.99927
R29434 a_18404_30344.n2 a_18404_30344.n1 8.0005
R29435 a_18404_30344.n3 a_18404_30344.t3 6.7165
R29436 a_18404_30344.n1 a_18404_30344.t6 5.96217
R29437 a_18404_30344.t0 a_18404_30344.n4 5.40498
R29438 a_18404_30344.n1 a_18404_30344.n0 1.33883
R29439 a_18404_30344.n4 a_18404_30344.n2 0.333109
R29440 _417_.A2.n9 _417_.A2.n5 19.7318
R29441 _417_.A2.n7 _417_.A2.t12 19.5645
R29442 _417_.A2.n3 _417_.A2.t9 19.4185
R29443 _417_.A2.n10 _417_.A2.t7 18.6885
R29444 _417_.A2.n7 _417_.A2.t8 18.4938
R29445 _417_.A2.n1 _417_.A2.t3 17.484
R29446 _417_.A2.n6 _417_.A2.t11 16.7662
R29447 _417_.A2.n3 _417_.A2.t10 16.535
R29448 _417_.A2.n5 _417_.A2.n2 15.5072
R29449 _417_.A2.n6 _417_.A2.t5 14.3815
R29450 _417_.A2 _417_.A2.n12 13.1405
R29451 _417_.A2.n10 _417_.A2.t4 11.9603
R29452 _417_.A2.n1 _417_.A2.t6 11.863
R29453 _417_.A2.n9 _417_.A2.n8 11.5205
R29454 _417_.A2.n12 _417_.A2.n11 9.0005
R29455 _417_.A2.n8 _417_.A2.n6 8.57871
R29456 _417_.A2 _417_.A2.t2 8.56922
R29457 _417_.A2 _417_.A2.n7 8.16594
R29458 _417_.A2.n2 _417_.A2.n1 8.0005
R29459 _417_.A2.n4 _417_.A2.n3 8.0005
R29460 _417_.A2.n5 _417_.A2.n4 4.68238
R29461 _417_.A2.n11 _417_.A2.n10 4.08017
R29462 _417_.A2 _417_.A2.n0 3.27068
R29463 _417_.A2.n0 _417_.A2.t1 1.61112
R29464 _417_.A2.n0 _417_.A2.t0 1.61112
R29465 _417_.A2.n8 _417_.A2 0.57628
R29466 _417_.A2.n12 _417_.A2.n9 0.4505
R29467 _417_.A2.n11 _417_.A2 0.165746
R29468 _417_.A2.n4 _417_.A2 0.103625
R29469 _417_.A2.n2 _417_.A2 0.0996525
R29470 a_49936_19325.n3 a_49936_19325.t3 121.874
R29471 a_49936_19325.t3 a_49936_19325.t5 61.5152
R29472 a_49936_19325.n0 a_49936_19325.t2 52.378
R29473 a_49936_19325.n0 a_49936_19325.t7 17.7882
R29474 a_49936_19325.n2 a_49936_19325.t1 11.1158
R29475 a_49936_19325.n4 a_49936_19325.n3 9.95623
R29476 a_49936_19325.t0 a_49936_19325.n4 8.02846
R29477 a_49936_19325.n2 a_49936_19325.n1 8.0005
R29478 a_49936_19325.n3 a_49936_19325.t4 6.7165
R29479 a_49936_19325.n1 a_49936_19325.t6 5.96217
R29480 a_49936_19325.n1 a_49936_19325.n0 1.33883
R29481 a_49936_19325.n4 a_49936_19325.n2 0.376152
R29482 _281_.ZN.n7 _281_.ZN.n6 20.9505
R29483 _281_.ZN.n4 _281_.ZN.t8 19.5645
R29484 _281_.ZN.n2 _281_.ZN.t5 19.4185
R29485 _281_.ZN.n1 _281_.ZN.t9 18.6885
R29486 _281_.ZN.n4 _281_.ZN.t7 17.1312
R29487 _281_.ZN.n2 _281_.ZN.t6 16.535
R29488 _281_.ZN.n1 _281_.ZN.t4 11.8873
R29489 _281_.ZN.n3 _281_.ZN 11.2205
R29490 _281_.ZN.n3 _281_.ZN 10.3689
R29491 _281_.ZN.n6 _281_.ZN.n3 9.6755
R29492 _281_.ZN.n7 _281_.ZN.t1 8.29806
R29493 _281_.ZN _281_.ZN.n2 8.10362
R29494 _281_.ZN.n5 _281_.ZN.n4 8.0005
R29495 _281_.ZN.n8 _281_.ZN.t0 4.50873
R29496 _281_.ZN.n6 _281_.ZN.n5 4.5005
R29497 _281_.ZN _281_.ZN.n1 4.24542
R29498 _281_.ZN _281_.ZN.n0 2.89216
R29499 _281_.ZN.n0 _281_.ZN.t3 1.84822
R29500 _281_.ZN.n0 _281_.ZN.t2 1.84822
R29501 _281_.ZN.n8 _281_.ZN.n7 0.542363
R29502 _281_.ZN _281_.ZN.n8 0.215857
R29503 _281_.ZN.n5 _281_.ZN 0.1125
R29504 _411_.A2.n9 _411_.A2 20.7036
R29505 _411_.A2.n6 _411_.A2.t12 19.5645
R29506 _411_.A2.n8 _411_.A2.t8 18.9805
R29507 _411_.A2.n10 _411_.A2.t10 18.6885
R29508 _411_.A2.n6 _411_.A2.t9 18.4938
R29509 _411_.A2.n5 _411_.A2.t11 16.7662
R29510 _411_.A2.n5 _411_.A2.t13 14.3815
R29511 _411_.A2.n10 _411_.A2.t15 11.8873
R29512 _411_.A2.n8 _411_.A2.t14 11.4372
R29513 _411_.A2.n11 _411_.A2 11.3405
R29514 _411_.A2.n12 _411_.A2.n11 10.2605
R29515 _411_.A2.n9 _411_.A2.n7 10.1705
R29516 _411_.A2.n7 _411_.A2.n5 8.38432
R29517 _411_.A2 _411_.A2.n6 8.16594
R29518 _411_.A2 _411_.A2.n8 8.11457
R29519 _411_.A2 _411_.A2.n13 6.79383
R29520 _411_.A2.n2 _411_.A2.n0 5.98178
R29521 _411_.A2.n4 _411_.A2.n3 5.2005
R29522 _411_.A2.n2 _411_.A2.n1 5.2005
R29523 _411_.A2 _411_.A2.n10 4.24542
R29524 _411_.A2.n11 _411_.A2.n9 2.3405
R29525 _411_.A2.n13 _411_.A2.t2 1.99806
R29526 _411_.A2.n13 _411_.A2.t3 1.99806
R29527 _411_.A2.n0 _411_.A2.t5 1.84822
R29528 _411_.A2.n0 _411_.A2.t7 1.84822
R29529 _411_.A2.n3 _411_.A2.t6 1.84822
R29530 _411_.A2.n3 _411_.A2.t4 1.84822
R29531 _411_.A2.n1 _411_.A2.t0 1.84822
R29532 _411_.A2.n1 _411_.A2.t1 1.84822
R29533 _411_.A2.n7 _411_.A2 0.816321
R29534 _411_.A2.n12 _411_.A2.n4 0.800989
R29535 _411_.A2.n4 _411_.A2.n2 0.781777
R29536 _411_.A2 _411_.A2.n12 0.631974
R29537 _294_.A2 _294_.A2.n9 20.8805
R29538 _294_.A2.n5 _294_.A2.n4 20.6511
R29539 _294_.A2.n0 _294_.A2.t2 18.6885
R29540 _294_.A2.n6 _294_.A2.t7 18.6885
R29541 _294_.A2.n1 _294_.A2.t9 18.6885
R29542 _294_.A2.n3 _294_.A2.t6 18.6885
R29543 _294_.A2.n6 _294_.A2.t4 11.9603
R29544 _294_.A2.n3 _294_.A2.t3 11.9603
R29545 _294_.A2.n0 _294_.A2.t8 11.8873
R29546 _294_.A2.n1 _294_.A2.t5 11.8873
R29547 _294_.A2.n9 _294_.A2.n8 10.0237
R29548 _294_.A2 _294_.A2.t1 9.70112
R29549 _294_.A2.n8 _294_.A2.n5 9.12366
R29550 _294_.A2.n8 _294_.A2.n7 9.08607
R29551 _294_.A2.n5 _294_.A2.n2 5.39607
R29552 _294_.A2.n9 _294_.A2 4.66575
R29553 _294_.A2 _294_.A2.t0 4.43672
R29554 _294_.A2 _294_.A2.n0 4.24542
R29555 _294_.A2.n7 _294_.A2.n6 4.0005
R29556 _294_.A2.n2 _294_.A2.n1 4.0005
R29557 _294_.A2.n4 _294_.A2.n3 4.0005
R29558 _294_.A2.n7 _294_.A2 0.245418
R29559 _294_.A2.n2 _294_.A2 0.245418
R29560 _294_.A2.n4 _294_.A2 0.245418
R29561 a_21652_27591.n0 a_21652_27591.t7 121.874
R29562 a_21652_27591.t7 a_21652_27591.t4 61.5152
R29563 a_21652_27591.n1 a_21652_27591.t2 52.378
R29564 a_21652_27591.n1 a_21652_27591.t3 17.7152
R29565 a_21652_27591.n3 a_21652_27591.t1 11.1158
R29566 a_21652_27591.n4 a_21652_27591.n0 9.95623
R29567 a_21652_27591.t0 a_21652_27591.n4 8.02846
R29568 a_21652_27591.n3 a_21652_27591.n2 8.0005
R29569 a_21652_27591.n0 a_21652_27591.t5 6.7165
R29570 a_21652_27591.n2 a_21652_27591.t6 6.023
R29571 a_21652_27591.n2 a_21652_27591.n1 1.33883
R29572 a_21652_27591.n4 a_21652_27591.n3 0.376152
R29573 a_32740_22504.n3 a_32740_22504.t3 121.874
R29574 a_32740_22504.t3 a_32740_22504.t6 61.5152
R29575 a_32740_22504.n0 a_32740_22504.t5 52.378
R29576 a_32740_22504.n0 a_32740_22504.t2 17.7882
R29577 a_32740_22504.n2 a_32740_22504.t1 11.1158
R29578 a_32740_22504.n4 a_32740_22504.n3 9.95623
R29579 a_32740_22504.t0 a_32740_22504.n4 8.02846
R29580 a_32740_22504.n2 a_32740_22504.n1 8.0005
R29581 a_32740_22504.n3 a_32740_22504.t7 6.7165
R29582 a_32740_22504.n1 a_32740_22504.t4 5.96217
R29583 a_32740_22504.n1 a_32740_22504.n0 1.33883
R29584 a_32740_22504.n4 a_32740_22504.n2 0.376152
R29585 a_31508_29159.n0 a_31508_29159.t3 121.874
R29586 a_31508_29159.t3 a_31508_29159.t6 61.5152
R29587 a_31508_29159.n1 a_31508_29159.t7 52.378
R29588 a_31508_29159.n1 a_31508_29159.t5 17.7152
R29589 a_31508_29159.n3 a_31508_29159.t1 11.1158
R29590 a_31508_29159.n4 a_31508_29159.n0 9.95623
R29591 a_31508_29159.t0 a_31508_29159.n4 8.02846
R29592 a_31508_29159.n3 a_31508_29159.n2 8.0005
R29593 a_31508_29159.n0 a_31508_29159.t4 6.7165
R29594 a_31508_29159.n2 a_31508_29159.t2 6.023
R29595 a_31508_29159.n2 a_31508_29159.n1 1.33883
R29596 a_31508_29159.n4 a_31508_29159.n3 0.376152
R29597 a_35092_19368.n3 a_35092_19368.t7 121.874
R29598 a_35092_19368.t7 a_35092_19368.t3 61.5152
R29599 a_35092_19368.n0 a_35092_19368.t2 52.378
R29600 a_35092_19368.n0 a_35092_19368.t6 17.7882
R29601 a_35092_19368.n2 a_35092_19368.t1 11.1158
R29602 a_35092_19368.n4 a_35092_19368.n3 9.95623
R29603 a_35092_19368.t0 a_35092_19368.n4 8.02846
R29604 a_35092_19368.n2 a_35092_19368.n1 8.0005
R29605 a_35092_19368.n3 a_35092_19368.t5 6.7165
R29606 a_35092_19368.n1 a_35092_19368.t4 5.96217
R29607 a_35092_19368.n1 a_35092_19368.n0 1.33883
R29608 a_35092_19368.n4 a_35092_19368.n2 0.376152
R29609 a_33748_20936.n3 a_33748_20936.t2 121.874
R29610 a_33748_20936.t2 a_33748_20936.t7 61.5152
R29611 a_33748_20936.n0 a_33748_20936.t6 52.378
R29612 a_33748_20936.n0 a_33748_20936.t5 17.7882
R29613 a_33748_20936.n2 a_33748_20936.t1 11.1158
R29614 a_33748_20936.n4 a_33748_20936.n3 9.95623
R29615 a_33748_20936.t0 a_33748_20936.n4 8.02846
R29616 a_33748_20936.n2 a_33748_20936.n1 8.0005
R29617 a_33748_20936.n3 a_33748_20936.t4 6.7165
R29618 a_33748_20936.n1 a_33748_20936.t3 5.96217
R29619 a_33748_20936.n1 a_33748_20936.n0 1.33883
R29620 a_33748_20936.n4 a_33748_20936.n2 0.376152
R29621 _363_.Z.n0 _363_.Z.t3 20.5135
R29622 _363_.Z.n1 _363_.Z.t9 18.5425
R29623 _363_.Z.n3 _363_.Z.t2 16.3282
R29624 _363_.Z.n5 _363_.Z.t4 15.3305
R29625 _363_.Z.n5 _363_.Z.t8 15.0872
R29626 _363_.Z.n3 _363_.Z.t7 14.6735
R29627 _363_.Z.n1 _363_.Z.t5 14.053
R29628 _363_.Z _363_.Z.n8 11.7455
R29629 _363_.Z.n0 _363_.Z.t6 11.4372
R29630 _363_.Z.n8 _363_.Z.n7 10.4405
R29631 _363_.Z.n8 _363_.Z.n2 10.4405
R29632 _363_.Z _363_.Z.n0 8.96449
R29633 _363_.Z.n2 _363_.Z.n1 8.89427
R29634 _363_.Z _363_.Z.t1 8.62678
R29635 _363_.Z.n6 _363_.Z.n5 8.10306
R29636 _363_.Z.n4 _363_.Z.n3 8.0005
R29637 _363_.Z.n7 _363_.Z.n4 6.51366
R29638 _363_.Z.n7 _363_.Z.n6 4.50259
R29639 _363_.Z _363_.Z.t0 4.30606
R29640 _363_.Z.n2 _363_.Z 0.187167
R29641 _363_.Z.n6 _363_.Z 0.0878529
R29642 _363_.Z.n4 _363_.Z 0.00997368
R29643 a_28596_27916.n9 a_28596_27916.n8 5.2005
R29644 a_28596_27916.n7 a_28596_27916.n6 5.2005
R29645 a_28596_27916.n5 a_28596_27916.n4 5.2005
R29646 a_28596_27916.n3 a_28596_27916.n2 5.2005
R29647 a_28596_27916.t3 a_28596_27916.n9 4.99956
R29648 a_28596_27916.n1 a_28596_27916.t7 4.88774
R29649 a_28596_27916.n2 a_28596_27916.t6 3.1505
R29650 a_28596_27916.n1 a_28596_27916.n0 2.6005
R29651 a_28596_27916.n2 a_28596_27916.t1 1.51717
R29652 a_28596_27916.n4 a_28596_27916.t10 1.51717
R29653 a_28596_27916.n4 a_28596_27916.t8 1.51717
R29654 a_28596_27916.n6 a_28596_27916.t0 1.51717
R29655 a_28596_27916.n6 a_28596_27916.t2 1.51717
R29656 a_28596_27916.n8 a_28596_27916.t9 1.51717
R29657 a_28596_27916.n8 a_28596_27916.t11 1.51717
R29658 a_28596_27916.n0 a_28596_27916.t4 1.51717
R29659 a_28596_27916.n0 a_28596_27916.t5 1.51717
R29660 a_28596_27916.n3 a_28596_27916.n1 0.902492
R29661 a_28596_27916.n9 a_28596_27916.n7 0.798761
R29662 a_28596_27916.n7 a_28596_27916.n5 0.798761
R29663 a_28596_27916.n5 a_28596_27916.n3 0.798761
R29664 a_32180_25640.n3 a_32180_25640.t6 121.874
R29665 a_32180_25640.t6 a_32180_25640.t4 61.5152
R29666 a_32180_25640.n0 a_32180_25640.t3 52.378
R29667 a_32180_25640.n0 a_32180_25640.t2 17.7882
R29668 a_32180_25640.n2 a_32180_25640.t1 11.1158
R29669 a_32180_25640.n4 a_32180_25640.n3 9.95623
R29670 a_32180_25640.t0 a_32180_25640.n4 8.02846
R29671 a_32180_25640.n2 a_32180_25640.n1 8.0005
R29672 a_32180_25640.n3 a_32180_25640.t5 6.7165
R29673 a_32180_25640.n1 a_32180_25640.t7 5.96217
R29674 a_32180_25640.n1 a_32180_25640.n0 1.33883
R29675 a_32180_25640.n4 a_32180_25640.n2 0.376152
R29676 _284_.A2.n8 _284_.A2 30.713
R29677 _284_.A2.n7 _284_.A2.t9 15.7077
R29678 _284_.A2.n0 _284_.A2.t3 15.5617
R29679 _284_.A2.n2 _284_.A2.t5 14.7465
R29680 _284_.A2.n5 _284_.A2.t8 14.7465
R29681 _284_.A2.n0 _284_.A2.t4 14.7465
R29682 _284_.A2.n7 _284_.A2.t2 14.6005
R29683 _284_.A2.n4 _284_.A2.n3 13.3198
R29684 _284_.A2.n3 _284_.A2.t7 12.0455
R29685 _284_.A2.n4 _284_.A2.t6 12.0455
R29686 _284_.A2.n1 _284_.A2.n0 9.40137
R29687 _284_.A2 _284_.A2.n7 8.81272
R29688 _284_.A2 _284_.A2.t1 8.52139
R29689 _284_.A2.n6 _284_.A2.n5 8.0005
R29690 _284_.A2.n2 _284_.A2.n1 8.0005
R29691 _284_.A2.n8 _284_.A2.t0 4.09844
R29692 _284_.A2.n3 _284_.A2.n2 1.99583
R29693 _284_.A2.n5 _284_.A2.n4 1.99583
R29694 _284_.A2.n6 _284_.A2.n1 0.39963
R29695 _284_.A2 _284_.A2.n6 0.373002
R29696 _284_.A2 _284_.A2.n8 0.218
R29697 a_53744_22851.n0 a_53744_22851.t6 121.874
R29698 a_53744_22851.t6 a_53744_22851.t3 61.5152
R29699 a_53744_22851.n1 a_53744_22851.t4 52.378
R29700 a_53744_22851.n1 a_53744_22851.t5 17.7152
R29701 a_53744_22851.n3 a_53744_22851.t1 11.1158
R29702 a_53744_22851.n4 a_53744_22851.n0 9.95623
R29703 a_53744_22851.t0 a_53744_22851.n4 8.02846
R29704 a_53744_22851.n3 a_53744_22851.n2 8.0005
R29705 a_53744_22851.n0 a_53744_22851.t7 6.7165
R29706 a_53744_22851.n2 a_53744_22851.t2 6.023
R29707 a_53744_22851.n2 a_53744_22851.n1 1.33883
R29708 a_53744_22851.n4 a_53744_22851.n3 0.376152
R29709 ui_in[1].n0 ui_in[1].t1 20.1607
R29710 ui_in[1].n1 ui_in[1] 16.3517
R29711 ui_in[1].n0 ui_in[1].t0 10.8288
R29712 ui_in[1].n1 ui_in[1].n0 8.0005
R29713 ui_in[1] ui_in[1].n1 0.065101
R29714 _397_.A1.n1 _397_.A1.t13 25.4288
R29715 _397_.A1.n13 _397_.A1.t3 22.1195
R29716 _397_.A1.n14 _397_.A1.t2 19.5645
R29717 _397_.A1.n3 _397_.A1.t15 18.9805
R29718 _397_.A1.n14 _397_.A1.t9 18.4938
R29719 _397_.A1.n5 _397_.A1 17.5536
R29720 _397_.A1.n0 _397_.A1.t12 17.5205
R29721 _397_.A1.n6 _397_.A1.n5 17.2805
R29722 _397_.A1.n9 _397_.A1.t8 16.7783
R29723 _397_.A1.n8 _397_.A1.t14 16.7783
R29724 _397_.A1.n9 _397_.A1.n8 16.5048
R29725 _397_.A1.n4 _397_.A1.t4 16.2795
R29726 _397_.A1.n4 _397_.A1.t11 15.2818
R29727 _397_.A1.n6 _397_.A1.n2 14.608
R29728 _397_.A1.n17 _397_.A1 11.8556
R29729 _397_.A1.n0 _397_.A1.t10 11.5588
R29730 _397_.A1.n10 _397_.A1.t6 11.5588
R29731 _397_.A1.n7 _397_.A1.t5 11.5588
R29732 _397_.A1.n3 _397_.A1.t17 11.4372
R29733 _397_.A1.n1 _397_.A1.t7 10.5247
R29734 _397_.A1.n12 _397_.A1 9.1805
R29735 _397_.A1.n13 _397_.A1.t16 9.02817
R29736 _397_.A1 _397_.A1.n17 9.0005
R29737 _397_.A1 _397_.A1.t1 8.69622
R29738 _397_.A1 _397_.A1.n13 8.35407
R29739 _397_.A1.n15 _397_.A1.n14 8.33318
R29740 _397_.A1.n11 _397_.A1.n7 8.28737
R29741 _397_.A1 _397_.A1.n4 8.17653
R29742 _397_.A1 _397_.A1.n3 8.11576
R29743 _397_.A1 _397_.A1.n0 8.05312
R29744 _397_.A1.n11 _397_.A1.n10 8.0005
R29745 _397_.A1.n2 _397_.A1.n1 8.0005
R29746 _397_.A1.n16 _397_.A1.n12 6.8405
R29747 _397_.A1 _397_.A1.t0 6.72245
R29748 _397_.A1.n17 _397_.A1.n16 6.1205
R29749 _397_.A1.n5 _397_.A1 4.64874
R29750 _397_.A1.n16 _397_.A1.n15 4.5005
R29751 _397_.A1.n12 _397_.A1.n6 1.4405
R29752 _397_.A1 _397_.A1.n11 0.950062
R29753 _397_.A1.n10 _397_.A1.n9 0.3655
R29754 _397_.A1.n8 _397_.A1.n7 0.3655
R29755 _397_.A1.n15 _397_.A1 0.1805
R29756 _397_.A1.n2 _397_.A1 0.113
R29757 ui_in[7].n1 ui_in[7].t1 28.5995
R29758 ui_in[7].n0 ui_in[7].t0 18.7493
R29759 ui_in[7].n2 ui_in[7] 17.157
R29760 ui_in[7].n0 ui_in[7].t2 12.1672
R29761 ui_in[7].n2 ui_in[7].n1 2.66717
R29762 ui_in[7].n1 ui_in[7].n0 1.0005
R29763 ui_in[7] ui_in[7].n2 0.0290366
R29764 ui_in[2].n0 ui_in[2].t0 20.1607
R29765 ui_in[2].n1 ui_in[2] 17.6117
R29766 ui_in[2].n0 ui_in[2].t1 10.8288
R29767 ui_in[2].n1 ui_in[2].n0 8.0005
R29768 ui_in[2] ui_in[2].n1 0.065101
R29769 uio_oe[0] uio_oe[0].t0 8.31126
R29770 _451_.Q.n14 _451_.Q.t3 20.2945
R29771 _451_.Q.n11 _451_.Q.t13 19.7105
R29772 _451_.Q.n4 _451_.Q.t4 19.1995
R29773 _451_.Q.n1 _451_.Q.t6 18.6885
R29774 _451_.Q.n7 _451_.Q.n3 17.8205
R29775 _451_.Q.n0 _451_.Q.t15 17.7395
R29776 _451_.Q.n5 _451_.Q.t9 17.5692
R29777 _451_.Q.n13 _451_.Q.t5 16.3282
R29778 _451_.Q.n8 _451_.Q.t17 16.3282
R29779 _451_.Q.n5 _451_.Q.t2 16.1335
R29780 _451_.Q.n13 _451_.Q.t12 15.6955
R29781 _451_.Q.n8 _451_.Q.t14 14.7465
R29782 _451_.Q.n11 _451_.Q.t11 14.3085
R29783 _451_.Q.n4 _451_.Q.t7 13.6637
R29784 _451_.Q.n0 _451_.Q.t8 12.6782
R29785 _451_.Q.n14 _451_.Q.t16 12.301
R29786 _451_.Q.n1 _451_.Q.t10 11.8873
R29787 _451_.Q.n3 _451_.Q 11.7005
R29788 _451_.Q.n6 _451_.Q 10.0805
R29789 _451_.Q _451_.Q.n16 10.0805
R29790 _451_.Q.n16 _451_.Q.n15 9.73236
R29791 _451_.Q.n3 _451_.Q.n2 9.44607
R29792 _451_.Q.n6 _451_.Q 9.1805
R29793 _451_.Q _451_.Q.t1 8.69622
R29794 _451_.Q _451_.Q.n13 8.4405
R29795 _451_.Q.n10 _451_.Q.n7 8.2805
R29796 _451_.Q _451_.Q.n4 8.1405
R29797 _451_.Q.n9 _451_.Q.n8 8.13432
R29798 _451_.Q _451_.Q.n5 8.02303
R29799 _451_.Q _451_.Q.n11 8.00997
R29800 _451_.Q.n15 _451_.Q.n14 8.0005
R29801 _451_.Q _451_.Q.t0 6.72245
R29802 _451_.Q.n12 _451_.Q 5.89313
R29803 _451_.Q.n16 _451_.Q.n12 5.2205
R29804 _451_.Q.n10 _451_.Q.n9 4.59844
R29805 _451_.Q _451_.Q.n0 4.07694
R29806 _451_.Q.n2 _451_.Q.n1 4.0005
R29807 _451_.Q.n7 _451_.Q.n6 1.8005
R29808 _451_.Q.n15 _451_.Q 0.311585
R29809 _451_.Q.n2 _451_.Q 0.245418
R29810 _451_.Q.n12 _451_.Q.n10 0.1805
R29811 _451_.Q.n9 _451_.Q 0.00286842
R29812 a_52064_19715.n0 a_52064_19715.t5 121.874
R29813 a_52064_19715.t5 a_52064_19715.t7 61.5152
R29814 a_52064_19715.n1 a_52064_19715.t2 52.378
R29815 a_52064_19715.n1 a_52064_19715.t4 17.7152
R29816 a_52064_19715.n3 a_52064_19715.t1 11.1158
R29817 a_52064_19715.n4 a_52064_19715.n0 9.95623
R29818 a_52064_19715.t0 a_52064_19715.n4 8.02846
R29819 a_52064_19715.n3 a_52064_19715.n2 8.0005
R29820 a_52064_19715.n0 a_52064_19715.t3 6.7165
R29821 a_52064_19715.n2 a_52064_19715.t6 6.023
R29822 a_52064_19715.n2 a_52064_19715.n1 1.33883
R29823 a_52064_19715.n4 a_52064_19715.n3 0.376152
R29824 _337_.A3.n8 _337_.A3.n7 30.4701
R29825 _337_.A3.n2 _337_.A3.n1 30.4701
R29826 _337_.A3.n13 _337_.A3.t7 20.1161
R29827 _337_.A3.n8 _337_.A3.t14 19.0535
R29828 _337_.A3.n7 _337_.A3.t15 19.0535
R29829 _337_.A3.n1 _337_.A3.t13 19.0535
R29830 _337_.A3.n2 _337_.A3.t9 19.0535
R29831 _337_.A3.n13 _337_.A3.t10 18.2505
R29832 _337_.A3.n11 _337_.A3.t12 17.8003
R29833 _337_.A3.n14 _337_.A3.t5 17.3623
R29834 _337_.A3.n16 _337_.A3.n15 17.0026
R29835 _337_.A3.n12 _337_.A3 15.7596
R29836 _337_.A3.n11 _337_.A3.t4 14.7465
R29837 _337_.A3.n14 _337_.A3.t2 14.6735
R29838 _337_.A3.n9 _337_.A3.t11 10.5612
R29839 _337_.A3.n6 _337_.A3.t6 10.5612
R29840 _337_.A3.n0 _337_.A3.t3 10.5612
R29841 _337_.A3.n3 _337_.A3.t8 10.5612
R29842 _337_.A3 _337_.A3.n13 9.79005
R29843 _337_.A3 _337_.A3.t1 8.69622
R29844 _337_.A3.n4 _337_.A3.n0 8.54637
R29845 _337_.A3 _337_.A3.n11 8.11418
R29846 _337_.A3.n15 _337_.A3.n14 8.0005
R29847 _337_.A3.n4 _337_.A3.n3 8.0005
R29848 _337_.A3.n6 _337_.A3.n5 8.0005
R29849 _337_.A3.n10 _337_.A3.n9 8.0005
R29850 _337_.A3 _337_.A3.t0 6.72245
R29851 _337_.A3.n12 _337_.A3 6.2105
R29852 _337_.A3 _337_.A3.n16 4.5005
R29853 _337_.A3.n9 _337_.A3.n8 4.2345
R29854 _337_.A3.n7 _337_.A3.n6 4.2345
R29855 _337_.A3.n1 _337_.A3.n0 4.2345
R29856 _337_.A3.n3 _337_.A3.n2 4.2345
R29857 _337_.A3.n16 _337_.A3.n12 1.2605
R29858 _337_.A3.n5 _337_.A3.n4 1.19007
R29859 _337_.A3.n10 _337_.A3.n5 0.518884
R29860 _337_.A3 _337_.A3.n10 0.0873675
R29861 _337_.A3.n15 _337_.A3 0.0217143
R29862 a_35204_24455.n0 a_35204_24455.t6 121.874
R29863 a_35204_24455.t6 a_35204_24455.t4 61.5152
R29864 a_35204_24455.n1 a_35204_24455.t2 52.378
R29865 a_35204_24455.n1 a_35204_24455.t3 17.7152
R29866 a_35204_24455.n3 a_35204_24455.t1 11.1158
R29867 a_35204_24455.n4 a_35204_24455.n0 9.95623
R29868 a_35204_24455.t0 a_35204_24455.n4 8.02846
R29869 a_35204_24455.n3 a_35204_24455.n2 8.0005
R29870 a_35204_24455.n0 a_35204_24455.t7 6.7165
R29871 a_35204_24455.n2 a_35204_24455.t5 6.023
R29872 a_35204_24455.n2 a_35204_24455.n1 1.33883
R29873 a_35204_24455.n4 a_35204_24455.n3 0.376152
R29874 _325_.A2.n6 _325_.A2.t6 27.9595
R29875 _325_.A2.n2 _325_.A2.t7 17.484
R29876 _325_.A2.n0 _325_.A2.t2 16.3282
R29877 _325_.A2.n4 _325_.A2.t11 16.3282
R29878 _325_.A2.n9 _325_.A2.t9 15.3305
R29879 _325_.A2.n9 _325_.A2.t8 15.148
R29880 _325_.A2.n4 _325_.A2.t4 14.7465
R29881 _325_.A2.n0 _325_.A2.t3 14.6735
R29882 _325_.A2.n5 _325_.A2 12.1955
R29883 _325_.A2.n2 _325_.A2.t5 11.863
R29884 _325_.A2.n11 _325_.A2.n10 10.8005
R29885 _325_.A2.n12 _325_.A2.n11 9.56943
R29886 _325_.A2.n8 _325_.A2.n7 9.1805
R29887 _325_.A2.n12 _325_.A2.t1 8.31032
R29888 _325_.A2 _325_.A2.n2 8.09965
R29889 _325_.A2.n10 _325_.A2.n9 8.01109
R29890 _325_.A2.n1 _325_.A2.n0 8.0005
R29891 _325_.A2.n7 _325_.A2.n6 8.0005
R29892 _325_.A2 _325_.A2.n4 8.0005
R29893 _325_.A2.n11 _325_.A2.n8 6.8405
R29894 _325_.A2.n6 _325_.A2.t10 5.8405
R29895 _325_.A2.n5 _325_.A2.n3 5.3555
R29896 _325_.A2.n3 _325_.A2.n1 5.29866
R29897 _325_.A2.n3 _325_.A2 4.67135
R29898 _325_.A2 _325_.A2.t0 4.31594
R29899 _325_.A2.n8 _325_.A2.n5 3.6005
R29900 _325_.A2 _325_.A2.n12 0.211571
R29901 _325_.A2.n10 _325_.A2 0.148735
R29902 _325_.A2.n7 _325_.A2 0.0921364
R29903 _325_.A2.n1 _325_.A2 0.00997368
R29904 a_29828_24455.n0 a_29828_24455.t6 121.874
R29905 a_29828_24455.t6 a_29828_24455.t5 61.5152
R29906 a_29828_24455.n1 a_29828_24455.t4 52.378
R29907 a_29828_24455.n1 a_29828_24455.t7 17.7152
R29908 a_29828_24455.n3 a_29828_24455.t1 11.1158
R29909 a_29828_24455.n4 a_29828_24455.n0 9.95623
R29910 a_29828_24455.t0 a_29828_24455.n4 8.02846
R29911 a_29828_24455.n3 a_29828_24455.n2 8.0005
R29912 a_29828_24455.n0 a_29828_24455.t3 6.7165
R29913 a_29828_24455.n2 a_29828_24455.t2 6.023
R29914 a_29828_24455.n2 a_29828_24455.n1 1.33883
R29915 a_29828_24455.n4 a_29828_24455.n3 0.376152
R29916 a_15828_27208.n3 a_15828_27208.t7 121.874
R29917 a_15828_27208.t7 a_15828_27208.t4 61.5152
R29918 a_15828_27208.n0 a_15828_27208.t2 52.378
R29919 a_15828_27208.n0 a_15828_27208.t5 17.7882
R29920 a_15828_27208.n2 a_15828_27208.t1 11.1158
R29921 a_15828_27208.n4 a_15828_27208.n3 9.99927
R29922 a_15828_27208.n2 a_15828_27208.n1 8.0005
R29923 a_15828_27208.n3 a_15828_27208.t3 6.7165
R29924 a_15828_27208.n1 a_15828_27208.t6 5.96217
R29925 a_15828_27208.t0 a_15828_27208.n4 5.40498
R29926 a_15828_27208.n1 a_15828_27208.n0 1.33883
R29927 a_15828_27208.n4 a_15828_27208.n2 0.333109
R29928 _311_.A2.n6 _311_.A2.t7 27.9595
R29929 _311_.A2.n1 _311_.A2.t5 26.7915
R29930 _311_.A2.n4 _311_.A2.t4 19.1995
R29931 _311_.A2.n3 _311_.A2.t3 18.6885
R29932 _311_.A2.n10 _311_.A2.n9 15.6155
R29933 _311_.A2.n0 _311_.A2.t11 15.3305
R29934 _311_.A2.n0 _311_.A2.t8 15.0872
R29935 _311_.A2.n5 _311_.A2 14.5805
R29936 _311_.A2.n4 _311_.A2.t10 13.6637
R29937 _311_.A2.n3 _311_.A2.t6 11.9603
R29938 _311_.A2.n9 _311_.A2.n2 11.6012
R29939 _311_.A2.n8 _311_.A2.n7 10.8905
R29940 _311_.A2 _311_.A2.t1 8.52139
R29941 _311_.A2 _311_.A2.n0 8.15932
R29942 _311_.A2 _311_.A2.n4 8.1405
R29943 _311_.A2.n2 _311_.A2.n1 8.11425
R29944 _311_.A2.n7 _311_.A2.n6 8.0005
R29945 _311_.A2.n8 _311_.A2.n5 7.0205
R29946 _311_.A2.n1 _311_.A2.t2 6.37583
R29947 _311_.A2.n6 _311_.A2.t9 5.8405
R29948 _311_.A2.n10 _311_.A2 5.27874
R29949 _311_.A2.n11 _311_.A2.n10 4.703
R29950 _311_.A2.n5 _311_.A2 4.6405
R29951 _311_.A2 _311_.A2.n3 4.24542
R29952 _311_.A2.n11 _311_.A2.t0 4.09844
R29953 _311_.A2.n9 _311_.A2.n8 3.2405
R29954 _311_.A2 _311_.A2.n11 0.218
R29955 _311_.A2.n2 _311_.A2 0.103735
R29956 _311_.A2.n7 _311_.A2 0.0921364
R29957 uo_out[4].n6 uo_out[4] 16.1626
R29958 uo_out[4].n5 uo_out[4].n4 7.19999
R29959 uo_out[4].n8 uo_out[4].n1 6.36507
R29960 uo_out[4].n7 uo_out[4].n2 6.36507
R29961 uo_out[4].n5 uo_out[4].n3 6.30441
R29962 uo_out[4] uo_out[4].n10 3.81667
R29963 uo_out[4].n4 uo_out[4].t4 2.89962
R29964 uo_out[4].n4 uo_out[4].t11 2.89962
R29965 uo_out[4].n1 uo_out[4].t8 2.89962
R29966 uo_out[4].n1 uo_out[4].t2 2.89962
R29967 uo_out[4].n2 uo_out[4].t3 2.89962
R29968 uo_out[4].n2 uo_out[4].t9 2.89962
R29969 uo_out[4].n3 uo_out[4].t10 2.89962
R29970 uo_out[4].n3 uo_out[4].t5 2.89962
R29971 uo_out[4].n9 uo_out[4].n0 2.70811
R29972 uo_out[4].n10 uo_out[4].t1 2.06607
R29973 uo_out[4].n10 uo_out[4].t7 2.06607
R29974 uo_out[4].n0 uo_out[4].t6 2.06607
R29975 uo_out[4].n0 uo_out[4].t0 2.06607
R29976 uo_out[4].n9 uo_out[4].n8 1.50949
R29977 uo_out[4].n8 uo_out[4].n7 0.877022
R29978 uo_out[4].n7 uo_out[4].n6 0.815785
R29979 uo_out[4] uo_out[4].n9 0.267929
R29980 uo_out[4].n6 uo_out[4].n5 0.0192013
R29981 uio_out[4] uio_out[4].t1 8.3895
R29982 uio_out[4] uio_out[4].t0 4.3844
R29983 a_52400_25987.n0 a_52400_25987.t7 121.874
R29984 a_52400_25987.t7 a_52400_25987.t5 61.5152
R29985 a_52400_25987.n1 a_52400_25987.t6 52.378
R29986 a_52400_25987.n1 a_52400_25987.t2 17.7152
R29987 a_52400_25987.n3 a_52400_25987.t1 11.1158
R29988 a_52400_25987.n4 a_52400_25987.n0 9.95623
R29989 a_52400_25987.t0 a_52400_25987.n4 8.02846
R29990 a_52400_25987.n3 a_52400_25987.n2 8.0005
R29991 a_52400_25987.n0 a_52400_25987.t3 6.7165
R29992 a_52400_25987.n2 a_52400_25987.t4 6.023
R29993 a_52400_25987.n2 a_52400_25987.n1 1.33883
R29994 a_52400_25987.n4 a_52400_25987.n3 0.376152
R29995 a_28820_30344.n3 a_28820_30344.t4 121.874
R29996 a_28820_30344.t4 a_28820_30344.t5 61.5152
R29997 a_28820_30344.n0 a_28820_30344.t3 52.378
R29998 a_28820_30344.n0 a_28820_30344.t6 17.7882
R29999 a_28820_30344.n2 a_28820_30344.t1 11.1158
R30000 a_28820_30344.n4 a_28820_30344.n3 9.95623
R30001 a_28820_30344.t0 a_28820_30344.n4 8.02846
R30002 a_28820_30344.n2 a_28820_30344.n1 8.0005
R30003 a_28820_30344.n3 a_28820_30344.t2 6.7165
R30004 a_28820_30344.n1 a_28820_30344.t7 5.96217
R30005 a_28820_30344.n1 a_28820_30344.n0 1.33883
R30006 a_28820_30344.n4 a_28820_30344.n2 0.376152
R30007 rst_n.n1 rst_n.t1 28.7301
R30008 rst_n.n0 rst_n.t0 18.7615
R30009 rst_n.n2 rst_n 16.8044
R30010 rst_n.n0 rst_n.t2 13.4447
R30011 rst_n.n2 rst_n.n1 2.66717
R30012 rst_n.n1 rst_n.n0 1.01439
R30013 rst_n rst_n.n2 0.0312895
R30014 a_23892_27208.n3 a_23892_27208.t4 121.874
R30015 a_23892_27208.t4 a_23892_27208.t7 61.5152
R30016 a_23892_27208.n0 a_23892_27208.t5 52.378
R30017 a_23892_27208.n0 a_23892_27208.t3 17.7882
R30018 a_23892_27208.n2 a_23892_27208.t1 11.1158
R30019 a_23892_27208.n4 a_23892_27208.n3 9.95623
R30020 a_23892_27208.t0 a_23892_27208.n4 8.02846
R30021 a_23892_27208.n2 a_23892_27208.n1 8.0005
R30022 a_23892_27208.n3 a_23892_27208.t2 6.7165
R30023 a_23892_27208.n1 a_23892_27208.t6 5.96217
R30024 a_23892_27208.n1 a_23892_27208.n0 1.33883
R30025 a_23892_27208.n4 a_23892_27208.n2 0.376152
R30026 _288_.ZN.n8 _288_.ZN.t5 21.5355
R30027 _288_.ZN.n1 _288_.ZN.t6 21.5355
R30028 _288_.ZN.n5 _288_.ZN.n4 18.9805
R30029 _288_.ZN.n10 _288_.ZN.n9 18.9464
R30030 _288_.ZN.n4 _288_.ZN.t7 15.8172
R30031 _288_.ZN.n5 _288_.ZN.t10 15.8172
R30032 _288_.ZN.n8 _288_.ZN.t3 9.91633
R30033 _288_.ZN.n3 _288_.ZN.t9 9.91633
R30034 _288_.ZN.n6 _288_.ZN.t8 9.91633
R30035 _288_.ZN.n1 _288_.ZN.t4 9.91633
R30036 _288_.ZN.n2 _288_.ZN.n1 9.26624
R30037 _288_.ZN.n7 _288_.ZN.n6 8.0005
R30038 _288_.ZN.n3 _288_.ZN.n2 8.0005
R30039 _288_.ZN.n9 _288_.ZN.n8 8.0005
R30040 _288_.ZN.n10 _288_.ZN.n0 6.58318
R30041 _288_.ZN.n4 _288_.ZN.n3 5.23217
R30042 _288_.ZN.n6 _288_.ZN.n5 5.23217
R30043 _288_.ZN _288_.ZN.t0 4.34603
R30044 _288_.ZN.n0 _288_.ZN.t2 2.89962
R30045 _288_.ZN.n0 _288_.ZN.t1 2.89962
R30046 _288_.ZN _288_.ZN.n7 1.17906
R30047 _288_.ZN.n7 _288_.ZN.n2 0.425606
R30048 _288_.ZN _288_.ZN.n10 0.245128
R30049 _288_.ZN.n9 _288_.ZN 0.0177059
R30050 uio_out[3] uio_out[3].t0 8.31126
R30051 a_35316_29159.n0 a_35316_29159.t3 121.874
R30052 a_35316_29159.t3 a_35316_29159.t4 61.5152
R30053 a_35316_29159.n1 a_35316_29159.t2 52.378
R30054 a_35316_29159.n1 a_35316_29159.t7 17.7152
R30055 a_35316_29159.n3 a_35316_29159.t1 11.1158
R30056 a_35316_29159.n4 a_35316_29159.n0 9.95623
R30057 a_35316_29159.t0 a_35316_29159.n4 8.02846
R30058 a_35316_29159.n3 a_35316_29159.n2 8.0005
R30059 a_35316_29159.n0 a_35316_29159.t6 6.7165
R30060 a_35316_29159.n2 a_35316_29159.t5 6.023
R30061 a_35316_29159.n2 a_35316_29159.n1 1.33883
R30062 a_35316_29159.n4 a_35316_29159.n3 0.376152
R30063 ui_in[0].n1 ui_in[0].t0 28.7301
R30064 ui_in[0].n0 ui_in[0].t1 18.7615
R30065 ui_in[0].n2 ui_in[0] 15.5444
R30066 ui_in[0].n0 ui_in[0].t2 13.5055
R30067 ui_in[0].n2 ui_in[0].n1 2.66717
R30068 ui_in[0].n1 ui_in[0].n0 1.01439
R30069 ui_in[0] ui_in[0].n2 0.0312895
R30070 ui_in[4].n0 ui_in[4].t1 29.2005
R30071 ui_in[4].n1 ui_in[4] 16.5226
R30072 ui_in[4].n0 ui_in[4].t0 12.1428
R30073 ui_in[4].n1 ui_in[4].n0 8.07362
R30074 ui_in[4] ui_in[4].n1 0.1265
R30075 a_42484_18183.n0 a_42484_18183.t7 121.874
R30076 a_42484_18183.t7 a_42484_18183.t5 61.5152
R30077 a_42484_18183.n1 a_42484_18183.t4 52.378
R30078 a_42484_18183.n1 a_42484_18183.t2 17.7152
R30079 a_42484_18183.n3 a_42484_18183.t1 11.1158
R30080 a_42484_18183.n4 a_42484_18183.n0 9.95623
R30081 a_42484_18183.t0 a_42484_18183.n4 8.02846
R30082 a_42484_18183.n3 a_42484_18183.n2 8.0005
R30083 a_42484_18183.n0 a_42484_18183.t3 6.7165
R30084 a_42484_18183.n2 a_42484_18183.t6 6.023
R30085 a_42484_18183.n2 a_42484_18183.n1 1.33883
R30086 a_42484_18183.n4 a_42484_18183.n3 0.376152
R30087 a_41028_28776.n3 a_41028_28776.t5 121.874
R30088 a_41028_28776.t5 a_41028_28776.t4 61.5152
R30089 a_41028_28776.n0 a_41028_28776.t3 52.378
R30090 a_41028_28776.n0 a_41028_28776.t2 17.7882
R30091 a_41028_28776.n2 a_41028_28776.t1 11.1158
R30092 a_41028_28776.n4 a_41028_28776.n3 9.95623
R30093 a_41028_28776.t0 a_41028_28776.n4 8.02846
R30094 a_41028_28776.n2 a_41028_28776.n1 8.0005
R30095 a_41028_28776.n3 a_41028_28776.t7 6.7165
R30096 a_41028_28776.n1 a_41028_28776.t6 5.96217
R30097 a_41028_28776.n1 a_41028_28776.n0 1.33883
R30098 a_41028_28776.n4 a_41028_28776.n2 0.376152
R30099 uio_oe[3] uio_oe[3].t0 8.31126
R30100 _256_.A2.n0 _256_.A2.t3 19.7835
R30101 _256_.A2.n0 _256_.A2.t2 14.3085
R30102 _256_.A2.n1 _256_.A2.t1 8.92356
R30103 _256_.A2 _256_.A2.n0 8.0005
R30104 _256_.A2.n1 _256_.A2.t0 4.12916
R30105 _256_.A2 _256_.A2.n1 0.023
R30106 _268_.A2.n1 _268_.A2.t5 26.7915
R30107 _268_.A2.n0 _268_.A2.t6 16.0362
R30108 _268_.A2.n3 _268_.A2.t9 16.0118
R30109 _268_.A2.n5 _268_.A2.t8 15.3305
R30110 _268_.A2.n5 _268_.A2.t3 15.148
R30111 _268_.A2.n0 _268_.A2.t7 14.7465
R30112 _268_.A2.n2 _268_.A2 14.378
R30113 _268_.A2.n3 _268_.A2.t4 13.2622
R30114 _268_.A2.n7 _268_.A2.n6 12.4205
R30115 _268_.A2.n4 _268_.A2 10.9207
R30116 _268_.A2.n6 _268_.A2 9.68874
R30117 _268_.A2.n7 _268_.A2.t1 9.61569
R30118 _268_.A2.n2 _268_.A2 9.3605
R30119 _268_.A2 _268_.A2.n5 8.15932
R30120 _268_.A2 _268_.A2.n0 8.158
R30121 _268_.A2 _268_.A2.n1 8.13682
R30122 _268_.A2 _268_.A2.n3 8.13034
R30123 _268_.A2.n1 _268_.A2.t2 6.37583
R30124 _268_.A2 _268_.A2.t0 4.43672
R30125 _268_.A2.n6 _268_.A2.n4 1.9805
R30126 _268_.A2.n4 _268_.A2.n2 0.7205
R30127 _268_.A2 _268_.A2.n7 0.0859237
R30128 a_45456_30301.n3 a_45456_30301.t4 121.874
R30129 a_45456_30301.t4 a_45456_30301.t5 61.5152
R30130 a_45456_30301.n0 a_45456_30301.t7 52.378
R30131 a_45456_30301.n0 a_45456_30301.t6 17.7882
R30132 a_45456_30301.n2 a_45456_30301.t1 11.1158
R30133 a_45456_30301.n4 a_45456_30301.n3 9.95623
R30134 a_45456_30301.t0 a_45456_30301.n4 8.02846
R30135 a_45456_30301.n2 a_45456_30301.n1 8.0005
R30136 a_45456_30301.n3 a_45456_30301.t3 6.7165
R30137 a_45456_30301.n1 a_45456_30301.t2 5.96217
R30138 a_45456_30301.n1 a_45456_30301.n0 1.33883
R30139 a_45456_30301.n4 a_45456_30301.n2 0.376152
R30140 uio_oe[1] uio_oe[1].t0 8.31126
R30141 ena.n0 ena.t0 29.2005
R30142 ena.n0 ena.t1 12.1428
R30143 ena ena.n0 8.19963
R30144 uio_oe[2] uio_oe[2].t0 8.31126
R30145 uio_in[1].n0 uio_in[1].t0 19.7105
R30146 uio_in[1].n1 uio_in[1] 15.6533
R30147 uio_in[1].n0 uio_in[1].t1 13.3108
R30148 uio_in[1].n1 uio_in[1].n0 4.0005
R30149 uio_in[1] uio_in[1].n1 0.0737
R30150 uio_oe[6] uio_oe[6].t0 4.13855
R30151 uio_oe[4] uio_oe[4].t0 4.13855
R30152 uio_out[0] uio_out[0].t0 8.31126
R30153 uio_oe[7] uio_oe[7].t0 4.13855
R30154 uio_out[1] uio_out[1].t0 8.31126
R30155 ui_in[3].n0 ui_in[3].t0 29.2005
R30156 ui_in[3].n0 ui_in[3].t1 12.1428
R30157 ui_in[3] ui_in[3].n0 8.19963
R30158 uio_out[2] uio_out[2].t0 8.31126
C0 _260_.A1 a_41440_23208# 0.01383f
C1 a_4516_26724# a_4604_26680# 0.28563f
C2 _336_.A2 a_28552_25940# 0.01094f
C3 _474_.CLK a_48708_29816# 0.02156f
C4 a_37084_1159# a_37532_1159# 0.0131f
C5 a_67572_10664# a_68020_10664# 0.01328f
C6 _355_.B a_27328_25227# 0.05263f
C7 a_1468_20408# VPWR 0.29679f
C8 _371_.ZN a_28432_29535# 0.00156f
C9 _336_.A2 a_25884_24679# 0.00595f
C10 _304_.B _381_.Z 0.0403f
C11 _388_.B a_45508_31048# 0.00286f
C12 _452_.Q a_42982_21730# 0.00875f
C13 a_65756_2727# VPWR 0.31963f
C14 a_45820_12568# VPWR 0.29679f
C15 a_61748_16936# a_62196_16936# 0.01328f
C16 a_67012_2824# a_67100_1159# 0.0027f
C17 _284_.ZN a_41160_29083# 0.0175f
C18 a_4828_29383# a_4740_29480# 0.28563f
C19 a_41028_15368# a_41476_15368# 0.01328f
C20 a_34644_20072# VPWR 0.2434f
C21 _416_.A1 a_44864_27165# 0.01991f
C22 _250_.C a_61948_27815# 0.00101f
C23 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN 0.63209f
C24 a_66316_10567# VPWR 0.32291f
C25 a_43132_15271# a_43044_15368# 0.28563f
C26 a_27004_27815# a_26916_27912# 0.28563f
C27 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN 0.66543f
C28 a_65308_17272# a_65332_16936# 0.00172f
C29 a_28260_23208# VPWR 0.20595f
C30 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN a_65756_26247# 0.00412f
C31 _275_.A2 a_51457_29861# 0.02556f
C32 a_54444_19975# a_54892_19975# 0.01222f
C33 a_44476_15271# a_44924_15271# 0.0131f
C34 _336_.A2 a_28256_25597# 0.03141f
C35 a_16052_22020# a_16500_22020# 0.01328f
C36 a_57020_2727# a_56932_2824# 0.28563f
C37 a_63876_15748# VPWR 0.20595f
C38 _327_.Z a_40580_20072# 0.05783f
C39 a_1020_16839# a_1468_16839# 0.0131f
C40 a_55340_23544# clk 0.00613f
C41 a_22660_23208# a_22748_21543# 0.00151f
C42 _330_.A1 a_38852_25156# 0.00557f
C43 a_49600_30180# _324_.C 0.00134f
C44 a_7876_1256# VPWR 0.20968f
C45 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I 0.07209f
C46 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN a_61500_17272# 0.00576f
C47 a_2276_7908# VPWR 0.20634f
C48 a_26132_23588# a_25772_23544# 0.0869f
C49 a_22636_23544# a_23084_23544# 0.0131f
C50 _417_.A2 a_47552_19715# 0.00667f
C51 a_10452_31048# VPWR 0.21152f
C52 a_37892_1256# a_38340_1256# 0.01328f
C53 a_20980_25156# a_20620_25112# 0.08707f
C54 a_4068_4772# VPWR 0.2157f
C55 a_52876_13703# a_53236_13800# 0.08707f
C56 _251_.A1 a_62644_26724# 0.04979f
C57 a_66764_13703# a_67212_13703# 0.0131f
C58 _317_.A2 VPWR 1.42648f
C59 a_17148_2727# a_17596_2727# 0.0131f
C60 _424_.A2 a_52036_22504# 0.00207f
C61 _419_.A4 a_46352_22021# 0.0041f
C62 VPWR ui_in[1] 0.36276f
C63 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I 0.00124f
C64 a_39660_16839# a_40020_16936# 0.08707f
C65 a_46628_10664# a_46628_9476# 0.05841f
C66 a_66092_16839# VPWR 0.35504f
C67 a_34084_1636# VPWR 0.20902f
C68 _447_.Q _438_.ZN 0.44955f
C69 a_4068_1636# a_3708_1592# 0.08707f
C70 a_44028_27815# VPWR 0.32555f
C71 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I 0.00886f
C72 a_62756_27912# vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN 0.00141f
C73 a_2276_29860# a_2724_29860# 0.01328f
C74 a_4068_17316# a_4516_17316# 0.01328f
C75 a_2276_17316# a_1916_17272# 0.08717f
C76 _330_.A1 a_36016_20893# 0.00145f
C77 a_5052_11000# a_4940_10567# 0.02634f
C78 a_57044_23588# clk 0.00219f
C79 a_54108_11000# a_54556_11000# 0.01288f
C80 a_58052_11044# a_58140_11000# 0.28563f
C81 a_53012_16936# a_53460_16936# 0.01328f
C82 a_47388_1592# a_47972_1636# 0.01675f
C83 a_44500_25156# VPWR 0.00866f
C84 a_57492_17316# a_57132_17272# 0.0869f
C85 a_1380_20072# a_1380_18884# 0.05841f
C86 _294_.A2 _290_.ZN 0.3879f
C87 a_19948_26680# a_20396_26680# 0.01222f
C88 a_54892_26680# a_54780_26247# 0.02634f
C89 a_47252_18884# VPWR 0.00664f
C90 a_1828_25156# VPWR 0.20348f
C91 a_1468_27815# a_1828_27912# 0.08717f
C92 a_15692_27815# a_16140_27815# 0.0131f
C93 a_60656_29612# VPWR 0.00983f
C94 _381_.Z VPWR 1.14615f
C95 a_25012_20452# VPWR 0.20692f
C96 a_59484_12568# VPWR 0.31547f
C97 a_3172_15748# a_3260_15704# 0.28563f
C98 a_60212_25156# a_60416_25156# 0.03324f
C99 a_17956_2824# a_18404_2824# 0.01328f
C100 a_15580_29383# a_16164_29480# 0.01675f
C101 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_56236_24679# 0.00264f
C102 _350_.A2 _459_.CLK 0.13206f
C103 a_55452_21543# a_55364_21640# 0.28563f
C104 a_60180_10664# VPWR 0.20896f
C105 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I a_60180_14180# 0.03156f
C106 a_5388_7431# a_5300_7528# 0.28563f
C107 a_54108_15271# a_54468_15368# 0.08717f
C108 a_4156_8999# a_4068_9096# 0.28563f
C109 a_65756_4295# a_65668_4392# 0.28563f
C110 _324_.C _238_.I 0.08706f
C111 a_64860_5863# a_64772_5960# 0.28563f
C112 _362_.B _452_.CLK 0.3944f
C113 _294_.A2 a_37396_29860# 0.00304f
C114 a_51540_24776# VPWR 0.00636f
C115 a_33412_15368# VPWR 0.20644f
C116 a_51048_26680# a_51436_27208# 0.00334f
C117 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.00129f
C118 _474_.CLK vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN 0.03121f
C119 a_52920_22760# _281_.A1 0.00996f
C120 a_36860_15271# VPWR 0.32932f
C121 a_2276_14180# a_1916_14136# 0.08717f
C122 a_4068_14180# a_4516_14180# 0.01328f
C123 a_44038_21236# a_44270_21790# 0.00209f
C124 a_64748_23111# vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN 0.00161f
C125 a_32180_23588# a_31820_23544# 0.08663f
C126 a_30276_1256# VPWR 0.20348f
C127 a_65308_7431# VPWR 0.30378f
C128 _255_.ZN a_58340_29860# 0.00132f
C129 a_14004_31048# uio_oe[2] 0.0965f
C130 a_67100_4295# VPWR 0.29679f
C131 _260_.ZN a_42168_22504# 0.03405f
C132 a_58588_21543# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.05735f
C133 a_63852_13703# a_63764_13800# 0.28563f
C134 a_61412_26344# VPWR 0.2093f
C135 _346_.B a_22064_27912# 0.00116f
C136 a_38584_28292# a_38523_27967# 0.01684f
C137 _474_.CLK _402_.A1 0.77911f
C138 a_36548_17316# a_36524_16839# 0.00172f
C139 a_32604_17272# a_32604_16839# 0.05841f
C140 a_13452_30951# VPWR 0.32115f
C141 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN a_62844_27815# 0.02475f
C142 a_39300_31048# VPWR 0.01802f
C143 a_50860_16839# a_50772_16936# 0.28563f
C144 _358_.A3 a_32292_26344# 0.01996f
C145 a_63876_18504# VPWR 0.20348f
C146 a_2724_23208# a_2724_22020# 0.05841f
C147 _359_.B a_30795_29977# 0.0018f
C148 a_45620_16936# VPWR 0.20681f
C149 a_40220_1592# VPWR 0.33352f
C150 a_9532_1159# a_9892_1256# 0.08717f
C151 _452_.Q _304_.A1 2.26526f
C152 _260_.A2 _305_.A2 0.0864f
C153 a_2724_29480# a_3172_29480# 0.01328f
C154 a_10564_1636# a_11012_1636# 0.01328f
C155 _434_.ZN VPWR 1.00811f
C156 a_53772_12135# a_54220_12135# 0.01288f
C157 a_67772_12568# a_67660_12135# 0.02634f
C158 a_24876_23544# a_24988_23111# 0.02634f
C159 a_46984_23588# a_47412_23588# 0.00223f
C160 a_41440_28363# a_42320_28777# 0.00306f
C161 a_32068_17316# a_31708_17272# 0.08707f
C162 a_61412_11044# a_61500_11000# 0.28563f
C163 a_51644_11000# a_51532_10567# 0.02634f
C164 a_10340_2824# VPWR 0.21189f
C165 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN 0.00432f
C166 _248_.B1 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.0828f
C167 a_54692_1636# a_54332_1592# 0.08707f
C168 _393_.A3 a_47700_28292# 0.00246f
C169 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I a_58388_20452# 0.01061f
C170 _397_.A2 a_47525_29480# 0.00603f
C171 _365_.ZN a_34084_28776# 0.0227f
C172 a_11100_29816# uio_oe[4] 0.00114f
C173 a_36996_26724# VPWR 0.20348f
C174 a_16140_24679# a_16588_24679# 0.0131f
C175 _416_.A2 a_46476_20937# 0.00141f
C176 a_59484_1159# a_59932_1159# 0.0131f
C177 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN a_53460_18504# 0.00168f
C178 a_54444_18407# a_54356_18504# 0.28563f
C179 a_66764_20408# a_67212_20408# 0.012f
C180 a_63876_15368# VPWR 0.20897f
C181 a_57492_18504# VPWR 0.21569f
C182 a_52640_29860# VPWR 0.01437f
C183 a_20172_25112# VPWR 0.31547f
C184 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.06757f
C185 a_32964_15748# a_33052_15704# 0.28563f
C186 a_36548_15748# a_36996_15748# 0.01328f
C187 _427_.ZN a_53796_20452# 0.00422f
C188 a_46268_12135# VPWR 0.29679f
C189 _359_.ZN a_35204_26344# 0.00469f
C190 a_20956_2727# a_21092_1636# 0.00154f
C191 _324_.C hold2.I 0.03387f
C192 a_46628_18504# a_46492_17272# 0.00154f
C193 a_50324_18504# a_50436_17316# 0.02666f
C194 a_36772_23208# VPWR 0.12511f
C195 a_60416_25156# VPWR 0.00966f
C196 _251_.A1 a_63952_29480# 0.14256f
C197 uo_out[5] uo_out[6] 0.06365f
C198 a_38304_20072# VPWR 0.01426f
C199 _383_.ZN _381_.Z 0.08848f
C200 _452_.CLK a_43020_16839# 0.01498f
C201 _384_.ZN _395_.A1 0.39915f
C202 a_4156_15704# VPWR 0.30552f
C203 _250_.C a_62308_27912# 0.00134f
C204 _381_.Z a_50068_27508# 0.02379f
C205 a_55812_15368# VPWR 0.20348f
C206 _301_.A1 a_38529_22804# 0.00482f
C207 _359_.B a_34155_25273# 0.00833f
C208 a_64300_23544# vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN 0.00227f
C209 a_26132_22020# a_26220_21976# 0.28563f
C210 _350_.A2 _371_.A3 0.05264f
C211 a_54804_24776# clk 0.0155f
C212 _247_.B a_59172_27912# 0.01027f
C213 a_23084_29383# _345_.A2 0.00212f
C214 a_47948_16839# a_48396_16839# 0.01288f
C215 a_46628_14180# a_46268_14136# 0.08707f
C216 a_40556_16839# VPWR 0.31208f
C217 a_52676_1256# VPWR 0.20348f
C218 a_37196_23544# a_37644_23544# 0.01255f
C219 a_60292_1256# a_60740_1256# 0.01328f
C220 _397_.A2 a_51084_28248# 0.00511f
C221 _274_.A3 VPWR 0.60718f
C222 a_57940_17316# VPWR 0.21952f
C223 a_60628_13800# a_61076_13800# 0.01328f
C224 a_39548_2727# a_39996_2727# 0.0131f
C225 _474_.CLK a_53996_25112# 0.04103f
C226 _459_.CLK a_29804_23544# 0.00127f
C227 _251_.A1 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN 0.0375f
C228 a_31260_17272# VPWR 0.29679f
C229 a_20420_23208# a_20532_22020# 0.02666f
C230 _402_.A1 _265_.ZN 0.07989f
C231 _349_.A4 VPWR 1.90478f
C232 a_36016_20893# a_35723_20569# 0.49319f
C233 a_20956_1159# a_20868_1256# 0.28563f
C234 a_53884_1592# VPWR 0.32982f
C235 _408_.ZN _407_.ZN 0.63647f
C236 a_51084_12135# a_50996_12232# 0.28563f
C237 a_12356_29860# a_12444_29816# 0.28563f
C238 _355_.C a_20191_29611# 0.00358f
C239 _252_.ZN a_60852_28292# 0.01349f
C240 _317_.A2 a_36636_21543# 0.00396f
C241 a_39236_17316# a_40040_17675# 0.00302f
C242 a_5300_15368# a_5388_13703# 0.0027f
C243 _336_.A2 a_27476_23588# 0.00702f
C244 a_58588_11000# a_58476_10567# 0.02634f
C245 a_1020_10567# a_1468_10567# 0.0131f
C246 a_32740_2824# VPWR 0.20348f
C247 a_57604_1636# a_57692_1592# 0.28563f
C248 a_61188_1636# a_61636_1636# 0.01328f
C249 a_30388_28776# VPWR 0.02697f
C250 _281_.ZN clk 0.26811f
C251 _384_.A3 _427_.B2 0.20344f
C252 _383_.A2 VPWR 0.64982f
C253 a_27004_23111# a_27452_23111# 0.01288f
C254 a_14796_23111# a_15156_23208# 0.08717f
C255 a_18716_24679# a_19076_24776# 0.08707f
C256 _444_.D a_36300_23544# 0.00277f
C257 a_4516_9476# VPWR 0.20862f
C258 _350_.A2 uo_out[7] 0.05713f
C259 a_45820_14136# VPWR 0.29679f
C260 a_10788_2824# a_10876_1159# 0.0027f
C261 a_51332_2824# a_51196_1592# 0.00154f
C262 a_55140_2824# a_55140_1636# 0.05841f
C263 a_31260_18407# a_31172_18504# 0.28563f
C264 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I VPWR 0.96949f
C265 a_3620_31048# a_3620_29860# 0.05841f
C266 a_68108_12135# VPWR 0.35526f
C267 _304_.B _324_.C 2.01097f
C268 _467_.D VPWR 0.58126f
C269 _373_.A2 a_28054_30196# 0.06366f
C270 a_53704_23219# a_54040_22366# 0.00983f
C271 a_40356_2824# a_40804_2824# 0.01328f
C272 _304_.B a_40220_20408# 0.00426f
C273 a_4068_24776# VPWR 0.22146f
C274 vgaringosc.workerclkbuff_notouch_.I _397_.A2 0.04722f
C275 a_20003_29611# _375_.Z 0.18628f
C276 a_59955_30600# _237_.A1 0.26253f
C277 _334_.A1 _459_.CLK 0.09506f
C278 a_28708_21640# a_28820_20452# 0.02666f
C279 a_2364_19975# a_2724_20072# 0.08717f
C280 vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I clk 0.28668f
C281 a_43044_15748# VPWR 0.21514f
C282 a_43008_26795# a_44571_26841# 0.41635f
C283 a_41099_26841# a_41384_26841# 0.00277f
C284 a_45732_9476# a_45372_9432# 0.08717f
C285 a_47076_9476# a_47524_9476# 0.01328f
C286 a_32180_22020# a_31820_21976# 0.08663f
C287 a_53124_14180# a_53572_14180# 0.01328f
C288 a_40436_26841# VPWR 0.00246f
C289 _459_.CLK _457_.D 0.01122f
C290 a_36960_27912# a_38523_27967# 0.41635f
C291 _443_.D a_37516_27599# 0.26504f
C292 _230_.I ui_in[0] 0.00366f
C293 a_30388_25156# VPWR 0.23063f
C294 a_1828_12612# a_1916_12568# 0.28563f
C295 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I a_66228_20452# 0.05859f
C296 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_64884_26724# 0.01986f
C297 a_51756_18407# a_51780_17316# 0.0016f
C298 _459_.CLK _454_.Q 0.46771f
C299 a_34304_24029# a_33932_24073# 0.10745f
C300 _256_.A2 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN 0.01826f
C301 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I _248_.B1 0.0292f
C302 _284_.ZN a_40038_28720# 0.08269f
C303 _402_.A1 _398_.C 0.69008f
C304 _251_.A1 a_65084_30951# 0.00464f
C305 _252_.ZN _238_.I 0.03154f
C306 _279_.Z clkbuf_1_0__f_clk.I 0.07935f
C307 a_27364_23208# a_27476_22020# 0.02666f
C308 a_50884_17316# VPWR 0.21315f
C309 a_23556_23208# a_23532_21976# 0.0016f
C310 a_67684_1636# VPWR 0.21497f
C311 a_57828_25156# VPWR 0.20103f
C312 a_31932_1159# a_32292_1256# 0.08717f
C313 a_21652_31048# uio_out[4] 0.00506f
C314 a_47524_12232# a_47972_12232# 0.01328f
C315 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN a_64100_27912# 0.02582f
C316 a_61612_12135# a_61972_12232# 0.08707f
C317 a_59036_12568# a_58948_11044# 0.00151f
C318 _378_.I a_21652_29480# 0.19396f
C319 a_16700_1592# a_17148_1592# 0.01288f
C320 a_20644_1636# a_20732_1592# 0.28563f
C321 a_16028_29816# _459_.CLK 0.0028f
C322 a_23644_21543# VPWR 0.31547f
C323 a_32292_26344# a_31803_24831# 0.00139f
C324 a_22996_28292# _345_.A2 0.00794f
C325 a_55140_2824# VPWR 0.20348f
C326 a_55452_11000# a_55476_10664# 0.00172f
C327 a_41028_1636# a_40892_1159# 0.00168f
C328 a_1828_2824# a_1828_1636# 0.05841f
C329 _470_.D _284_.A2 0.14042f
C330 _411_.A2 a_49764_26724# 0.01153f
C331 _470_.Q a_45128_26031# 0.00159f
C332 a_25884_23111# a_25796_23208# 0.28563f
C333 a_20868_24776# a_21316_24776# 0.01328f
C334 a_54244_9476# VPWR 0.20692f
C335 a_61412_14180# VPWR 0.20897f
C336 _452_.CLK a_34308_24776# 0.01014f
C337 _274_.ZN vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.00226f
C338 _474_.Q _324_.B 0.24712f
C339 _397_.A1 _384_.ZN 0.171f
C340 _383_.A2 _383_.ZN 0.21489f
C341 _324_.C VPWR 5.40483f
C342 a_61972_12232# VPWR 0.20622f
C343 _335_.ZN _223_.ZN 1.76736f
C344 a_42684_15704# a_43132_15704# 0.01288f
C345 a_40220_20408# VPWR 0.29679f
C346 a_64996_31048# VPWR 0.17093f
C347 _474_.CLK _424_.B1 0.06624f
C348 a_66116_18884# a_66092_18407# 0.00172f
C349 _288_.ZN a_37291_29535# 0.01047f
C350 a_67348_20072# VPWR 0.20595f
C351 _319_.A3 _319_.ZN 0.04234f
C352 a_11772_2727# a_12356_2824# 0.01675f
C353 a_59332_29816# _324_.C 0.23981f
C354 _452_.Q a_39684_20072# 0.01108f
C355 a_24864_29931# _340_.ZN 0.00307f
C356 a_63964_19975# a_64412_19975# 0.0131f
C357 a_49180_15704# VPWR 0.3009f
C358 _416_.ZN VPWR 0.43823f
C359 a_17732_31048# uio_out[7] 0.00733f
C360 _495_.I _265_.ZN 0.01037f
C361 a_46940_17272# a_46852_15748# 0.00151f
C362 a_2276_20452# a_2724_20452# 0.01328f
C363 a_22636_25112# a_22548_23588# 0.00151f
C364 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN VPWR 0.79686f
C365 _324_.B a_43892_20072# 0.00368f
C366 _402_.A1 a_39884_27815# 0.00714f
C367 _474_.CLK _386_.ZN 0.00117f
C368 a_46180_12612# a_46268_12568# 0.28563f
C369 a_49764_12612# a_50212_12612# 0.01328f
C370 a_61948_2727# a_62396_2727# 0.0131f
C371 _424_.A2 _412_.ZN 0.40125f
C372 _284_.A2 _412_.B2 0.00196f
C373 a_67100_18840# a_67012_17316# 0.00151f
C374 a_43356_1159# a_43268_1256# 0.28563f
C375 a_62396_12568# a_62308_11044# 0.00151f
C376 a_65220_7528# a_65220_6340# 0.05841f
C377 a_64324_9096# a_64324_7908# 0.05841f
C378 a_30724_20072# a_31172_20072# 0.01328f
C379 a_18044_1159# VPWR 0.30075f
C380 a_66116_5960# a_66116_4772# 0.05841f
C381 a_67012_4392# a_67012_3204# 0.05841f
C382 _402_.A1 _393_.A3 0.03511f
C383 a_20868_21640# VPWR 0.20641f
C384 a_35740_26247# a_36188_26247# 0.01255f
C385 a_50524_17272# a_50972_17272# 0.01288f
C386 _452_.CLK a_39684_26344# 0.00546f
C387 a_48508_10567# a_49204_10664# 0.01227f
C388 a_3260_1159# a_3708_1159# 0.0131f
C389 a_62508_10567# a_62956_10567# 0.01288f
C390 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN a_63852_23544# 0.00305f
C391 _330_.A1 _325_.A2 0.61658f
C392 _330_.A1 a_36524_18407# 0.02186f
C393 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN 0.12881f
C394 a_24452_23208# a_24900_23208# 0.01328f
C395 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN a_61724_18407# 0.00105f
C396 _304_.B a_40332_21543# 0.0125f
C397 a_65220_9476# VPWR 0.21249f
C398 a_51428_20452# VPWR 0.00975f
C399 a_18292_23588# VPWR 0.21304f
C400 a_67908_6340# VPWR 0.21437f
C401 a_54804_20072# VPWR 0.20622f
C402 a_19164_21543# a_19076_21640# 0.28563f
C403 _251_.A1 ui_in[4] 0.01253f
C404 a_31036_21543# a_31484_21543# 0.01288f
C405 a_65756_3160# VPWR 0.31505f
C406 a_48060_13703# VPWR 0.29679f
C407 a_4740_29480# a_4604_28248# 0.00154f
C408 a_67012_2824# a_66876_1592# 0.00154f
C409 _455_.Q a_23920_27555# 0.02122f
C410 _334_.A1 uo_out[7] 2.0048f
C411 a_18180_31048# _459_.CLK 0.00192f
C412 _459_.CLK a_23284_26724# 0.00112f
C413 a_49988_15748# a_49628_15704# 0.08707f
C414 _316_.ZN _316_.A3 0.04078f
C415 a_51108_11044# VPWR 0.20627f
C416 a_12892_29816# a_12892_29383# 0.05841f
C417 a_62756_2824# a_63204_2824# 0.01328f
C418 _304_.ZN a_42252_20936# 1.5247f
C419 a_62308_27912# a_62284_26680# 0.0016f
C420 a_56964_26724# a_58140_26680# 0.00689f
C421 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I 0.00479f
C422 _451_.Q _438_.ZN 0.05896f
C423 _459_.CLK a_41140_27912# 0.0026f
C424 a_1828_26344# VPWR 0.20348f
C425 a_54692_26344# VPWR 0.13408f
C426 a_42908_30951# vgaringosc.workerclkbuff_notouch_.I 0.00116f
C427 a_23196_2727# a_23108_2824# 0.28563f
C428 a_53884_20408# VPWR 0.32236f
C429 _267_.A2 a_53616_29480# 0.00162f
C430 _384_.A1 a_54892_23544# 0.00447f
C431 _252_.ZN a_60212_25156# 0.00125f
C432 _438_.A2 a_37472_24419# 0.18149f
C433 _324_.C a_50068_27508# 0.0023f
C434 _223_.I _352_.A2 0.0171f
C435 _474_.CLK a_52676_17316# 0.002f
C436 a_5052_9432# a_4940_8999# 0.02634f
C437 a_56124_9432# a_56796_9432# 0.00544f
C438 a_58052_9476# a_58500_9476# 0.01328f
C439 a_3172_28292# VPWR 0.20993f
C440 a_4068_1256# a_4740_1256# 0.00347f
C441 a_4740_31048# a_5188_31048# 0.01328f
C442 a_61500_14136# a_61948_14136# 0.01288f
C443 a_1380_3204# a_1828_3204# 0.01328f
C444 a_65444_14180# a_65084_14136# 0.08707f
C445 a_16052_20452# a_16140_20408# 0.28563f
C446 a_34080_22461# a_33708_22505# 0.10745f
C447 a_17820_30951# uio_out[7] 0.00877f
C448 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I 0.02306f
C449 _450_.D _331_.ZN 0.00152f
C450 a_21628_1592# a_21764_1256# 0.00168f
C451 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I 0.63145f
C452 a_51892_13800# a_51980_12135# 0.00151f
C453 _397_.A2 a_48292_26369# 0.0048f
C454 a_20379_29977# a_20624_30345# 0.00232f
C455 _459_.CLK a_18816_29931# 0.00136f
C456 a_40444_1159# VPWR 0.3289f
C457 a_54332_1159# a_54692_1256# 0.08717f
C458 a_1828_11044# a_2276_11044# 0.01328f
C459 a_30364_1592# a_30812_1592# 0.01288f
C460 a_62284_16839# a_62732_16839# 0.0131f
C461 a_47776_20893# a_47483_20569# 0.49319f
C462 _419_.Z a_51108_21640# 0.01574f
C463 _229_.I a_60068_27912# 0.00254f
C464 a_59820_10567# a_59732_10664# 0.28563f
C465 _304_.B _281_.A1 0.11234f
C466 a_41564_24679# _226_.ZN 0.00226f
C467 a_2276_18504# a_2276_17316# 0.05841f
C468 _304_.B a_41996_28777# 0.00657f
C469 a_19188_22020# VPWR 0.22891f
C470 a_40332_21543# VPWR 0.31247f
C471 a_42340_28409# VPWR 0.00258f
C472 a_25772_23544# VPWR 0.31768f
C473 a_20508_2727# VPWR 0.31143f
C474 a_54192_22851# VPWR 0.3991f
C475 a_2276_13800# VPWR 0.20634f
C476 a_2812_18840# a_3260_18840# 0.0131f
C477 _460_.Q uo_out[6] 0.00689f
C478 a_29692_21543# a_30052_21640# 0.08707f
C479 _470_.Q a_48580_27508# 0.0041f
C480 a_5412_29860# VPWR 0.2085f
C481 a_63068_15704# a_63068_15271# 0.05841f
C482 a_57244_11000# VPWR 0.32088f
C483 a_40220_26247# a_40580_26344# 0.0869f
C484 vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I 0.01821f
C485 a_18268_30951# _459_.CLK 0.00208f
C486 _424_.B1 _398_.C 0.08141f
C487 _355_.C a_22560_30288# 0.00202f
C488 _370_.B a_30388_28776# 0.02522f
C489 a_67908_15748# a_67996_15704# 0.28563f
C490 _432_.ZN _325_.A1 0.48086f
C491 a_23627_27967# a_23912_27967# 0.00277f
C492 _363_.Z a_34586_27912# 0.00128f
C493 a_19948_27815# VPWR 0.3179f
C494 _474_.CLK a_53212_27815# 0.00744f
C495 a_61612_23111# a_61972_23208# 0.08717f
C496 a_34172_2727# a_34532_2824# 0.08717f
C497 _474_.Q a_50732_23233# 0.00179f
C498 _244_.Z vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN 0.00387f
C499 _397_.A4 a_47636_23588# 0.00694f
C500 a_64660_23588# a_65108_23588# 0.01328f
C501 a_43232_29480# a_44112_29167# 0.00306f
C502 a_49896_18909# a_50384_19204# 0.8399f
C503 a_53348_18884# a_52228_19368# 0.07589f
C504 a_49492_18840# a_49888_19369# 0.00232f
C505 _276_.A2 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN 0.01284f
C506 _251_.A1 a_59172_26724# 0.00116f
C507 a_63652_9476# a_63740_9432# 0.28563f
C508 _448_.Q a_38876_19975# 0.01649f
C509 a_54192_22851# a_54108_21543# 0.00144f
C510 _223_.I a_30912_27508# 0.0011f
C511 _300_.ZN _325_.A2 0.0019f
C512 a_1468_3160# a_1468_2727# 0.05841f
C513 a_64772_3204# a_64412_3160# 0.08717f
C514 _330_.A1 a_40244_18180# 0.02273f
C515 a_21292_20408# a_21740_20408# 0.0131f
C516 _252_.ZN VPWR 0.68794f
C517 a_45920_20523# a_47552_19715# 0.00205f
C518 a_7180_30951# a_7092_31048# 0.28563f
C519 _412_.ZN a_53716_26399# 0.00165f
C520 _365_.ZN a_36100_26724# 0.00163f
C521 a_13700_1636# VPWR 0.20348f
C522 a_55900_12568# a_56348_12568# 0.01288f
C523 a_59844_12612# a_59932_12568# 0.28563f
C524 a_52024_20083# a_53436_19759# 0.00393f
C525 a_20672_30301# uio_out[5] 0.82533f
C526 a_11100_29816# a_11236_29480# 0.00168f
C527 a_62844_1159# VPWR 0.3289f
C528 _350_.A2 _340_.A2 0.04081f
C529 a_65756_1159# a_65668_1256# 0.28563f
C530 a_2364_19975# VPWR 0.30029f
C531 a_60180_12232# a_60292_11044# 0.02666f
C532 a_56372_12232# a_56348_11000# 0.0016f
C533 a_37668_1636# a_37308_1592# 0.08707f
C534 a_3708_18407# VPWR 0.33374f
C535 _305_.A2 a_44500_22020# 0.00909f
C536 _311_.Z _317_.A2 0.01949f
C537 a_43940_27912# _330_.A1 0.00883f
C538 _345_.A2 a_22996_25156# 0.00193f
C539 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.00859f
C540 hold2.I a_44028_25156# 0.00249f
C541 _437_.A1 _430_.ZN 0.25319f
C542 _281_.A1 VPWR 1.35346f
C543 a_21396_26399# VPWR 0.00246f
C544 a_56372_10664# a_57044_10664# 0.00347f
C545 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN 0.00398f
C546 a_41996_28777# VPWR 0.42174f
C547 a_35988_18504# a_36100_17316# 0.02666f
C548 a_25660_1159# a_26108_1159# 0.0131f
C549 _350_.A2 _459_.Q 0.09789f
C550 a_18628_24776# a_18716_23111# 0.00151f
C551 a_25324_21976# VPWR 0.31533f
C552 a_53996_25112# a_53996_24679# 0.05841f
C553 a_18400_28733# VPWR 0.19184f
C554 _324_.C a_44744_26355# 0.0372f
C555 _452_.CLK a_32380_23111# 0.01311f
C556 _304_.ZN a_42154_21236# 0.04748f
C557 a_28260_21640# a_28708_21640# 0.01328f
C558 a_42908_2727# VPWR 0.33374f
C559 a_55588_2824# a_55676_1159# 0.0027f
C560 a_63764_13800# VPWR 0.20622f
C561 a_3708_26247# a_3620_26344# 0.28563f
C562 a_45396_22020# VPWR 0.02076f
C563 a_38472_30169# VPWR 0.99997f
C564 _474_.CLK _386_.A4 0.0059f
C565 _474_.CLK vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN 0.01479f
C566 a_4852_15368# a_5300_15368# 0.01328f
C567 _438_.A2 a_39669_21236# 0.00503f
C568 a_11548_29816# VPWR 0.37751f
C569 a_66452_16936# a_66564_15748# 0.02666f
C570 a_4156_10567# VPWR 0.3269f
C571 a_39796_22504# a_40780_21543# 0.00196f
C572 a_56124_2727# a_56260_1636# 0.00154f
C573 a_49112_29885# _383_.A2 0.00178f
C574 _443_.D a_37840_27599# 0.00106f
C575 _452_.CLK a_43888_19204# 0.00524f
C576 a_31708_15271# a_31620_15368# 0.28563f
C577 a_30140_23111# VPWR 0.33016f
C578 a_33052_15271# a_33500_15271# 0.0131f
C579 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN a_61276_15271# 0.00106f
C580 _229_.I a_62279_28293# 0.00199f
C581 a_59260_26680# a_59620_27208# 0.06541f
C582 _260_.A1 a_42084_24072# 0.00225f
C583 a_45596_2727# a_45508_2824# 0.28563f
C584 a_65668_17316# a_66116_17316# 0.01328f
C585 _452_.Q a_38644_19368# 0.00125f
C586 a_61500_17272# a_62172_17272# 0.00544f
C587 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN 0.02058f
C588 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I 0.01226f
C589 a_38852_18884# VPWR 0.01105f
C590 a_67436_16839# a_67796_16936# 0.08663f
C591 a_61500_26247# VPWR 0.33016f
C592 _459_.CLK _370_.ZN 0.03473f
C593 a_17932_23544# a_18380_23544# 0.01288f
C594 a_21876_23588# a_21964_23544# 0.28563f
C595 a_1916_8999# a_2364_8999# 0.0131f
C596 a_66204_7864# a_66204_7431# 0.05841f
C597 _474_.CLK a_53796_20452# 0.00377f
C598 a_2812_7431# a_3260_7431# 0.0131f
C599 a_3708_5863# a_4156_5863# 0.0131f
C600 _355_.C a_25884_27815# 0.01067f
C601 a_67100_6296# a_67100_5863# 0.05841f
C602 a_26468_1256# a_26916_1256# 0.01328f
C603 a_4940_4295# a_5388_4295# 0.01222f
C604 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I 0.00585f
C605 a_1916_13703# a_2276_13800# 0.08717f
C606 a_27028_20452# a_27116_20408# 0.28563f
C607 a_55564_13703# a_56012_13703# 0.01288f
C608 a_5724_2727# a_6172_2727# 0.0131f
C609 a_37780_16936# a_37756_15271# 0.00134f
C610 a_43736_25896# _435_.A3 0.00436f
C611 _274_.A2 a_56804_30344# 0.00592f
C612 _319_.A3 a_37360_19325# 0.00112f
C613 a_65756_26247# vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN 0.00383f
C614 a_37556_23588# VPWR 0.21206f
C615 a_3260_16839# a_3620_16936# 0.08717f
C616 a_19836_1592# VPWR 0.33243f
C617 a_63204_12612# a_63292_12568# 0.28563f
C618 a_1020_23544# a_1020_23111# 0.05841f
C619 a_9084_30951# a_9635_30644# 0.03643f
C620 _325_.A1 a_41804_19376# 0.00384f
C621 _325_.B _325_.ZN 0.01103f
C622 _223_.I _223_.ZN 0.63741f
C623 a_47271_21640# VPWR 0.50298f
C624 _267_.A1 _274_.A2 0.01608f
C625 a_66428_15271# a_66340_15368# 0.28563f
C626 a_50748_11000# a_51196_11000# 0.01288f
C627 a_41812_16936# a_42484_16936# 0.00347f
C628 a_67124_12232# a_67236_11044# 0.02666f
C629 a_40580_1636# a_40668_1592# 0.28563f
C630 a_44164_1636# a_44612_1636# 0.01328f
C631 _441_.B _301_.A1 0.00612f
C632 _386_.ZN _393_.A3 0.02391f
C633 _384_.ZN _389_.ZN 0.00327f
C634 _474_.CLK a_57020_23111# 0.00225f
C635 _304_.B a_44028_25156# 0.00352f
C636 _260_.A1 a_41216_23208# 0.01303f
C637 VPWR uio_in[3] 0.00114f
C638 a_4516_26724# a_4156_26680# 0.08674f
C639 a_1916_26680# a_2364_26680# 0.0131f
C640 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _416_.A1 0.12489f
C641 _395_.A2 a_50732_23233# 0.0162f
C642 _260_.A1 _325_.A1 0.81201f
C643 _294_.ZN _288_.ZN 0.00155f
C644 _243_.B2 a_58020_27508# 0.41657f
C645 _336_.A2 a_25436_24679# 0.0028f
C646 a_1020_20408# VPWR 0.30073f
C647 _397_.A1 a_51576_25896# 0.19571f
C648 a_65084_2727# VPWR 0.36385f
C649 _388_.B a_45060_31048# 0.00691f
C650 a_45372_12568# VPWR 0.30073f
C651 a_6620_29383# uio_oe[7] 0.00106f
C652 a_18628_26344# a_19076_26344# 0.01328f
C653 _452_.Q a_42778_21812# 0.11261f
C654 a_6620_2727# a_6756_1636# 0.00154f
C655 a_6532_2824# a_6980_2824# 0.01328f
C656 a_4156_29383# a_4740_29480# 0.01675f
C657 a_35008_27533# a_35140_26680# 0.00115f
C658 a_33860_20072# VPWR 0.21375f
C659 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I 0.00146f
C660 a_62420_22020# vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I 0.00466f
C661 a_1020_28248# a_1020_27815# 0.05841f
C662 a_61076_20452# a_61524_20452# 0.01328f
C663 a_26556_27815# a_26916_27912# 0.08674f
C664 a_65868_10567# VPWR 0.34668f
C665 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN a_61724_18407# 0.00499f
C666 a_42684_15271# a_43044_15368# 0.08717f
C667 a_30924_21976# a_31036_21543# 0.02634f
C668 a_37532_21543# a_37444_21640# 0.28563f
C669 a_27812_23208# VPWR 0.20595f
C670 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN a_64860_26247# 0.01912f
C671 a_41776_18504# _452_.D 0.00621f
C672 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN ui_in[1] 0.01609f
C673 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I a_61300_15748# 0.00211f
C674 _474_.D a_51220_18504# 0.00172f
C675 a_15156_28292# a_15604_28292# 0.01328f
C676 a_56572_2727# a_56932_2824# 0.08717f
C677 vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I 0.00725f
C678 a_40668_19975# a_40580_20072# 0.28563f
C679 a_54892_23544# clk 0.00613f
C680 a_63428_15748# VPWR 0.20595f
C681 a_60964_26344# a_60212_25156# 0.02619f
C682 _311_.Z a_36772_23208# 0.00646f
C683 a_33860_16936# a_33860_15748# 0.05841f
C684 _330_.A1 a_38628_25156# 0.00265f
C685 a_52564_18504# a_53012_18504# 0.01328f
C686 a_40244_18180# a_40040_17675# 0.00385f
C687 a_7428_1256# VPWR 0.20348f
C688 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN a_58924_17272# 0.0367f
C689 a_1828_7908# VPWR 0.20348f
C690 a_25684_23588# a_25772_23544# 0.28563f
C691 _417_.A2 a_47259_20127# 0.00104f
C692 a_10004_31048# VPWR 0.22654f
C693 a_16588_25112# a_17036_25112# 0.01288f
C694 a_3620_4772# VPWR 0.22347f
C695 a_20532_25156# a_20620_25112# 0.28563f
C696 a_30724_26020# _459_.D 0.00127f
C697 _324_.C _260_.ZN 0.00147f
C698 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I 0.65977f
C699 a_52920_22760# a_53704_23219# 0.02307f
C700 a_36148_21976# VPWR 0.81688f
C701 a_52876_13703# a_52788_13800# 0.28563f
C702 _251_.A1 a_62196_26724# 0.00446f
C703 a_32268_20408# a_32716_20408# 0.0131f
C704 a_37892_26344# _444_.D 0.00492f
C705 a_26108_30951# a_26556_30951# 0.01222f
C706 a_39660_16839# a_39572_16936# 0.28563f
C707 _355_.C _358_.A2 0.23834f
C708 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN 0.03547f
C709 _246_.B2 _247_.B 0.29777f
C710 _256_.A2 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN 0.08073f
C711 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I a_65072_29860# 0.03484f
C712 _251_.A1 a_59397_26344# 0.08384f
C713 a_65420_16839# VPWR 0.35266f
C714 a_33636_1636# VPWR 0.20713f
C715 a_2812_12135# a_3260_12135# 0.0131f
C716 a_60380_12568# a_60268_12135# 0.02634f
C717 a_3620_1636# a_3708_1592# 0.28563f
C718 a_7204_1636# a_7652_1636# 0.01328f
C719 a_17036_23544# a_17036_23111# 0.05841f
C720 _460_.Q a_35740_25112# 0.00415f
C721 a_43580_27815# VPWR 0.31205f
C722 a_20980_23588# a_20956_23111# 0.00172f
C723 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I VPWR 0.7305f
C724 a_45012_29816# a_45416_29885# 0.41635f
C725 _330_.A1 a_34716_20937# 0.0273f
C726 a_1828_17316# a_1916_17272# 0.28563f
C727 a_56596_23588# clk 0.00657f
C728 a_60628_12232# a_60716_10567# 0.0027f
C729 a_58052_11044# a_57692_11000# 0.08707f
C730 _330_.A1 a_37980_17272# 0.01775f
C731 a_44028_25156# VPWR 0.00979f
C732 _260_.A1 _327_.A2 0.92796f
C733 a_57044_17316# a_57132_17272# 0.28563f
C734 a_47525_29480# _393_.A1 0.07735f
C735 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I 0.00642f
C736 a_25124_28776# VPWR 0.03032f
C737 a_48060_1159# a_48508_1159# 0.0131f
C738 _301_.A1 _300_.A2 0.15634f
C739 a_36996_2824# a_36860_1592# 0.00154f
C740 a_47028_18884# VPWR 0.01378f
C741 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I 0.00482f
C742 a_65668_18884# a_66116_18884# 0.01328f
C743 a_1380_25156# VPWR 0.20348f
C744 _300_.A2 a_39236_20072# 0.0026f
C745 a_59796_29480# VPWR 0.00407f
C746 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN VPWR 0.77212f
C747 a_24564_20452# VPWR 0.20692f
C748 a_1468_27815# a_1380_27912# 0.28563f
C749 _459_.Q _334_.A1 0.07657f
C750 _375_.Z a_21287_29076# 0.00513f
C751 _451_.Q a_40692_21640# 0.02217f
C752 a_60212_25156# a_60064_25156# 0.00128f
C753 a_3172_15748# a_2812_15704# 0.08717f
C754 _355_.C _355_.ZN 0.26505f
C755 a_59036_12568# VPWR 0.31547f
C756 a_34844_15704# a_34980_15368# 0.00168f
C757 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN VPWR 0.72524f
C758 a_15580_29383# a_15492_29480# 0.28563f
C759 a_52004_15368# a_52452_15368# 0.01328f
C760 a_55004_21543# a_55364_21640# 0.08663f
C761 _437_.A1 _441_.A3 0.01574f
C762 _324_.C a_57156_27912# 0.00303f
C763 a_59732_10664# VPWR 0.20614f
C764 _340_.A2 _454_.Q 0.02608f
C765 a_3708_8999# a_4068_9096# 0.08717f
C766 a_4940_7431# a_5300_7528# 0.08674f
C767 a_54108_15271# a_54020_15368# 0.28563f
C768 a_64412_5863# a_64772_5960# 0.08717f
C769 _370_.ZN uo_out[7] 0.04986f
C770 _294_.A2 a_36948_29860# 0.0028f
C771 a_65308_4295# a_65668_4392# 0.08717f
C772 _476_.Q a_51620_19911# 0.00988f
C773 _362_.B a_35874_27937# 0.00515f
C774 _474_.Q a_49492_18840# 0.03909f
C775 a_32964_15368# VPWR 0.20348f
C776 a_55452_15271# a_55900_15271# 0.0131f
C777 a_50724_24908# VPWR 0.00571f
C778 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN 0.11044f
C779 a_51240_23340# _281_.A1 0.00747f
C780 a_18828_21976# a_19276_21976# 0.01288f
C781 a_67996_2727# a_67908_2824# 0.28563f
C782 _371_.A1 _336_.Z 0.01408f
C783 a_36412_15271# VPWR 0.32932f
C784 a_1828_14180# a_1916_14136# 0.28563f
C785 _459_.CLK _234_.ZN 0.03057f
C786 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN VPWR 0.88997f
C787 a_26220_23544# a_26132_22020# 0.0027f
C788 a_36972_16839# a_37420_16839# 0.01288f
C789 a_40916_16936# a_40804_15748# 0.02666f
C790 a_41948_17433# VPWR 0.00266f
C791 _230_.I _250_.ZN 0.30656f
C792 a_64300_23111# vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN 0.00705f
C793 _433_.ZN _304_.A1 0.03118f
C794 a_13452_30951# uio_oe[2] 0.04244f
C795 a_31732_23588# a_31820_23544# 0.28563f
C796 a_64860_7431# VPWR 0.30145f
C797 a_29828_1256# VPWR 0.20348f
C798 a_48868_1256# a_49316_1256# 0.01328f
C799 a_30476_23544# a_30924_23544# 0.01255f
C800 a_66652_4295# VPWR 0.29679f
C801 a_60964_26344# VPWR 0.20701f
C802 a_49652_13800# a_50100_13800# 0.01328f
C803 a_63404_13703# a_63764_13800# 0.08707f
C804 a_28124_2727# a_28572_2727# 0.0131f
C805 a_64324_3204# a_64188_2727# 0.00168f
C806 _346_.B a_21268_27912# 0.00183f
C807 _417_.A2 _419_.Z 0.06329f
C808 a_13004_30951# VPWR 0.31184f
C809 _334_.A1 _461_.D 0.04669f
C810 _359_.B a_31088_30301# 0.00363f
C811 a_50412_16839# a_50772_16936# 0.08717f
C812 a_21404_23111# a_21428_22020# 0.0016f
C813 a_63428_18504# VPWR 0.20348f
C814 a_53684_10664# a_53796_9476# 0.02666f
C815 _358_.A3 a_31844_26344# 0.13484f
C816 a_9532_1159# a_9444_1256# 0.28563f
C817 a_47300_1636# VPWR 0.2147f
C818 a_45172_16936# VPWR 0.20665f
C819 a_27924_23588# a_27900_23111# 0.00172f
C820 a_46984_23588# a_47172_23588# 0.00843f
C821 a_21964_25112# a_21852_24679# 0.02634f
C822 _427_.ZN a_55228_20408# 0.0032f
C823 a_5052_29816# a_5500_29816# 0.01288f
C824 a_41440_28363# a_41828_28777# 0.00393f
C825 a_35204_17316# a_35652_17316# 0.01328f
C826 a_31620_17316# a_31708_17272# 0.28563f
C827 a_47300_15368# a_47164_14136# 0.00154f
C828 a_51108_15368# a_51108_14180# 0.05841f
C829 a_9892_2824# VPWR 0.21003f
C830 a_26692_1636# a_26556_1159# 0.00168f
C831 a_50300_1592# a_50748_1592# 0.01288f
C832 a_54244_1636# a_54332_1592# 0.28563f
C833 _330_.A1 a_49764_26724# 0.03948f
C834 a_64548_11044# a_64996_11044# 0.01328f
C835 a_61412_11044# a_61052_11000# 0.08707f
C836 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I a_57940_20452# 0.00244f
C837 a_58500_21640# a_58388_20452# 0.02666f
C838 _393_.A3 a_47476_28292# 0.00228f
C839 a_15692_23111# a_16140_23111# 0.0131f
C840 a_36548_26724# VPWR 0.2056f
C841 a_10652_29816# uio_oe[4] 0.00113f
C842 a_21540_28292# a_22548_28292# 0.00196f
C843 _416_.A2 a_46848_20893# 0.00351f
C844 a_53996_18407# a_54356_18504# 0.08674f
C845 a_67124_20452# a_68020_20452# 0.0023f
C846 a_63428_15368# VPWR 0.20897f
C847 a_57044_18504# VPWR 0.20744f
C848 a_19724_25112# VPWR 0.32344f
C849 a_51457_29861# VPWR 0.98114f
C850 a_16052_27912# a_16500_27912# 0.01328f
C851 vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN VPWR 0.84115f
C852 a_54824_22045# a_54692_20452# 0.00128f
C853 a_45820_12135# VPWR 0.29679f
C854 _378_.I a_20396_27815# 0.00169f
C855 a_32964_15748# a_32604_15704# 0.08707f
C856 _359_.ZN a_34308_26344# 0.11567f
C857 a_28932_2824# a_29380_2824# 0.01328f
C858 _336_.Z a_30476_25112# 0.01569f
C859 a_36288_23208# VPWR 0.01381f
C860 _260_.A2 _325_.A1 0.02612f
C861 a_43580_15704# a_43580_15271# 0.05841f
C862 _251_.A1 a_61940_29076# 0.0012f
C863 a_60064_25156# VPWR 0.00645f
C864 _428_.Z a_52920_22760# 0.00187f
C865 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I 0.00562f
C866 a_21316_21640# a_21204_20452# 0.02666f
C867 a_19524_21640# a_19500_20408# 0.0016f
C868 _386_.A4 _393_.A3 0.12265f
C869 _362_.ZN a_32476_29167# 0.02057f
C870 a_3708_15704# VPWR 0.33374f
C871 a_55364_15368# VPWR 0.20348f
C872 _301_.A1 a_38325_22804# 0.00355f
C873 a_43824_18147# a_44459_18559# 0.02112f
C874 a_42896_18504# a_44752_18147# 0.02307f
C875 _359_.B a_34448_25597# 0.00623f
C876 a_54356_24776# clk 0.0155f
C877 a_26132_22020# a_25772_21976# 0.08707f
C878 a_4604_21976# a_4516_20452# 0.0027f
C879 a_31820_23544# a_31732_22020# 0.00151f
C880 a_46180_14180# a_46268_14136# 0.28563f
C881 a_49764_14180# a_50212_14180# 0.01328f
C882 a_37532_17272# a_37444_15748# 0.00151f
C883 a_40108_16839# VPWR 0.31253f
C884 a_47860_16936# a_47748_15748# 0.02666f
C885 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN _249_.A2 0.03625f
C886 a_27668_31048# a_26916_31048# 0.00282f
C887 a_52228_1256# VPWR 0.20348f
C888 _395_.A1 clkload0.Z 0.00559f
C889 _412_.ZN _478_.D 0.00152f
C890 a_57492_17316# VPWR 0.20944f
C891 a_64188_14136# a_64100_12612# 0.00151f
C892 _226_.ZN _302_.Z 0.03907f
C893 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN VPWR 0.88149f
C894 _402_.A1 a_41440_28363# 0.04794f
C895 a_30812_17272# VPWR 0.30073f
C896 a_61076_10664# a_60964_9476# 0.02666f
C897 a_28348_23111# a_28372_22020# 0.0016f
C898 a_53436_1592# VPWR 0.3289f
C899 a_56796_1592# a_56932_1256# 0.00168f
C900 a_20508_1159# a_20868_1256# 0.08717f
C901 a_50636_12135# a_50996_12232# 0.08707f
C902 a_13340_1592# a_13788_1592# 0.01288f
C903 a_13700_29480# a_14148_29480# 0.01328f
C904 a_23532_23544# a_23556_23208# 0.00172f
C905 a_64300_12135# a_64972_12135# 0.00544f
C906 _408_.ZN a_50704_27912# 0.00291f
C907 _229_.I _250_.A2 0.3279f
C908 _474_.CLK a_54692_18884# 0.01028f
C909 _252_.ZN a_60404_28292# 0.05367f
C910 _325_.B a_43468_16839# 0.03228f
C911 a_60276_29032# a_60852_28292# 0.00141f
C912 a_12356_29860# a_11996_29816# 0.08707f
C913 _317_.A2 a_35816_21192# 0.53413f
C914 _336_.A2 a_27028_23588# 0.00718f
C915 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_59732_14180# 0.00767f
C916 a_57604_1636# a_57244_1592# 0.08707f
C917 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN 0.03379f
C918 a_45080_29535# VPWR 0.00204f
C919 a_32292_2824# VPWR 0.20348f
C920 a_14796_23111# a_14708_23208# 0.28563f
C921 _393_.A3 _407_.A1 0.00208f
C922 a_18716_24679# a_18628_24776# 0.28563f
C923 _300_.ZN _302_.Z 0.07943f
C924 a_51332_24372# a_52852_24372# 0.01147f
C925 a_64324_9096# a_64772_9096# 0.01328f
C926 a_4068_9476# VPWR 0.2157f
C927 a_65220_7528# a_65668_7528# 0.01328f
C928 a_45372_14136# VPWR 0.30073f
C929 a_66116_5960# a_66564_5960# 0.01328f
C930 a_67012_4392# a_67460_4392# 0.01328f
C931 a_54780_26247# VPWR 0.32437f
C932 _384_.A1 _475_.Q 0.18516f
C933 a_30812_18407# a_31172_18504# 0.08717f
C934 _417_.A2 _424_.A1 0.0043f
C935 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I VPWR 0.77811f
C936 _362_.B a_33148_25641# 0.00123f
C937 a_35232_24029# a_36300_23544# 0.00506f
C938 _268_.A1 a_52764_27815# 0.00151f
C939 _373_.A2 a_26427_29977# 0.00392f
C940 _261_.ZN _304_.A1 0.0274f
C941 a_67660_12135# VPWR 0.31389f
C942 a_17060_29480# VPWR 0.20716f
C943 a_39460_15748# a_39908_15748# 0.01328f
C944 _304_.B a_39772_20408# 0.00374f
C945 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN a_62564_29032# 0.00263f
C946 _234_.ZN uo_out[7] 0.05433f
C947 a_3620_24776# VPWR 0.22347f
C948 a_20003_29611# a_20191_29611# 0.00762f
C949 a_58911_30644# _237_.A1 0.0121f
C950 a_2364_19975# a_2276_20072# 0.28563f
C951 a_42596_15748# VPWR 0.23951f
C952 _437_.A1 _330_.A1 0.7957f
C953 a_43936_27165# a_43564_27209# 0.10745f
C954 a_43008_26795# a_44864_27165# 0.02307f
C955 a_45284_9476# a_45372_9432# 0.28563f
C956 a_30476_21976# a_30924_21976# 0.01255f
C957 a_31732_22020# a_31820_21976# 0.28563f
C958 _402_.A1 a_50176_26724# 0.00468f
C959 _246_.B2 a_60793_29860# 0.00353f
C960 _327_.Z _330_.A2 0.83212f
C961 a_54804_16936# a_54692_15748# 0.02666f
C962 a_36960_27912# a_37516_27599# 0.8399f
C963 _443_.D a_37888_27555# 0.07535f
C964 _268_.A2 a_52756_29076# 0.30474f
C965 _241_.I0 a_56964_26724# 0.00671f
C966 a_50524_2727# a_50972_2727# 0.0131f
C967 a_3620_12612# a_4068_12612# 0.01328f
C968 a_7292_1592# a_7428_1256# 0.00168f
C969 a_1828_12612# a_1468_12568# 0.08717f
C970 a_25928_25273# VPWR 0.00218f
C971 a_53124_17316# a_53100_16839# 0.00172f
C972 a_29184_25597# a_28891_25273# 0.49319f
C973 a_49180_17272# a_49292_16839# 0.02634f
C974 _459_.CLK a_23084_28248# 0.00989f
C975 _251_.A1 a_63616_31128# 1.30158f
C976 a_60276_29032# _238_.I 0.43738f
C977 a_47297_25596# clkbuf_1_0__f_clk.I 0.00242f
C978 a_50436_17316# VPWR 0.24967f
C979 _419_.A4 a_47948_23111# 0.00174f
C980 a_67236_1636# VPWR 0.20952f
C981 a_31932_1159# a_31844_1256# 0.28563f
C982 a_65532_1592# a_65668_1256# 0.00168f
C983 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN a_62756_27912# 0.00369f
C984 a_61612_12135# a_61524_12232# 0.28563f
C985 a_21204_31048# uio_out[4] 0.00286f
C986 a_20644_1636# a_20284_1592# 0.08707f
C987 a_23196_21543# VPWR 0.31547f
C988 a_17148_29816# a_17596_29816# 0.01255f
C989 _421_.A1 _284_.B 0.04071f
C990 a_16052_26344# a_16052_25156# 0.05841f
C991 _324_.C vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN 0.02795f
C992 _416_.A1 _392_.A2 0.02849f
C993 a_47300_17316# a_47748_17316# 0.01328f
C994 a_65532_11000# a_65420_10567# 0.02634f
C995 a_51532_10567# a_51980_10567# 0.01288f
C996 a_54692_2824# VPWR 0.20348f
C997 a_64100_1636# a_64548_1636# 0.01328f
C998 _417_.A2 _416_.A2 0.00595f
C999 a_53124_27912# a_53572_27912# 0.01328f
C1000 a_25436_23111# a_25796_23208# 0.08663f
C1001 a_4068_23208# a_4852_23208# 0.00276f
C1002 _352_.A2 a_29575_28293# 0.10242f
C1003 a_53796_9476# VPWR 0.20692f
C1004 a_20060_21543# a_20508_21543# 0.01288f
C1005 a_60964_14180# VPWR 0.23032f
C1006 _264_.B a_41564_24679# 0.01874f
C1007 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN a_56596_18504# 0.00341f
C1008 a_21764_2824# a_21852_1159# 0.0027f
C1009 _474_.Q a_47860_23208# 0.04248f
C1010 a_35204_31048# _459_.CLK 0.00144f
C1011 a_61524_12232# VPWR 0.20622f
C1012 a_39772_20408# VPWR 0.29803f
C1013 a_51332_2824# a_51780_2824# 0.01328f
C1014 a_5276_30951# a_5412_29860# 0.00154f
C1015 _288_.ZN a_36284_29167# 0.00212f
C1016 a_32088_24831# VPWR 0.00204f
C1017 _319_.A2 a_37744_20452# 0.02791f
C1018 a_66900_20072# VPWR 0.20595f
C1019 _452_.Q _301_.A1 0.00107f
C1020 a_11772_2727# a_11684_2824# 0.28563f
C1021 _319_.A3 a_34160_20523# 0.02697f
C1022 _452_.Q a_39236_20072# 0.00438f
C1023 a_11548_30951# uio_oe[4] 0.00221f
C1024 a_48732_15704# VPWR 0.2987f
C1025 _397_.A1 clkload0.Z 0.00603f
C1026 a_45696_20072# VPWR 1.10648f
C1027 a_50524_9432# a_50972_9432# 0.0131f
C1028 a_52228_9476# a_52900_9476# 0.00347f
C1029 _288_.ZN _362_.B 0.00215f
C1030 _495_.I a_41440_28363# 0.00468f
C1031 a_28672_31048# _373_.A2 0.02497f
C1032 a_17284_31048# uio_out[7] 0.00506f
C1033 a_63428_15368# a_63404_13703# 0.00131f
C1034 a_56796_14136# a_57244_14136# 0.01222f
C1035 _325_.A2 _332_.Z 0.02808f
C1036 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN 0.00635f
C1037 a_4604_11000# a_4516_9476# 0.0027f
C1038 _373_.ZN _337_.A3 0.01442f
C1039 a_46180_12612# a_45820_12568# 0.08707f
C1040 _402_.A1 a_38816_27555# 0.01033f
C1041 a_62420_23208# vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I 0.00142f
C1042 _325_.A1 a_44276_20072# 0.10539f
C1043 _284_.A2 a_50792_26344# 0.00467f
C1044 a_20956_24679# a_20980_23588# 0.0016f
C1045 a_17596_1159# VPWR 0.29825f
C1046 a_42908_1159# a_43268_1256# 0.08717f
C1047 a_58388_12232# a_58836_12232# 0.01328f
C1048 _460_.D a_32980_25641# 0.00144f
C1049 a_4852_12232# a_4964_11044# 0.02666f
C1050 a_27140_1636# a_27588_1636# 0.01328f
C1051 a_20420_21640# VPWR 0.20641f
C1052 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I _249_.A2 0.15137f
C1053 a_62396_11000# a_62420_10664# 0.00172f
C1054 a_48508_10567# a_48420_10664# 0.28563f
C1055 a_42996_18840# a_43344_19001# 0.00277f
C1056 _452_.CLK a_39236_26344# 0.00667f
C1057 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN clk 0.02619f
C1058 _330_.A1 a_34732_19975# 0.01016f
C1059 _330_.A1 a_36076_18407# 0.0039f
C1060 a_54356_20072# a_54444_18407# 0.00151f
C1061 a_33164_24679# a_33612_24679# 0.01222f
C1062 a_64772_9476# VPWR 0.21055f
C1063 a_56348_30951# ui_in[4] 0.00362f
C1064 a_63876_20072# a_64324_20072# 0.01328f
C1065 a_67460_6340# VPWR 0.20348f
C1066 a_17844_23588# VPWR 0.20639f
C1067 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.0823f
C1068 a_18716_21543# a_19076_21640# 0.08707f
C1069 a_65308_3160# VPWR 0.33761f
C1070 a_47612_13703# VPWR 0.29679f
C1071 _455_.Q a_23627_27967# 0.00964f
C1072 _416_.A3 a_47164_18407# 0.01463f
C1073 _452_.CLK _330_.A2 0.04121f
C1074 _419_.A4 a_49448_20936# 0.00127f
C1075 _424_.A2 a_51240_20452# 0.00171f
C1076 a_54692_26344# a_54804_25156# 0.02666f
C1077 a_26160_27165# a_27140_26724# 0.00702f
C1078 _465_.D a_20672_30301# 0.00589f
C1079 _397_.A4 _282_.ZN 0.30239f
C1080 a_17732_31048# _459_.CLK 0.00656f
C1081 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN a_55140_27912# 0.01924f
C1082 a_53124_15748# a_53572_15748# 0.01328f
C1083 a_50660_11044# VPWR 0.22943f
C1084 a_49540_15748# a_49628_15704# 0.28563f
C1085 _337_.A3 a_28124_26680# 0.02721f
C1086 a_34084_28776# VPWR 0.02454f
C1087 a_33152_22091# _316_.A3 0.00528f
C1088 a_41788_2727# a_41924_1636# 0.00154f
C1089 _474_.CLK _424_.A2 0.38548f
C1090 a_56964_26724# a_57276_27208# 0.00685f
C1091 _287_.A1 _285_.Z 0.07674f
C1092 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN _250_.B 0.1232f
C1093 _451_.Q a_40580_20072# 0.03538f
C1094 a_1380_26344# VPWR 0.20348f
C1095 a_22748_2727# a_23108_2824# 0.08717f
C1096 _355_.C a_17844_27912# 0.00231f
C1097 a_39256_28292# uo_out[7] 0.0117f
C1098 _384_.A1 a_54444_23544# 0.0194f
C1099 _275_.ZN a_50996_28292# 0.00272f
C1100 _438_.A2 a_37179_24831# 0.00497f
C1101 _474_.CLK a_52228_17316# 0.00201f
C1102 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN 0.0588f
C1103 a_2724_28292# VPWR 0.20782f
C1104 a_44786_24120# a_44906_23588# 0.00165f
C1105 a_40676_25640# _264_.B 0.0091f
C1106 a_64996_14180# a_65084_14136# 0.28563f
C1107 a_16052_20452# a_15692_20408# 0.08717f
C1108 a_17396_20452# a_17844_20452# 0.01328f
C1109 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I a_65644_23544# 0.04641f
C1110 a_17372_30951# uio_out[7] 0.00619f
C1111 _327_.A2 a_44276_20072# 0.0105f
C1112 a_60285_30600# a_60909_30600# 0.10419f
C1113 a_52540_12568# a_53124_12612# 0.01675f
C1114 _260_.A1 hold2.I 0.00278f
C1115 _478_.D _427_.ZN 0.05297f
C1116 a_39996_1159# VPWR 0.32824f
C1117 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.02262f
C1118 a_54332_1159# a_54244_1256# 0.28563f
C1119 _218_.ZN a_50748_20408# 0.00156f
C1120 a_45920_20523# a_46800_20937# 0.00306f
C1121 _355_.C _351_.ZN 0.55542f
C1122 _229_.I a_59172_27912# 0.0073f
C1123 a_45284_10664# a_45732_10664# 0.01328f
C1124 a_59372_10567# a_59732_10664# 0.08707f
C1125 a_54780_1592# a_54780_1159# 0.05841f
C1126 a_14236_1159# a_14684_1159# 0.0131f
C1127 _381_.A2 _412_.B2 0.00426f
C1128 _304_.B a_42368_28733# 0.00243f
C1129 _459_.CLK a_41160_29083# 0.08209f
C1130 a_18740_22020# VPWR 0.21276f
C1131 a_38340_21327# VPWR 0.29435f
C1132 _432_.ZN VPWR 0.40459f
C1133 a_29692_21543# a_29604_21640# 0.28563f
C1134 a_16948_21640# a_17396_21640# 0.01328f
C1135 a_4964_18884# a_5052_18840# 0.28563f
C1136 a_25324_23544# VPWR 0.31486f
C1137 _424_.B1 a_50176_26724# 0.00131f
C1138 a_1828_13800# VPWR 0.20348f
C1139 a_53704_23219# VPWR 1.11195f
C1140 a_20060_2727# VPWR 0.3161f
C1141 _470_.Q a_48376_27508# 0.00647f
C1142 _230_.I a_63524_29098# 0.00271f
C1143 _285_.Z _293_.A2 1.20802f
C1144 a_4964_29860# VPWR 0.2085f
C1145 a_40244_18180# _332_.Z 0.17103f
C1146 a_56796_11000# VPWR 0.3337f
C1147 a_66116_15748# a_65980_15271# 0.00168f
C1148 _304_.ZN a_42168_22504# 0.11f
C1149 a_40220_26247# a_40132_26344# 0.28563f
C1150 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN a_58588_21543# 0.03498f
C1151 _340_.A2 uio_out[1] 0.40156f
C1152 a_17820_30951# _459_.CLK 0.00613f
C1153 _355_.C a_20672_30301# 0.00451f
C1154 _355_.C _337_.A3 0.37484f
C1155 _351_.ZN a_24636_25641# 0.00131f
C1156 _452_.Q a_42252_20936# 0.05428f
C1157 a_67908_15748# a_67548_15704# 0.08674f
C1158 a_19500_27815# VPWR 0.34697f
C1159 a_64412_15704# a_64860_15704# 0.0131f
C1160 _474_.CLK a_52764_27815# 0.00266f
C1161 a_34172_2727# a_34084_2824# 0.28563f
C1162 a_61612_23111# a_61524_23208# 0.28563f
C1163 _474_.Q a_50420_23233# 0.00461f
C1164 a_4604_7864# a_5052_7864# 0.01222f
C1165 a_61500_9432# a_61948_9432# 0.0131f
C1166 a_63652_9476# a_63292_9432# 0.08717f
C1167 _448_.Q a_37384_19624# 0.40385f
C1168 a_14708_23588# a_15156_23588# 0.01328f
C1169 a_15044_1256# a_15492_1256# 0.01328f
C1170 a_64324_6340# a_64772_6340# 0.01328f
C1171 a_65220_4772# a_65668_4772# 0.01328f
C1172 _330_.A1 a_39264_18147# 0.01316f
C1173 a_64324_3204# a_64412_3160# 0.28563f
C1174 a_66116_3204# a_66564_3204# 0.01328f
C1175 a_4940_13703# a_5388_13703# 0.01222f
C1176 a_60276_29032# VPWR 0.5896f
C1177 a_5724_29383# a_6172_29383# 0.0131f
C1178 a_6723_30644# a_7092_31048# 0.02397f
C1179 _416_.A1 a_46389_21236# 0.00141f
C1180 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I a_67772_24679# 0.01418f
C1181 a_13252_1636# VPWR 0.20348f
C1182 _304_.B _260_.A1 0.50752f
C1183 a_59844_12612# a_59484_12568# 0.08707f
C1184 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN 0.00718f
C1185 a_62420_13800# a_62508_12135# 0.00151f
C1186 _459_.CLK a_23084_25112# 0.01491f
C1187 a_20379_29977# uio_out[5] 0.05496f
C1188 _325_.A2 a_43452_18191# 0.01962f
C1189 a_66787_30600# vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.00587f
C1190 a_65084_1159# a_65668_1256# 0.01675f
C1191 _395_.A1 a_49764_23588# 0.00346f
C1192 _304_.B _428_.Z 0.20885f
C1193 a_62396_1159# VPWR 0.3289f
C1194 a_1916_19975# VPWR 0.297f
C1195 a_47524_11044# a_47972_11044# 0.01328f
C1196 _416_.ZN a_46576_19759# 0.00123f
C1197 a_3260_18407# VPWR 0.30487f
C1198 a_5412_1636# a_5276_1159# 0.00168f
C1199 a_1468_1592# a_1468_1159# 0.05841f
C1200 a_33276_1592# a_33724_1592# 0.01288f
C1201 a_37220_1636# a_37308_1592# 0.28563f
C1202 a_30724_16936# a_31172_16936# 0.01328f
C1203 input9.Z _267_.A2 0.00333f
C1204 _311_.Z a_36148_21976# 0.05872f
C1205 _305_.A2 a_44028_22020# 0.01071f
C1206 a_36016_20893# _325_.A2 0.00829f
C1207 a_43492_27912# _330_.A1 0.0035f
C1208 a_43940_27912# a_44388_27912# 0.01328f
C1209 _255_.I _243_.B2 0.00245f
C1210 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN 0.00199f
C1211 _437_.A1 a_38616_24328# 0.52361f
C1212 a_42368_28733# VPWR 0.21531f
C1213 a_22660_2824# a_22524_1592# 0.00154f
C1214 _467_.D _378_.I 0.00289f
C1215 _350_.A2 a_29804_30951# 0.01252f
C1216 a_24876_21976# VPWR 0.31436f
C1217 a_54432_31128# vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN 0.02048f
C1218 _452_.CLK a_31932_23111# 0.0048f
C1219 _279_.Z _473_.Q 0.04508f
C1220 a_42236_2727# VPWR 0.34979f
C1221 a_63316_13800# VPWR 0.20622f
C1222 a_31080_29977# VPWR 0.00204f
C1223 a_44948_22020# VPWR 0.0086f
C1224 a_17484_26247# a_17932_26247# 0.0131f
C1225 a_3260_26247# a_3620_26344# 0.08717f
C1226 _474_.CLK a_55228_20408# 0.05312f
C1227 a_11100_29816# VPWR 0.33743f
C1228 a_63092_16936# a_63068_15704# 0.0016f
C1229 a_3708_10567# VPWR 0.33374f
C1230 a_31260_15271# a_31620_15368# 0.08717f
C1231 a_29692_23111# VPWR 0.31431f
C1232 _452_.CLK a_43400_18909# 0.01963f
C1233 a_36960_27912# a_37840_27599# 0.00306f
C1234 _284_.ZN uo_out[3] 0.04003f
C1235 _424_.A2 _398_.C 0.42886f
C1236 _260_.A1 a_41880_24072# 0.00383f
C1237 a_45148_2727# a_45508_2824# 0.08717f
C1238 a_53908_24776# _384_.A1 0.03719f
C1239 _452_.CLK _304_.A1 0.00924f
C1240 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN a_56596_29861# 0.00198f
C1241 _452_.Q a_39268_18840# 0.03812f
C1242 _441_.A2 _438_.ZN 0.00874f
C1243 _399_.ZN _417_.A2 0.21113f
C1244 a_67436_16839# a_67348_16936# 0.28563f
C1245 a_65308_18407# a_66092_18407# 0.00443f
C1246 _459_.CLK a_29232_29931# 0.00773f
C1247 a_61052_26247# VPWR 0.3289f
C1248 a_64860_9432# a_64860_8999# 0.05841f
C1249 _355_.C a_21044_27508# 0.00689f
C1250 a_21876_23588# a_21516_23544# 0.08663f
C1251 _403_.ZN a_44571_26841# 0.00582f
C1252 a_4156_25112# a_4604_25112# 0.01222f
C1253 a_1916_13703# a_1828_13800# 0.28563f
C1254 a_27028_20452# a_26668_20408# 0.08717f
C1255 a_28372_20452# a_28820_20452# 0.01328f
C1256 _287_.A1 _371_.A1 0.07167f
C1257 _363_.Z _223_.ZN 0.03543f
C1258 a_62980_18504# a_62980_17316# 0.05841f
C1259 _330_.ZN a_38564_15748# 0.0011f
C1260 a_37108_23588# VPWR 0.20368f
C1261 a_3260_16839# a_3172_16936# 0.28563f
C1262 a_23196_29816# a_23644_29816# 0.01222f
C1263 _260_.A1 VPWR 1.81001f
C1264 a_19388_1592# VPWR 0.34002f
C1265 _419_.Z a_45920_20523# 0.00407f
C1266 a_35516_1592# a_35652_1256# 0.00168f
C1267 a_66340_12612# a_66788_12612# 0.01328f
C1268 a_63204_12612# a_62844_12568# 0.08707f
C1269 _459_.CLK _335_.ZN 0.00382f
C1270 _371_.A2 _352_.A2 0.89007f
C1271 a_47047_21640# VPWR 0.0065f
C1272 _428_.Z VPWR 0.55493f
C1273 a_63316_12232# a_63292_11000# 0.0016f
C1274 a_49652_12232# a_49740_10567# 0.00151f
C1275 a_65980_15271# a_66340_15368# 0.0869f
C1276 _474_.CLK a_56572_23111# 0.01139f
C1277 a_40580_1636# a_40220_1592# 0.08707f
C1278 a_4068_26724# a_4156_26680# 0.28563f
C1279 _395_.A2 a_50420_23233# 0.01931f
C1280 a_67124_10664# a_67572_10664# 0.01328f
C1281 a_36636_1159# a_37084_1159# 0.0131f
C1282 _452_.CLK _448_.D 0.07981f
C1283 hold2.I _260_.A2 0.85194f
C1284 a_58063_30644# _246_.B2 0.00241f
C1285 a_28124_26680# a_27328_25227# 0.00104f
C1286 _304_.B _470_.Q 0.30575f
C1287 a_4964_20452# VPWR 0.21167f
C1288 _397_.A1 a_50120_26476# 0.41478f
C1289 _388_.B a_44612_31048# 0.04305f
C1290 a_66564_2824# a_66652_1159# 0.0027f
C1291 _397_.Z a_48321_23208# 0.00267f
C1292 a_61300_16936# a_61748_16936# 0.01328f
C1293 _452_.Q a_42154_21236# 0.59984f
C1294 a_52452_12612# VPWR 0.21241f
C1295 a_64636_2727# VPWR 0.33348f
C1296 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN VPWR 0.79103f
C1297 a_4156_29383# a_4068_29480# 0.28563f
C1298 _416_.A3 _475_.Q 0.03057f
C1299 a_40580_15368# a_41028_15368# 0.01328f
C1300 a_33412_20072# VPWR 0.20644f
C1301 _355_.C _342_.ZN 0.53765f
C1302 _416_.A1 a_43936_27165# 0.00235f
C1303 a_4156_15704# a_4156_15271# 0.05841f
C1304 a_26556_27815# a_26468_27912# 0.28563f
C1305 a_65420_10567# VPWR 0.32173f
C1306 a_42684_15271# a_42596_15368# 0.28563f
C1307 a_27364_23208# VPWR 0.22345f
C1308 a_37084_21543# a_37444_21640# 0.08663f
C1309 a_64860_17272# a_64884_16936# 0.00172f
C1310 a_41572_18504# _452_.D 0.0018f
C1311 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I a_60852_15748# 0.01054f
C1312 _274_.A3 _274_.A2 0.17636f
C1313 a_44028_15271# a_44476_15271# 0.0131f
C1314 _336_.A1 VPWR 1.34865f
C1315 _249_.A2 VPWR 1.20474f
C1316 _448_.Q a_38676_20452# 0.00532f
C1317 a_15604_22020# a_16052_22020# 0.01328f
C1318 a_62980_15748# VPWR 0.20595f
C1319 _327_.Z a_39684_20072# 0.0113f
C1320 a_40220_19975# a_40580_20072# 0.08663f
C1321 a_56572_2727# a_56484_2824# 0.28563f
C1322 a_54444_23544# clk 0.00613f
C1323 a_60516_26344# a_60212_25156# 0.00283f
C1324 _311_.Z a_36288_23208# 0.01235f
C1325 _421_.A1 a_46984_23588# 0.06096f
C1326 _395_.A1 _404_.A1 0.29083f
C1327 a_38971_18559# a_39324_17272# 0.00158f
C1328 a_37444_1256# a_37892_1256# 0.01328f
C1329 a_22212_23208# a_22300_21543# 0.0027f
C1330 a_25684_23588# a_25324_23544# 0.08717f
C1331 a_6980_1256# VPWR 0.20348f
C1332 a_3172_4772# VPWR 0.20993f
C1333 a_20532_25156# a_20172_25112# 0.08707f
C1334 a_8996_31048# VPWR 0.23348f
C1335 a_1380_7908# VPWR 0.20348f
C1336 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN a_58476_17272# 0.00143f
C1337 a_16700_2727# a_17148_2727# 0.0131f
C1338 _251_.A1 a_61748_26724# 0.00116f
C1339 a_52428_13703# a_52788_13800# 0.08707f
C1340 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I a_58612_16936# 0.00323f
C1341 a_58700_16839# vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I 0.02518f
C1342 a_34960_22505# VPWR 0.00124f
C1343 a_66316_13703# a_66764_13703# 0.0131f
C1344 _324_.C a_65072_29860# 1.20192f
C1345 a_37444_26344# _444_.D 0.00481f
C1346 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN a_63092_26724# 0.00289f
C1347 a_39212_16839# a_39572_16936# 0.08707f
C1348 a_46180_10664# a_46180_9476# 0.05841f
C1349 a_64972_16839# VPWR 0.32113f
C1350 a_33188_1636# VPWR 0.2051f
C1351 a_64996_31048# a_65072_29860# 0.00135f
C1352 _327_.A2 a_41600_19376# 0.00102f
C1353 a_3620_1636# a_3260_1592# 0.08707f
C1354 a_43132_27815# VPWR 0.32469f
C1355 _261_.ZN a_40004_22020# 0.01325f
C1356 a_1828_29860# a_2276_29860# 0.01328f
C1357 a_62308_27912# a_62396_26247# 0.00151f
C1358 _330_.A1 a_35088_20893# 0.04415f
C1359 a_3620_17316# a_4068_17316# 0.01328f
C1360 a_1828_17316# a_1468_17272# 0.08717f
C1361 a_58500_21640# VPWR 0.16149f
C1362 _237_.A1 _243_.A1 0.00744f
C1363 a_57604_11044# a_57692_11000# 0.28563f
C1364 a_56148_23588# clk 0.00645f
C1365 a_53660_11000# a_54108_11000# 0.01288f
C1366 a_52564_16936# a_53012_16936# 0.01328f
C1367 a_46940_1592# a_47388_1592# 0.012f
C1368 a_31484_30951# _334_.A1 0.00108f
C1369 a_932_20072# a_932_18884# 0.05841f
C1370 a_57044_17316# a_56684_17272# 0.0869f
C1371 _384_.ZN _384_.A1 0.6288f
C1372 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_57044_23588# 0.00504f
C1373 _304_.B _260_.A2 0.67216f
C1374 a_65668_26344# vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I 0.00473f
C1375 _381_.Z _279_.Z 0.00123f
C1376 _300_.A2 a_38788_20072# 0.00187f
C1377 a_932_25156# VPWR 0.22176f
C1378 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I 0.022f
C1379 a_62564_29032# VPWR 0.48565f
C1380 vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I 0.00534f
C1381 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN _274_.A1 0.0336f
C1382 _336_.A1 a_28903_24776# 0.02535f
C1383 a_24116_20452# VPWR 0.20692f
C1384 a_15244_27815# a_15692_27815# 0.0131f
C1385 a_1020_27815# a_1380_27912# 0.08717f
C1386 _470_.Q VPWR 1.40608f
C1387 _375_.Z a_21103_29076# 0.00578f
C1388 _451_.Q a_40244_21640# 0.03187f
C1389 a_2724_15748# a_2812_15704# 0.28563f
C1390 a_58588_12568# VPWR 0.32371f
C1391 _355_.C a_27328_25227# 0.02611f
C1392 _474_.CLK _258_.I 0.00454f
C1393 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN 0.0033f
C1394 a_17508_2824# a_17956_2824# 0.01328f
C1395 a_15132_29383# a_15492_29480# 0.08717f
C1396 a_26556_30951# a_26720_30301# 0.00105f
C1397 a_55004_21543# a_54916_21640# 0.28563f
C1398 a_3708_8999# a_3620_9096# 0.28563f
C1399 a_59284_10664# VPWR 0.20614f
C1400 a_4940_7431# a_4852_7528# 0.28563f
C1401 a_53660_15271# a_54020_15368# 0.08717f
C1402 a_64412_5863# a_64324_5960# 0.28563f
C1403 a_44162_24120# a_44786_24120# 0.10711f
C1404 _294_.A2 a_36500_29860# 0.00351f
C1405 a_65308_4295# a_65220_4392# 0.28563f
C1406 a_29232_29931# uo_out[7] 0.01797f
C1407 _362_.B a_34586_27912# 0.00847f
C1408 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN 0.00669f
C1409 a_50464_24908# VPWR 0.0161f
C1410 _474_.Q a_48172_18840# 0.02634f
C1411 a_32516_15368# VPWR 0.20348f
C1412 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I a_58836_18884# 0.0056f
C1413 a_67548_2727# a_67908_2824# 0.08674f
C1414 a_35964_15271# VPWR 0.32932f
C1415 _416_.A1 _431_.A3 0.19886f
C1416 a_1828_14180# a_1468_14136# 0.08717f
C1417 _438_.A2 _448_.Q 0.18738f
C1418 _459_.CLK a_40038_28720# 0.0435f
C1419 a_3620_14180# a_4068_14180# 0.01328f
C1420 a_63092_26724# VPWR 0.20934f
C1421 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN ui_in[7] 0.00202f
C1422 a_40992_17433# VPWR 0.00205f
C1423 a_33776_29123# VPWR 0.69845f
C1424 a_31732_23588# a_31372_23544# 0.0869f
C1425 a_13004_30951# uio_oe[2] 0.00531f
C1426 _335_.ZN uo_out[7] 0.04668f
C1427 a_64412_7431# VPWR 0.3038f
C1428 a_25643_25273# a_25888_25641# 0.00232f
C1429 a_29380_1256# VPWR 0.20348f
C1430 a_66204_4295# VPWR 0.31657f
C1431 a_60516_26344# VPWR 0.16298f
C1432 a_63404_13703# a_63316_13800# 0.28563f
C1433 a_36100_17316# a_36076_16839# 0.00172f
C1434 a_32156_17272# a_32156_16839# 0.05841f
C1435 a_12548_31048# VPWR 0.3785f
C1436 a_50412_16839# a_50324_16936# 0.28563f
C1437 a_2276_23208# a_2276_22020# 0.05841f
C1438 _359_.B a_29788_30345# 0.01037f
C1439 a_62980_18504# VPWR 0.20348f
C1440 a_44724_16936# VPWR 0.20665f
C1441 a_46852_1636# VPWR 0.2085f
C1442 a_9084_1159# a_9444_1256# 0.08717f
C1443 a_53324_12135# a_53772_12135# 0.01288f
C1444 a_67324_12568# a_67212_12135# 0.02634f
C1445 a_2276_29480# a_2724_29480# 0.01328f
C1446 a_10116_1636# a_10564_1636# 0.01328f
C1447 _294_.A2 _462_.D 0.03155f
C1448 a_24428_23544# a_24540_23111# 0.02634f
C1449 _427_.ZN a_54780_20408# 0.00393f
C1450 a_26720_30301# a_28054_30196# 0.00639f
C1451 a_31620_17316# a_31260_17272# 0.08707f
C1452 _258_.I _247_.ZN 0.38813f
C1453 a_54244_1636# a_53884_1592# 0.08707f
C1454 a_60964_11044# a_61052_11000# 0.28563f
C1455 a_51196_11000# a_51084_10567# 0.02634f
C1456 a_9444_2824# VPWR 0.20815f
C1457 _393_.A3 a_46804_28292# 0.02035f
C1458 _274_.A2 _324_.C 0.00215f
C1459 a_36100_26724# VPWR 0.12999f
C1460 a_17472_28363# a_18352_28777# 0.00306f
C1461 a_21540_28292# a_21628_28248# 0.28563f
C1462 a_15692_24679# a_16140_24679# 0.0131f
C1463 a_57580_17272# vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I 0.00151f
C1464 _434_.ZN a_38529_22804# 0.00631f
C1465 _416_.A2 a_45920_20523# 0.01573f
C1466 a_53996_18407# a_53908_18504# 0.28563f
C1467 _260_.A2 VPWR 1.14741f
C1468 a_59036_1159# a_59484_1159# 0.0131f
C1469 a_66316_20408# a_66764_20408# 0.01222f
C1470 a_67124_20452# a_67212_20408# 0.28563f
C1471 a_62980_15368# VPWR 0.20897f
C1472 _303_.ZN _324_.B 0.05651f
C1473 a_50468_29977# VPWR 0.00127f
C1474 a_67548_18840# a_67996_18840# 0.01222f
C1475 a_56596_18504# VPWR 0.14909f
C1476 _304_.B a_52744_26031# 0.05911f
C1477 a_19276_25112# VPWR 0.35601f
C1478 vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN 0.0048f
C1479 a_45372_12135# VPWR 0.30073f
C1480 _378_.I a_19948_27815# 0.00344f
C1481 a_32516_15748# a_32604_15704# 0.28563f
C1482 a_36100_15748# a_36548_15748# 0.01328f
C1483 _336_.Z a_30388_25156# 0.03245f
C1484 a_20508_2727# a_20644_1636# 0.00154f
C1485 a_36084_23208# VPWR 0.00666f
C1486 a_59226_25156# VPWR 0.01435f
C1487 _459_.CLK _343_.A2 0.68137f
C1488 _251_.A1 a_59572_29076# 0.00753f
C1489 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN a_64188_27815# 0.01307f
C1490 _428_.Z a_51240_23340# 0.23097f
C1491 _427_.B1 _395_.A3 0.06709f
C1492 _397_.A1 _404_.A1 0.07135f
C1493 _383_.ZN _470_.Q 0.00112f
C1494 _452_.CLK a_41900_16839# 0.00239f
C1495 a_3260_15704# VPWR 0.30487f
C1496 _362_.ZN a_32848_29123# 0.01668f
C1497 a_54916_15368# VPWR 0.20348f
C1498 _301_.A1 a_38131_22804# 0.00101f
C1499 a_42896_18504# a_44459_18559# 0.41635f
C1500 a_43824_18147# a_43452_18191# 0.10745f
C1501 a_29268_22020# a_29716_22020# 0.01328f
C1502 a_53908_24776# clk 0.0155f
C1503 a_25684_22020# a_25772_21976# 0.28563f
C1504 a_46180_14180# a_45820_14136# 0.08707f
C1505 a_47500_16839# a_47948_16839# 0.01288f
C1506 _248_.B1 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I 0.00587f
C1507 a_39660_16839# VPWR 0.3281f
C1508 a_59844_1256# a_60292_1256# 0.01328f
C1509 _395_.A1 a_48384_26724# 0.01592f
C1510 a_36748_23544# a_37196_23544# 0.01255f
C1511 a_51780_1256# VPWR 0.20348f
C1512 a_27004_30951# a_26916_31048# 0.28563f
C1513 _412_.ZN a_51988_24776# 0.01557f
C1514 a_39100_2727# a_39548_2727# 0.0131f
C1515 a_60180_13800# a_60628_13800# 0.01328f
C1516 a_57044_17316# VPWR 0.20744f
C1517 _359_.ZN a_34155_25273# 0.0029f
C1518 _459_.CLK a_29716_23588# 0.00808f
C1519 a_37892_17316# VPWR 0.21341f
C1520 a_35088_20893# a_35723_20569# 0.02112f
C1521 a_19972_23208# a_20084_22020# 0.02666f
C1522 a_52988_1592# VPWR 0.3289f
C1523 a_64188_12568# a_64212_12232# 0.00172f
C1524 a_20508_1159# a_20420_1256# 0.28563f
C1525 _243_.A1 _242_.Z 0.26788f
C1526 a_50636_12135# a_50548_12232# 0.28563f
C1527 _229_.I a_60940_28248# 0.02131f
C1528 _474_.CLK a_54244_18884# 0.01949f
C1529 a_15492_29860# a_15940_29860# 0.01328f
C1530 a_11908_29860# a_11996_29816# 0.28563f
C1531 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I 0.09666f
C1532 _325_.B a_43020_16839# 0.0022f
C1533 _358_.A3 a_34396_24679# 0.00285f
C1534 _336_.A2 a_26580_23588# 0.00484f
C1535 a_54780_26247# a_54804_25156# 0.0016f
C1536 a_36148_21976# a_35816_21192# 0.00136f
C1537 _317_.A2 a_35268_21640# 0.00443f
C1538 a_4852_15368# a_4940_13703# 0.00151f
C1539 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_59284_14180# 0.01133f
C1540 _268_.A2 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I 0.03409f
C1541 a_58140_11000# a_58028_10567# 0.02634f
C1542 a_31844_2824# VPWR 0.20839f
C1543 a_60740_1636# a_61188_1636# 0.01328f
C1544 a_57156_1636# a_57244_1592# 0.28563f
C1545 a_44132_29535# VPWR 0.00246f
C1546 _300_.ZN a_39172_22504# 0.00111f
C1547 _247_.B a_60276_26724# 0.01172f
C1548 a_17932_24679# a_18628_24776# 0.01227f
C1549 a_26556_23111# a_27004_23111# 0.01288f
C1550 a_3620_9476# VPWR 0.22347f
C1551 _251_.A1 _257_.B 0.00693f
C1552 a_54692_2824# a_54692_1636# 0.05841f
C1553 a_50884_2824# a_50748_1592# 0.00154f
C1554 a_10340_2824# a_10428_1159# 0.0027f
C1555 a_52452_14180# VPWR 0.20968f
C1556 a_52744_26031# VPWR 0.18592f
C1557 a_30812_18407# a_30724_18504# 0.28563f
C1558 a_64188_27815# VPWR 0.32292f
C1559 _474_.CLK _478_.D 0.01103f
C1560 a_3172_31048# a_3172_29860# 0.05841f
C1561 _373_.A2 a_26720_30301# 0.00234f
C1562 _250_.B VPWR 0.41198f
C1563 a_67212_12135# VPWR 0.31389f
C1564 a_16612_29480# VPWR 0.20703f
C1565 a_39908_2824# a_40356_2824# 0.01328f
C1566 a_43750_23544# a_44302_23588# 0.00212f
C1567 _419_.A4 _281_.ZN 0.06099f
C1568 a_3172_24776# VPWR 0.20993f
C1569 a_40038_28720# uo_out[7] 0.8159f
C1570 a_932_6340# VPWR 0.22176f
C1571 _452_.CLK _424_.A2 0.53547f
C1572 _223_.I _459_.CLK 0.185f
C1573 a_28260_21640# a_28372_20452# 0.02666f
C1574 a_58687_31220# _237_.A1 0.00223f
C1575 a_42148_15748# VPWR 0.21644f
C1576 a_1916_19975# a_2276_20072# 0.08717f
C1577 a_57132_23544# a_57020_23111# 0.02634f
C1578 a_43008_26795# a_43564_27209# 0.8399f
C1579 a_46628_9476# a_47076_9476# 0.01328f
C1580 a_31732_22020# a_31372_21976# 0.0869f
C1581 _402_.A1 a_49952_26724# 0.00177f
C1582 a_52540_14136# a_53124_14180# 0.01675f
C1583 _327_.Z a_38644_19368# 0.02593f
C1584 a_36960_27912# a_37888_27555# 1.16391f
C1585 a_24980_25273# VPWR 0.00246f
C1586 vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I 0.63458f
C1587 a_1380_12612# a_1468_12568# 0.28563f
C1588 a_51308_18407# a_51332_17316# 0.0016f
C1589 _459_.CLK a_22636_28248# 0.00575f
C1590 a_40468_25157# _435_.ZN 0.00246f
C1591 _251_.A1 a_62532_30736# 0.00121f
C1592 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN a_61076_20452# 0.00102f
C1593 a_23108_23208# a_23084_21976# 0.0016f
C1594 a_26916_23208# a_27028_22020# 0.02666f
C1595 a_49988_17316# VPWR 0.21666f
C1596 a_31484_1159# a_31844_1256# 0.08717f
C1597 a_58588_12568# a_58500_11044# 0.00151f
C1598 a_61164_12135# a_61524_12232# 0.08707f
C1599 a_47076_12232# a_47524_12232# 0.01328f
C1600 a_66788_1636# VPWR 0.20952f
C1601 a_20196_1636# a_20284_1592# 0.28563f
C1602 _359_.B _288_.ZN 0.13803f
C1603 a_17956_29860# a_18044_29816# 0.28563f
C1604 a_22748_21543# VPWR 0.31547f
C1605 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN a_53212_27815# 0.0058f
C1606 a_45128_26031# _284_.B 0.00697f
C1607 a_55004_11000# a_55028_10664# 0.00172f
C1608 a_40580_1636# a_40444_1159# 0.00168f
C1609 a_54244_2824# VPWR 0.22423f
C1610 a_1380_2824# a_1380_1636# 0.05841f
C1611 a_20420_24776# a_20868_24776# 0.01328f
C1612 a_25436_23111# a_25348_23208# 0.28563f
C1613 _384_.ZN clk 0.10592f
C1614 a_53348_9476# VPWR 0.20692f
C1615 a_60268_14136# VPWR 0.31817f
C1616 _260_.A1 _260_.ZN 0.41941f
C1617 _229_.I _246_.B2 0.10684f
C1618 a_35988_18504# a_36436_18504# 0.01328f
C1619 _452_.CLK a_33524_24776# 0.00648f
C1620 _424_.B1 a_50300_20408# 0.00108f
C1621 _324_.C _279_.Z 0.00157f
C1622 a_11460_31048# a_11460_29860# 0.05841f
C1623 a_42236_15704# a_42684_15704# 0.01288f
C1624 a_61076_12232# VPWR 0.20622f
C1625 _474_.D a_51620_19911# 0.00489f
C1626 a_31140_24831# VPWR 0.00246f
C1627 a_56516_26344# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.03312f
C1628 a_66452_20072# VPWR 0.21172f
C1629 a_11324_2727# a_11684_2824# 0.08717f
C1630 a_11091_30644# uio_oe[4] 0.04236f
C1631 _395_.A3 _422_.ZN 0.00868f
C1632 _397_.A1 a_48384_26724# 0.02636f
C1633 a_48284_15704# VPWR 0.29679f
C1634 _452_.Q a_38788_20072# 0.00217f
C1635 a_63516_19975# a_63964_19975# 0.0131f
C1636 a_44276_20072# VPWR 0.64143f
C1637 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I a_64100_27912# 0.00285f
C1638 _355_.C a_20496_26344# 0.00261f
C1639 a_52228_9476# a_52316_9432# 0.28563f
C1640 _442_.ZN _435_.A3 0.00949f
C1641 _252_.ZN a_60740_26724# 0.01976f
C1642 a_1828_20452# a_2276_20452# 0.01328f
C1643 a_46492_17272# a_46404_15748# 0.00151f
C1644 _447_.Q a_42982_21730# 0.00289f
C1645 _412_.A1 _412_.ZN 1.08416f
C1646 _223_.I _371_.A3 0.41162f
C1647 _459_.CLK a_24952_29032# 0.02894f
C1648 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN VPWR 0.94344f
C1649 a_61276_2727# a_61948_2727# 0.00544f
C1650 a_49316_12612# a_49764_12612# 0.01328f
C1651 a_45732_12612# a_45820_12568# 0.28563f
C1652 a_66652_18840# a_66564_17316# 0.00151f
C1653 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.00345f
C1654 a_17148_1159# VPWR 0.29679f
C1655 a_42908_1159# a_42820_1256# 0.28563f
C1656 a_932_7908# a_1020_7864# 0.28563f
C1657 a_65668_5960# a_65668_4772# 0.05841f
C1658 a_61948_12568# a_61860_11044# 0.00151f
C1659 a_64772_7528# a_64772_6340# 0.05841f
C1660 a_22996_29480# _345_.A2 0.00125f
C1661 a_66564_4392# a_66564_3204# 0.05841f
C1662 a_35292_26247# a_35740_26247# 0.01255f
C1663 a_19972_21640# VPWR 0.20677f
C1664 a_50076_17272# a_50524_17272# 0.01288f
C1665 a_62060_10567# a_62508_10567# 0.01288f
C1666 a_48060_10567# a_48420_10664# 0.08717f
C1667 _454_.Q a_26556_27815# 0.02988f
C1668 a_2812_1159# a_3260_1159# 0.0131f
C1669 _330_.A1 a_35628_18407# 0.00188f
C1670 a_24004_23208# a_24452_23208# 0.01328f
C1671 a_56932_23208# VPWR 0.21824f
C1672 _251_.A1 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I 0.12987f
C1673 _395_.A1 _399_.A2 0.00773f
C1674 a_64324_9476# VPWR 0.22973f
C1675 a_17396_23588# VPWR 0.20348f
C1676 a_67012_6340# VPWR 0.20348f
C1677 a_66564_2824# a_66428_1592# 0.00154f
C1678 a_47164_13703# VPWR 0.29679f
C1679 a_18716_21543# a_18628_21640# 0.28563f
C1680 a_64860_3160# VPWR 0.33437f
C1681 a_30588_21543# a_31036_21543# 0.01288f
C1682 _238_.I _252_.B 0.02916f
C1683 _455_.Q a_22620_27599# 0.00753f
C1684 ui_in[2] ui_in[1] 0.2231f
C1685 a_26160_27165# a_25867_26841# 0.49319f
C1686 _465_.D a_20379_29977# 0.02945f
C1687 _424_.A2 a_50748_20408# 0.00145f
C1688 _223_.I uo_out[7] 0.02702f
C1689 a_17284_31048# _459_.CLK 0.0062f
C1690 _398_.C _478_.D 0.73268f
C1691 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN a_53572_27912# 0.00308f
C1692 a_49540_15748# a_49180_15704# 0.08707f
C1693 _311_.A2 VPWR 2.38091f
C1694 a_50212_11044# VPWR 0.22223f
C1695 a_12444_29816# a_12444_29383# 0.05841f
C1696 a_62308_2824# a_62756_2824# 0.01328f
C1697 _324_.C _304_.ZN 0.00325f
C1698 _443_.D uo_out[7] 0.00149f
C1699 _337_.A3 a_27676_26680# 0.0199f
C1700 _459_.Q a_29232_29931# 0.05686f
C1701 a_56964_26724# a_56836_27208# 0.00284f
C1702 a_61860_27912# a_61836_26680# 0.0016f
C1703 _474_.CLK a_46198_27060# 0.01911f
C1704 _441_.ZN a_40468_25157# 0.00176f
C1705 a_37067_19001# VPWR 0.3704f
C1706 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN a_63952_29480# 0.00316f
C1707 a_932_26344# VPWR 0.22176f
C1708 _451_.Q a_40132_20072# 0.00989f
C1709 a_22748_2727# a_22660_2824# 0.28563f
C1710 a_38772_28292# uo_out[7] 0.00102f
C1711 _267_.A2 a_52964_29480# 0.00167f
C1712 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN a_55228_20408# 0.03478f
C1713 a_2276_28292# VPWR 0.20634f
C1714 a_57604_9476# a_58052_9476# 0.01328f
C1715 _474_.CLK a_51780_17316# 0.00198f
C1716 a_3620_1256# a_4068_1256# 0.01328f
C1717 _474_.CLK clkbuf_1_0__f_clk.I 0.00384f
C1718 _459_.Q _335_.ZN 0.1807f
C1719 a_38523_27967# a_38808_27967# 0.00277f
C1720 a_4068_31048# a_4740_31048# 0.00347f
C1721 a_64996_14180# a_64636_14136# 0.08707f
C1722 a_15604_20452# a_15692_20408# 0.28563f
C1723 a_61052_14136# a_61500_14136# 0.01288f
C1724 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I a_65196_23544# 0.00218f
C1725 _284_.A2 a_46156_25112# 0.00353f
C1726 a_16916_31048# uio_out[7] 0.00401f
C1727 a_21180_1592# a_21316_1256# 0.00168f
C1728 _397_.Z _399_.A1 0.01489f
C1729 a_51444_13800# a_51532_12135# 0.00151f
C1730 _416_.A1 a_44688_26399# 0.00126f
C1731 _352_.A2 a_25524_26344# 0.01909f
C1732 _261_.ZN _301_.A1 0.54211f
C1733 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN 0.93238f
C1734 a_53660_1159# a_54244_1256# 0.01675f
C1735 a_39548_1159# VPWR 0.29679f
C1736 _218_.ZN a_50300_20408# 0.03805f
C1737 a_1380_11044# a_1828_11044# 0.01328f
C1738 a_61836_16839# a_62284_16839# 0.0131f
C1739 a_29916_1592# a_30364_1592# 0.01288f
C1740 a_48868_31048# a_48104_30219# 0.01115f
C1741 _454_.Q a_23834_28292# 0.00253f
C1742 a_46848_20893# a_47483_20569# 0.02112f
C1743 a_45920_20523# a_46308_20937# 0.00393f
C1744 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.01046f
C1745 _355_.C a_24304_26795# 0.02179f
C1746 a_59372_10567# a_59284_10664# 0.28563f
C1747 a_1828_18504# a_1828_17316# 0.05841f
C1748 _304_.B _476_.Q 0.14441f
C1749 _459_.CLK a_37584_29123# 0.0325f
C1750 _381_.A2 a_50792_26344# 0.00242f
C1751 a_18292_22020# VPWR 0.21304f
C1752 _389_.ZN _404_.A1 0.03476f
C1753 a_37444_21640# VPWR 0.20784f
C1754 a_24876_23544# VPWR 0.31389f
C1755 a_4964_18884# a_4604_18840# 0.08674f
C1756 a_19388_2727# VPWR 0.38777f
C1757 _461_.D _335_.ZN 0.01166f
C1758 a_2364_18840# a_2812_18840# 0.0131f
C1759 a_29244_21543# a_29604_21640# 0.08707f
C1760 _294_.ZN _223_.ZN 0.22507f
C1761 a_1380_13800# VPWR 0.20348f
C1762 a_40692_21640# a_40580_20452# 0.02666f
C1763 _447_.Q _304_.A1 0.48684f
C1764 _285_.Z a_37968_31048# 0.00898f
C1765 a_4516_29860# VPWR 0.20847f
C1766 _393_.ZN VPWR 0.59026f
C1767 a_37408_18504# a_37796_18191# 0.00393f
C1768 a_39772_26247# a_40132_26344# 0.0869f
C1769 a_33396_26344# a_33188_25940# 0.01342f
C1770 a_56348_11000# VPWR 0.31471f
C1771 a_62620_15704# a_62620_15271# 0.05841f
C1772 _245_.Z a_60212_25156# 0.00564f
C1773 _355_.C a_20379_29977# 0.04479f
C1774 _424_.B1 _384_.A3 0.45875f
C1775 a_17372_30951# _459_.CLK 0.00613f
C1776 _474_.Q a_51620_19911# 0.00109f
C1777 _351_.ZN a_25008_25597# 0.00349f
C1778 a_67460_15748# a_67548_15704# 0.28563f
C1779 _400_.ZN _470_.D 0.18404f
C1780 a_17932_27815# VPWR 0.3491f
C1781 _403_.ZN _397_.A4 0.05216f
C1782 a_22620_27599# a_22964_27967# 0.00275f
C1783 a_60604_26247# a_60212_25156# 0.0016f
C1784 _260_.A2 _260_.ZN 0.18524f
C1785 a_49600_30180# a_50012_29977# 0.00275f
C1786 a_33724_2727# a_34084_2824# 0.08717f
C1787 a_61164_23111# a_61524_23208# 0.08717f
C1788 _474_.Q a_48321_23208# 0.04642f
C1789 a_64212_23588# a_64660_23588# 0.01328f
C1790 _435_.A3 _435_.ZN 0.12393f
C1791 _330_.A1 _312_.ZN 0.00129f
C1792 _251_.A1 a_56964_26724# 0.29761f
C1793 a_49492_18840# a_50280_19369# 0.02112f
C1794 a_63204_9476# a_63292_9432# 0.28563f
C1795 uio_in[6] uio_in[5] 0.01021f
C1796 _330_.A1 a_38971_18559# 0.01046f
C1797 a_1020_3160# a_1020_2727# 0.05841f
C1798 a_20844_20408# a_21292_20408# 0.0131f
C1799 a_6172_30951# a_7092_31048# 0.00794f
C1800 a_6723_30644# a_6084_31048# 0.00397f
C1801 _351_.A2 a_25867_26841# 0.00486f
C1802 a_55452_12568# a_55900_12568# 0.01288f
C1803 a_59396_12612# a_59484_12568# 0.28563f
C1804 a_54804_26724# a_54780_26247# 0.00172f
C1805 a_12804_1636# VPWR 0.20348f
C1806 _447_.Q _448_.D 0.00273f
C1807 _459_.CLK a_22636_25112# 0.00116f
C1808 _325_.A2 a_43824_18147# 0.02204f
C1809 a_10652_29816# a_10788_29480# 0.00168f
C1810 a_61948_1159# VPWR 0.33352f
C1811 a_36436_18504# a_36524_16839# 0.00151f
C1812 a_45696_20072# a_46576_19759# 0.00306f
C1813 a_1468_19975# VPWR 0.29679f
C1814 a_65084_1159# a_64996_1256# 0.28563f
C1815 a_2812_18407# VPWR 0.30213f
C1816 a_37220_1636# a_36860_1592# 0.08707f
C1817 _474_.CLK vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I 0.00501f
C1818 a_59732_12232# a_59844_11044# 0.02666f
C1819 a_37444_25156# a_37532_25112# 0.28563f
C1820 a_55924_12232# a_55900_11000# 0.0016f
C1821 _381_.A2 _281_.ZN 0.29273f
C1822 _416_.A3 a_49068_20408# 0.00244f
C1823 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN a_61836_23544# 0.00637f
C1824 a_43044_27912# _330_.A1 0.00848f
C1825 _476_.Q VPWR 1.41019f
C1826 a_55924_10664# a_56372_10664# 0.01328f
C1827 a_27676_26247# VPWR 0.31075f
C1828 a_25212_1159# a_25660_1159# 0.0131f
C1829 a_35540_18504# a_35652_17316# 0.02666f
C1830 a_932_1636# a_1380_1636# 0.01328f
C1831 a_24428_21976# VPWR 0.31436f
C1832 _337_.A3 a_26916_27912# 0.05508f
C1833 _324_.C a_44340_26183# 0.03391f
C1834 a_52024_20083# a_52944_19759# 0.00306f
C1835 _452_.CLK a_31484_23111# 0.00241f
C1836 a_27812_21640# a_28260_21640# 0.01328f
C1837 a_62868_13800# VPWR 0.20622f
C1838 input9.Z _276_.A2 0.12281f
C1839 a_30132_29977# VPWR 0.00246f
C1840 a_41788_2727# VPWR 0.31731f
C1841 a_44500_22020# VPWR 0.00866f
C1842 a_3260_26247# a_3172_26344# 0.28563f
C1843 _474_.CLK a_54780_20408# 0.02021f
C1844 a_4068_15368# a_4852_15368# 0.00276f
C1845 a_10652_29816# VPWR 0.33458f
C1846 a_3260_10567# VPWR 0.30487f
C1847 a_66004_16936# a_66116_15748# 0.02666f
C1848 a_31260_15271# a_31172_15368# 0.28563f
C1849 a_55676_2727# a_55812_1636# 0.00154f
C1850 _452_.Q a_42168_22504# 0.02296f
C1851 a_29244_23111# VPWR 0.31916f
C1852 a_32604_15271# a_33052_15271# 0.0131f
C1853 _441_.B _434_.ZN 0.18566f
C1854 _245_.Z VPWR 0.58573f
C1855 a_45148_2727# a_45060_2824# 0.28563f
C1856 _294_.A2 a_31964_28292# 0.00349f
C1857 _346_.A2 a_21876_25156# 0.00192f
C1858 a_65220_17316# a_65668_17316# 0.01328f
C1859 a_51620_19911# a_51968_20127# 0.00277f
C1860 a_60604_26247# VPWR 0.32908f
C1861 a_66988_16839# a_67348_16936# 0.0869f
C1862 a_1468_8999# a_1916_8999# 0.0131f
C1863 a_53996_24679# _478_.D 0.00116f
C1864 a_26020_1256# a_26468_1256# 0.01328f
C1865 a_17484_23544# a_17932_23544# 0.01288f
C1866 a_65756_7864# a_65756_7431# 0.05841f
C1867 _398_.C clkbuf_1_0__f_clk.I 0.27276f
C1868 a_2364_7431# a_2812_7431# 0.0131f
C1869 a_21428_23588# a_21516_23544# 0.28563f
C1870 a_3260_5863# a_3708_5863# 0.0131f
C1871 a_4156_4295# a_4940_4295# 0.00443f
C1872 a_67548_4728# a_67548_4295# 0.05841f
C1873 a_66652_6296# a_66652_5863# 0.05841f
C1874 _403_.ZN a_44864_27165# 0.00484f
C1875 a_5276_2727# a_5724_2727# 0.0131f
C1876 a_55116_13703# a_55564_13703# 0.01288f
C1877 a_1468_13703# a_1828_13800# 0.08717f
C1878 a_37332_16936# a_37308_15271# 0.00134f
C1879 a_26580_20452# a_26668_20408# 0.28563f
C1880 a_16700_29383# a_17148_29383# 0.012f
C1881 a_36660_23588# VPWR 0.20417f
C1882 a_64860_26247# a_65756_26247# 0.00373f
C1883 _287_.A1 a_30388_28776# 0.024f
C1884 _459_.Q a_30596_28292# 0.00689f
C1885 a_2812_16839# a_3172_16936# 0.08717f
C1886 a_18940_1592# VPWR 0.30582f
C1887 a_62756_12612# a_62844_12568# 0.28563f
C1888 a_8627_30644# a_9084_30951# 0.00916f
C1889 _325_.B a_43888_19204# 0.00177f
C1890 _325_.A1 a_42392_19243# 0.32337f
C1891 _371_.A2 a_28364_28776# 0.00374f
C1892 a_37584_29123# uo_out[7] 0.01411f
C1893 a_50084_24328# VPWR 0.60884f
C1894 a_65980_15271# a_65892_15368# 0.28563f
C1895 _249_.A2 _248_.B1 0.77561f
C1896 _304_.A1 a_40004_23233# 0.00496f
C1897 a_50300_11000# a_50748_11000# 0.01288f
C1898 a_66676_12232# a_66788_11044# 0.02666f
C1899 a_41364_16936# a_41812_16936# 0.01328f
C1900 a_43716_1636# a_44164_1636# 0.01328f
C1901 a_40132_1636# a_40220_1592# 0.28563f
C1902 _474_.CLK a_56124_23111# 0.02157f
C1903 _340_.A2 _343_.A2 0.02362f
C1904 a_67548_15704# a_67684_15368# 0.00168f
C1905 a_1468_26680# a_1916_26680# 0.0131f
C1906 a_4068_26724# a_3708_26680# 0.08717f
C1907 _384_.A3 _218_.ZN 0.17872f
C1908 _268_.A2 _416_.A1 0.32747f
C1909 _252_.B VPWR 1.1402f
C1910 _334_.A1 uo_out[4] 0.0242f
C1911 a_4516_20452# VPWR 0.20862f
C1912 _435_.A3 _441_.ZN 0.05536f
C1913 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I 0.01521f
C1914 _388_.B a_44164_31048# 0.02836f
C1915 _397_.A2 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.00432f
C1916 _452_.Q a_40780_21543# 0.00915f
C1917 a_64188_2727# VPWR 0.32977f
C1918 a_52004_12612# VPWR 0.20622f
C1919 a_17844_26344# a_18628_26344# 0.00276f
C1920 a_6172_2727# a_6308_1636# 0.00154f
C1921 a_6084_2824# a_6532_2824# 0.01328f
C1922 a_32964_20072# VPWR 0.20348f
C1923 a_58924_17272# vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I 0.00138f
C1924 a_3708_29383# a_4068_29480# 0.08717f
C1925 _355_.C a_24864_29931# 0.00133f
C1926 _416_.A1 a_43008_26795# 0.03627f
C1927 _427_.B1 _422_.ZN 0.16957f
C1928 a_64972_10567# VPWR 0.32368f
C1929 a_42236_15271# a_42596_15368# 0.08717f
C1930 a_23627_27967# a_23872_27599# 0.00232f
C1931 a_30476_21976# a_30588_21543# 0.02634f
C1932 a_25884_27815# a_26468_27912# 0.01675f
C1933 a_37084_21543# a_36996_21640# 0.28563f
C1934 _436_.B a_41384_26841# 0.00103f
C1935 a_26916_23208# VPWR 0.22387f
C1936 a_54804_16936# a_54780_15704# 0.0016f
C1937 _452_.CLK hold1.Z 0.07091f
C1938 a_14708_28292# a_15156_28292# 0.01328f
C1939 a_35156_29860# uo_out[4] 0.01597f
C1940 _451_.Q _330_.A2 0.05576f
C1941 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I VPWR 0.88122f
C1942 _448_.Q a_38228_20452# 0.02583f
C1943 a_56124_2727# a_56484_2824# 0.08717f
C1944 a_62532_15748# VPWR 0.20595f
C1945 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I _241_.Z 0.00491f
C1946 _416_.A1 a_46852_17316# 0.0016f
C1947 _327_.Z a_39236_20072# 0.00153f
C1948 a_40220_19975# a_40132_20072# 0.28563f
C1949 a_21964_23544# a_21876_22020# 0.00151f
C1950 a_33412_16936# a_33412_15748# 0.05841f
C1951 _311_.Z a_36084_23208# 0.00396f
C1952 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN a_64772_20072# 0.00173f
C1953 a_39264_18147# a_39236_17316# 0.00687f
C1954 a_52116_18504# a_52564_18504# 0.01328f
C1955 a_6532_1256# VPWR 0.20348f
C1956 a_7540_31048# VPWR 0.21155f
C1957 a_25236_23588# a_25324_23544# 0.28563f
C1958 a_20084_25156# a_20172_25112# 0.28563f
C1959 a_2724_4772# VPWR 0.20782f
C1960 a_16140_25112# a_16588_25112# 0.01288f
C1961 a_52428_13703# a_52340_13800# 0.28563f
C1962 a_58700_16839# a_58612_16936# 0.28563f
C1963 _476_.Q _424_.B2 0.06761f
C1964 _268_.A1 _267_.A1 0.06979f
C1965 a_52920_22760# a_53300_23047# 0.49319f
C1966 a_31820_20408# a_32268_20408# 0.0131f
C1967 a_25652_31048# a_26108_30951# 0.0065f
C1968 a_36996_26344# _444_.D 0.00481f
C1969 _359_.B a_34586_27912# 0.00173f
C1970 a_39212_16839# a_39124_16936# 0.28563f
C1971 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN a_62644_26724# 0.00142f
C1972 _327_.A2 a_42392_19243# 0.00674f
C1973 a_32740_1636# VPWR 0.20348f
C1974 a_64524_16839# VPWR 0.31934f
C1975 a_42684_27815# VPWR 0.34216f
C1976 a_20532_23588# a_20508_23111# 0.00172f
C1977 a_59932_12568# a_59820_12135# 0.02634f
C1978 a_3172_1636# a_3260_1592# 0.28563f
C1979 a_6756_1636# a_7204_1636# 0.01328f
C1980 a_16588_23544# a_16588_23111# 0.05841f
C1981 a_2364_12135# a_2812_12135# 0.0131f
C1982 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_62564_29032# 0.04353f
C1983 a_1380_17316# a_1468_17272# 0.28563f
C1984 _447_.Q a_39684_20072# 0.00131f
C1985 a_55364_21640# VPWR 0.21043f
C1986 a_57604_11044# a_57244_11000# 0.08707f
C1987 a_4156_11000# a_4156_10567# 0.05841f
C1988 a_55700_23588# clk 0.00532f
C1989 a_60180_12232# a_60268_10567# 0.00151f
C1990 _274_.A1 _267_.A2 1.20293f
C1991 a_67772_24679# vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I 0.00285f
C1992 a_56596_17316# a_56684_17272# 0.28563f
C1993 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_56596_23588# 0.02731f
C1994 a_47612_1159# a_48060_1159# 0.0131f
C1995 a_17484_27815# a_16240_26795# 0.00102f
C1996 a_36548_2824# a_36412_1592# 0.00154f
C1997 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN 0.66087f
C1998 a_65220_18884# a_65668_18884# 0.01328f
C1999 a_1020_27815# a_932_27912# 0.28563f
C2000 a_53212_29816# _274_.A1 0.37347f
C2001 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I 0.00575f
C2002 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I 0.65153f
C2003 a_23668_20452# VPWR 0.20692f
C2004 _336_.A1 a_28679_24776# 0.00213f
C2005 _459_.Q _223_.I 0.20549f
C2006 a_58140_12568# VPWR 0.35527f
C2007 a_2724_15748# a_2364_15704# 0.08717f
C2008 a_4516_15748# a_4964_15748# 0.01328f
C2009 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_63092_26724# 0.00452f
C2010 a_34396_15704# a_34532_15368# 0.00168f
C2011 a_15132_29383# a_15044_29480# 0.28563f
C2012 _390_.ZN _395_.A2 0.38239f
C2013 a_51556_15368# a_52004_15368# 0.01328f
C2014 a_54556_21543# a_54916_21640# 0.0869f
C2015 a_58836_10664# VPWR 0.20677f
C2016 a_53660_15271# a_53572_15368# 0.28563f
C2017 a_3260_8999# a_3620_9096# 0.08717f
C2018 a_43750_23544# a_44786_24120# 0.00135f
C2019 a_4156_7431# a_4852_7528# 0.01227f
C2020 a_932_5960# a_1380_5960# 0.01328f
C2021 a_64860_4295# a_65220_4392# 0.08717f
C2022 a_4852_21640# a_4964_20452# 0.02666f
C2023 a_62560_25112# vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I 0.15173f
C2024 _294_.A2 a_35818_29860# 0.01186f
C2025 _474_.Q a_47724_18840# 0.00163f
C2026 _402_.A1 _402_.B 1.32102f
C2027 _251_.A1 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN 0.01982f
C2028 a_55004_15271# a_55452_15271# 0.0131f
C2029 a_32068_15368# VPWR 0.20348f
C2030 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN a_65556_23588# 0.00359f
C2031 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I a_58388_18884# 0.00143f
C2032 _475_.D a_46352_20569# 0.00165f
C2033 a_67548_2727# a_67460_2824# 0.28563f
C2034 a_51240_23340# _476_.Q 0.00183f
C2035 _416_.A1 a_38752_26344# 0.00114f
C2036 a_18380_21976# a_18828_21976# 0.01288f
C2037 _459_.CLK a_38584_28292# 0.00139f
C2038 a_35516_15271# VPWR 0.32974f
C2039 a_62644_26724# VPWR 0.20657f
C2040 a_36524_16839# a_36972_16839# 0.01288f
C2041 a_1380_14180# a_1468_14136# 0.28563f
C2042 a_40468_16936# a_40356_15748# 0.02666f
C2043 a_25772_23544# a_25684_22020# 0.00151f
C2044 a_43814_21236# a_44038_21236# 0.75472f
C2045 a_67908_17316# VPWR 0.21197f
C2046 a_33483_29535# VPWR 0.3773f
C2047 a_32740_23208# a_32828_21543# 0.00108f
C2048 a_48420_1256# a_48868_1256# 0.01328f
C2049 a_28932_1256# VPWR 0.20348f
C2050 a_5388_7431# VPWR 0.35526f
C2051 a_31284_23588# a_31372_23544# 0.28563f
C2052 a_12548_31048# uio_oe[2] 0.00261f
C2053 a_65756_4295# VPWR 0.31505f
C2054 a_27676_2727# a_28124_2727# 0.0131f
C2055 a_62956_13703# a_63316_13800# 0.08707f
C2056 a_60013_26344# VPWR 0.00671f
C2057 a_49204_13800# a_49652_13800# 0.01328f
C2058 a_11548_30951# VPWR 0.37844f
C2059 a_49740_16839# a_50324_16936# 0.01675f
C2060 _223_.I _461_.D 0.00844f
C2061 _337_.ZN _371_.A1 1.8464f
C2062 _359_.B a_30160_30301# 0.00614f
C2063 a_20956_23111# a_20980_22020# 0.0016f
C2064 a_62532_18504# VPWR 0.20348f
C2065 a_44276_16936# VPWR 0.20665f
C2066 a_46404_1636# VPWR 0.20847f
C2067 _442_.ZN a_40084_25156# 0.0018f
C2068 a_9084_1159# a_8996_1256# 0.28563f
C2069 _395_.A1 _411_.A2 0.59231f
C2070 a_22059_26399# a_22304_26031# 0.00232f
C2071 a_53236_10664# a_53348_9476# 0.02666f
C2072 a_27476_23588# a_27452_23111# 0.00172f
C2073 a_21516_25112# a_21404_24679# 0.02634f
C2074 _427_.ZN a_54332_20408# 0.00393f
C2075 a_4604_29816# a_5052_29816# 0.01288f
C2076 a_26720_30301# a_26427_29977# 0.49319f
C2077 _265_.ZN a_43003_28409# 0.00347f
C2078 _407_.A1 _384_.A3 0.00776f
C2079 a_31172_17316# a_31260_17272# 0.28563f
C2080 a_34756_17316# a_35204_17316# 0.01328f
C2081 a_60380_11000# a_61052_11000# 0.00544f
C2082 a_64100_11044# a_64548_11044# 0.01328f
C2083 a_46852_15368# a_46716_14136# 0.00154f
C2084 a_52267_30644# uio_in[0] 0.00145f
C2085 a_50660_15368# a_50660_14180# 0.05841f
C2086 a_64412_15271# a_64548_14180# 0.00154f
C2087 a_8996_2824# VPWR 0.20815f
C2088 a_26244_1636# a_26108_1159# 0.00168f
C2089 a_49852_1592# a_50300_1592# 0.01288f
C2090 a_53796_1636# a_53884_1592# 0.28563f
C2091 _393_.A3 a_46580_28292# 0.00175f
C2092 a_48104_30219# _390_.ZN 0.00562f
C2093 _434_.ZN a_38325_22804# 0.00263f
C2094 a_35140_26680# VPWR 0.77503f
C2095 a_15244_23111# a_15692_23111# 0.0131f
C2096 a_17472_28363# a_17860_28777# 0.00393f
C2097 _378_.ZN a_18028_28777# 0.22974f
C2098 a_53548_18407# a_53908_18504# 0.08674f
C2099 _325_.A1 a_43828_16936# 0.00172f
C2100 a_67124_20452# a_66764_20408# 0.08663f
C2101 a_62532_15368# VPWR 0.20897f
C2102 _304_.B a_52848_25987# 0.0187f
C2103 a_54804_18504# VPWR 0.20457f
C2104 a_50012_29977# VPWR 0.00268f
C2105 a_15604_27912# a_16052_27912# 0.01328f
C2106 a_18828_25112# VPWR 0.32368f
C2107 _319_.ZN VPWR 0.83715f
C2108 _371_.ZN VPWR 0.7646f
C2109 a_32516_15748# a_32156_15704# 0.08707f
C2110 a_5388_12135# VPWR 0.35526f
C2111 _378_.I a_19500_27815# 0.01862f
C2112 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN 0.6322f
C2113 a_41340_15704# a_41476_15368# 0.00168f
C2114 _340_.A2 a_24952_29032# 0.47652f
C2115 a_28484_2824# a_28932_2824# 0.01328f
C2116 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN 0.00117f
C2117 _397_.A1 a_49212_26369# 0.00448f
C2118 a_36860_23111# VPWR 0.31803f
C2119 _474_.CLK a_56236_22505# 0.00103f
C2120 a_43132_15704# a_43132_15271# 0.05841f
C2121 _459_.CLK a_23084_29383# 0.00898f
C2122 a_19076_21640# a_19052_20408# 0.0016f
C2123 a_20868_21640# a_20756_20452# 0.02666f
C2124 _324_.C _328_.A2 0.46889f
C2125 _452_.CLK a_41452_16839# 0.00239f
C2126 a_2812_15704# VPWR 0.30213f
C2127 _362_.ZN a_31920_29480# 0.01818f
C2128 a_54468_15368# VPWR 0.20348f
C2129 a_42896_18504# a_43452_18191# 0.8399f
C2130 a_54088_22895# _427_.ZN 0.00303f
C2131 a_25684_22020# a_25324_21976# 0.08707f
C2132 _432_.ZN a_41476_24776# 0.02645f
C2133 _419_.A4 a_47636_25940# 0.02313f
C2134 a_53460_24776# clk 0.0155f
C2135 a_37084_17272# a_36996_15748# 0.00151f
C2136 a_49316_14180# a_49764_14180# 0.01328f
C2137 a_45732_14180# a_45820_14136# 0.28563f
C2138 a_47412_16936# a_47300_15748# 0.02666f
C2139 a_31372_23544# a_31284_22020# 0.00151f
C2140 a_39212_16839# VPWR 0.31397f
C2141 _248_.B1 a_64188_27815# 0.00335f
C2142 a_26556_30951# a_26916_31048# 0.08663f
C2143 a_51332_1256# VPWR 0.20348f
C2144 a_56596_17316# VPWR 0.14909f
C2145 a_63740_14136# a_63652_12612# 0.00151f
C2146 _359_.ZN a_34448_25597# 0.00391f
C2147 a_27900_23111# a_27924_22020# 0.0016f
C2148 a_20664_29977# VPWR 0.0018f
C2149 _451_.Q _304_.A1 0.06779f
C2150 a_37444_17316# VPWR 0.20348f
C2151 a_20060_1159# a_20420_1256# 0.08717f
C2152 a_56348_1592# a_56484_1256# 0.00168f
C2153 a_60628_10664# a_60516_9476# 0.02666f
C2154 a_52540_1592# VPWR 0.3289f
C2155 _229_.I a_60492_28248# 0.0156f
C2156 a_63852_12135# a_64300_12135# 0.012f
C2157 a_13252_29480# a_13700_29480# 0.01328f
C2158 a_50188_12135# a_50548_12232# 0.08707f
C2159 _395_.A1 _399_.ZN 0.10122f
C2160 a_12892_1592# a_13340_1592# 0.01288f
C2161 a_23084_23544# a_23108_23208# 0.00172f
C2162 _313_.ZN a_33724_23111# 0.02323f
C2163 _474_.CLK a_53436_18840# 0.02611f
C2164 a_11908_29860# a_11548_29816# 0.08707f
C2165 _355_.C a_18264_29480# 0.00245f
C2166 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_64188_27815# 0.01356f
C2167 vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I a_62620_19975# 0.00156f
C2168 a_37179_24831# a_37424_24463# 0.00232f
C2169 _358_.A3 a_33612_24679# 0.00283f
C2170 _317_.A2 a_35044_21640# 0.01232f
C2171 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_58836_14180# 0.04881f
C2172 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN _250_.B 0.03219f
C2173 _393_.A1 a_47733_29098# 0.00641f
C2174 a_31396_2824# VPWR 0.22891f
C2175 a_57156_1636# a_56796_1592# 0.08707f
C2176 a_5388_23111# a_5300_23208# 0.28563f
C2177 a_17932_24679# a_17844_24776# 0.28563f
C2178 a_27172_24328# a_28012_24679# 0.00611f
C2179 a_3172_9476# VPWR 0.20993f
C2180 a_64772_7528# a_65220_7528# 0.01328f
C2181 a_65668_5960# a_66116_5960# 0.01328f
C2182 a_66564_4392# a_67012_4392# 0.01328f
C2183 a_52004_14180# VPWR 0.20348f
C2184 a_67996_6296# a_67908_4772# 0.0027f
C2185 a_36076_18407# a_36524_18407# 0.012f
C2186 a_52848_25987# VPWR 0.39596f
C2187 _363_.Z _459_.CLK 0.02605f
C2188 a_39012_15748# a_39460_15748# 0.01328f
C2189 a_16164_29480# VPWR 0.22779f
C2190 a_66764_12135# VPWR 0.31389f
C2191 _460_.D VPWR 0.34605f
C2192 a_63952_29480# VPWR 0.59428f
C2193 a_38584_28292# uo_out[7] 0.03261f
C2194 a_2724_24776# VPWR 0.20782f
C2195 a_67460_7528# VPWR 0.20924f
C2196 a_31396_31048# _459_.CLK 0.00107f
C2197 a_41700_15748# VPWR 0.21074f
C2198 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN 0.9161f
C2199 a_1916_19975# a_1828_20072# 0.28563f
C2200 _255_.I a_59572_29076# 0.11039f
C2201 a_20396_27815# uio_out[6] 0.00381f
C2202 a_43008_26795# a_43936_27165# 1.16391f
C2203 a_40092_27209# a_40436_26841# 0.00275f
C2204 a_54892_18407# vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN 0.09198f
C2205 _311_.A2 _311_.Z 0.05683f
C2206 a_31284_22020# a_31372_21976# 0.28563f
C2207 _327_.Z a_39268_18840# 0.49075f
C2208 a_54356_16936# a_54244_15748# 0.02666f
C2209 _452_.CLK clkbuf_1_0__f_clk.I 0.00198f
C2210 _397_.A1 _411_.A2 1.05553f
C2211 a_49852_2727# a_50524_2727# 0.00544f
C2212 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN VPWR 0.99986f
C2213 a_6844_1592# a_6980_1256# 0.00168f
C2214 a_1380_12612# a_1020_12568# 0.08717f
C2215 a_3172_12612# a_3620_12612# 0.01328f
C2216 a_48732_17272# a_48844_16839# 0.02634f
C2217 a_52676_17316# a_52652_16839# 0.00172f
C2218 _459_.CLK a_22996_28292# 0.00585f
C2219 a_28256_25597# a_28891_25273# 0.02112f
C2220 a_49540_17316# VPWR 0.21427f
C2221 a_33724_23111# _316_.ZN 0.00246f
C2222 a_66340_1636# VPWR 0.2187f
C2223 a_5052_26680# a_4964_25156# 0.00151f
C2224 a_31484_1159# a_31396_1256# 0.28563f
C2225 a_61164_12135# a_61076_12232# 0.28563f
C2226 a_30795_29977# _371_.A1 0.00184f
C2227 a_20196_1636# a_19836_1592# 0.08707f
C2228 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN a_56036_28292# 0.00138f
C2229 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN 0.08594f
C2230 _287_.A1 a_38472_30169# 1.18488f
C2231 _474_.CLK _267_.A1 0.04326f
C2232 a_16700_29816# a_17148_29816# 0.01255f
C2233 a_17956_29860# a_17596_29816# 0.0869f
C2234 _324_.C a_61297_30300# 0.00401f
C2235 a_22300_21543# VPWR 0.33016f
C2236 a_45232_25987# _284_.B 0.00505f
C2237 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN a_52764_27815# 0.00163f
C2238 _452_.Q _434_.ZN 0.00511f
C2239 a_15604_26344# a_15604_25156# 0.05841f
C2240 a_46852_17316# a_47300_17316# 0.01328f
C2241 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN 0.00129f
C2242 a_63652_1636# a_64100_1636# 0.01328f
C2243 a_53572_2824# VPWR 0.21435f
C2244 a_51084_10567# a_51532_10567# 0.01288f
C2245 a_65084_11000# a_64972_10567# 0.02634f
C2246 a_52676_27912# a_53124_27912# 0.01328f
C2247 _474_.Q _399_.A1 0.49435f
C2248 a_3620_23208# a_4068_23208# 0.01328f
C2249 a_24988_23111# a_25348_23208# 0.08707f
C2250 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I a_63316_20452# 0.05647f
C2251 _281_.A1 a_52036_22504# 0.00112f
C2252 a_52900_9476# VPWR 0.22767f
C2253 a_21316_2824# a_21404_1159# 0.0027f
C2254 a_59820_14136# VPWR 0.29679f
C2255 a_19612_21543# a_20060_21543# 0.01288f
C2256 _260_.A1 a_41476_24776# 0.03308f
C2257 _452_.CLK a_33076_24776# 0.00825f
C2258 _255_.I _257_.B 0.05397f
C2259 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN 0.72747f
C2260 a_60628_12232# VPWR 0.20862f
C2261 a_45732_15748# a_46404_15748# 0.00347f
C2262 a_60404_28292# _252_.B 0.00974f
C2263 a_38764_20408# VPWR 0.31725f
C2264 a_50884_2824# a_51332_2824# 0.01328f
C2265 a_4828_30951# a_4964_29860# 0.00154f
C2266 _288_.ZN a_35728_29480# 0.00163f
C2267 a_66004_20072# VPWR 0.27016f
C2268 a_11324_2727# a_11236_2824# 0.28563f
C2269 a_47836_15704# VPWR 0.29679f
C2270 a_10540_30951# uio_oe[4] 0.00469f
C2271 a_64188_27815# a_64100_27912# 0.28563f
C2272 a_39536_26795# _435_.A3 0.0016f
C2273 a_52228_9476# a_51868_9432# 0.08717f
C2274 a_50076_9432# a_50524_9432# 0.0131f
C2275 a_26916_31048# _373_.A2 0.00119f
C2276 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN a_57156_14180# 0.00162f
C2277 a_62980_15368# a_62956_13703# 0.00131f
C2278 _272_.B1 ui_in[4] 0.02967f
C2279 _274_.A1 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.00243f
C2280 a_56348_14136# a_56796_14136# 0.01222f
C2281 _447_.Q a_42778_21812# 0.00155f
C2282 _473_.Q a_48084_18884# 0.00484f
C2283 _459_.CLK a_24304_29480# 0.00452f
C2284 _397_.A1 _399_.ZN 0.02574f
C2285 _373_.ZN _455_.Q 0.01603f
C2286 a_65084_30951# VPWR 0.347f
C2287 _452_.Q a_40556_16839# 0.00421f
C2288 _293_.A2 a_38472_30169# 0.1106f
C2289 a_45732_12612# a_45372_12568# 0.08707f
C2290 a_58588_21543# vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.00203f
C2291 a_20508_24679# a_20532_23588# 0.0016f
C2292 a_42236_1159# a_42820_1256# 0.01675f
C2293 a_16700_1159# VPWR 0.29679f
C2294 _330_.A1 _323_.A3 0.00948f
C2295 a_57940_12232# a_58388_12232# 0.01328f
C2296 a_26692_1636# a_27140_1636# 0.01328f
C2297 _427_.A2 a_54040_22366# 0.00655f
C2298 a_19524_21640# VPWR 0.23495f
C2299 a_53572_17316# vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN 0.00199f
C2300 a_43400_18909# a_44812_19369# 0.00393f
C2301 a_61948_11000# a_61972_10664# 0.00172f
C2302 a_48060_10567# a_47972_10664# 0.28563f
C2303 _454_.Q a_25884_27815# 0.03331f
C2304 _363_.Z uo_out[7] 0.09635f
C2305 _402_.A1 a_46352_22021# 0.10959f
C2306 a_56484_23208# VPWR 0.20488f
C2307 _330_.A1 a_35180_18407# 0.00112f
C2308 _251_.A1 a_64324_29860# 0.00853f
C2309 _438_.A2 a_39760_23588# 0.0144f
C2310 _437_.A1 a_38628_25156# 0.00375f
C2311 a_32096_24419# a_33164_24679# 0.00506f
C2312 a_52924_20127# VPWR 0.00246f
C2313 a_63740_9432# VPWR 0.33981f
C2314 a_16948_23588# VPWR 0.20348f
C2315 a_66564_6340# VPWR 0.20631f
C2316 a_46716_13703# VPWR 0.29679f
C2317 a_17932_21543# a_18628_21640# 0.01227f
C2318 _459_.CLK uo_out[3] 0.26814f
C2319 _474_.CLK _412_.A1 0.19734f
C2320 a_64412_3160# VPWR 0.33858f
C2321 a_63428_20072# a_63876_20072# 0.01328f
C2322 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I 0.00437f
C2323 _455_.Q a_22992_27555# 0.01479f
C2324 _398_.C a_51988_24776# 0.00122f
C2325 _397_.A4 _421_.A1 0.51551f
C2326 a_49092_15748# a_49180_15704# 0.28563f
C2327 a_52676_15748# a_53124_15748# 0.01328f
C2328 a_37532_25112# VPWR 0.34746f
C2329 a_49764_11044# VPWR 0.2124f
C2330 a_41340_2727# a_41476_1636# 0.00154f
C2331 _337_.A3 a_27228_26680# 0.02423f
C2332 a_36960_27912# uo_out[7] 0.00402f
C2333 a_12548_31048# a_12356_29860# 0.00285f
C2334 a_29804_30951# a_29232_29931# 0.00105f
C2335 a_50996_28292# _407_.A1 0.1068f
C2336 a_37360_19325# VPWR 0.524f
C2337 _441_.ZN a_40084_25156# 0.02168f
C2338 a_22300_2727# a_22660_2824# 0.08717f
C2339 _324_.C _412_.ZN 0.00579f
C2340 _267_.A2 a_52292_29480# 0.00109f
C2341 _395_.A2 _399_.A1 0.1873f
C2342 a_1828_28292# VPWR 0.20348f
C2343 a_4156_9432# a_4156_8999# 0.05841f
C2344 _371_.ZN _370_.B 0.00543f
C2345 a_64548_14180# a_64636_14136# 0.28563f
C2346 a_15604_20452# a_15244_20408# 0.08717f
C2347 a_16948_20452# a_17396_20452# 0.01328f
C2348 _284_.A2 a_46068_25156# 0.00634f
C2349 _397_.Z VPWR 0.5223f
C2350 _459_.CLK _371_.A2 0.14777f
C2351 a_40580_20072# _331_.ZN 0.00235f
C2352 _397_.A2 _395_.A1 0.59176f
C2353 _430_.ZN _435_.ZN 0.0044f
C2354 _460_.Q _358_.A3 1.29895f
C2355 a_52092_12568# a_52540_12568# 0.012f
C2356 _252_.ZN a_61948_27815# 0.00223f
C2357 _256_.A2 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I 0.00519f
C2358 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I 0.00286f
C2359 a_39100_1159# VPWR 0.30141f
C2360 a_53660_1159# a_53572_1256# 0.28563f
C2361 a_48420_31048# a_48104_30219# 0.00246f
C2362 a_38752_26344# _431_.A3 0.02375f
C2363 a_45920_20523# a_47483_20569# 0.41635f
C2364 _355_.C a_21600_26725# 0.00114f
C2365 a_13788_1159# a_14236_1159# 0.0131f
C2366 a_54332_1592# a_54332_1159# 0.05841f
C2367 a_58924_10567# a_59284_10664# 0.08707f
C2368 _459_.CLK a_37291_29535# 0.02583f
C2369 _381_.A2 a_47636_25940# 0.03881f
C2370 VPWR ui_in[4] 0.56355f
C2371 a_17844_22020# VPWR 0.20639f
C2372 a_45484_28248# _404_.A1 0.03319f
C2373 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I 0.25638f
C2374 a_36996_21640# VPWR 0.20921f
C2375 _294_.A2 uo_out[0] 0.00144f
C2376 a_24428_23544# VPWR 0.31389f
C2377 a_18940_2727# VPWR 0.32049f
C2378 a_53300_23047# VPWR 0.37452f
C2379 a_29244_21543# a_29156_21640# 0.28563f
C2380 a_932_13800# VPWR 0.22176f
C2381 a_4516_18884# a_4604_18840# 0.28563f
C2382 a_16500_21640# a_16948_21640# 0.01328f
C2383 _399_.A1 a_50196_22805# 0.4875f
C2384 _304_.B a_44028_22020# 0.00485f
C2385 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I 0.01482f
C2386 _424_.B1 _417_.Z 0.04089f
C2387 _285_.Z a_37386_31048# 0.00898f
C2388 a_4068_29860# VPWR 0.21569f
C2389 a_65668_27912# vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I 0.00186f
C2390 a_39264_18147# a_40244_18180# 0.00239f
C2391 a_45800_30345# VPWR 0.18775f
C2392 a_65668_15748# a_65532_15271# 0.00168f
C2393 a_55900_11000# VPWR 0.31436f
C2394 a_39772_26247# a_39684_26344# 0.28563f
C2395 _355_.C a_18044_29816# 0.00238f
C2396 _324_.C _452_.Q 0.01198f
C2397 _351_.ZN a_24080_25227# 0.00336f
C2398 a_63964_15704# a_64412_15704# 0.0131f
C2399 a_23627_27967# a_23920_27555# 0.49319f
C2400 _355_.C _455_.Q 1.31054f
C2401 a_67460_15748# a_67100_15704# 0.08674f
C2402 _452_.Q a_40220_20408# 0.03465f
C2403 _474_.Q a_49448_20072# 0.04886f
C2404 a_17484_27815# VPWR 0.32772f
C2405 _400_.ZN a_44961_27912# 0.07734f
C2406 _260_.A2 a_41476_24776# 0.0342f
C2407 _229_.I vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.11814f
C2408 a_61164_23111# a_61076_23208# 0.28563f
C2409 a_33724_2727# a_33636_2824# 0.28563f
C2410 _419_.A4 _475_.Q 0.09459f
C2411 a_61052_9432# a_61500_9432# 0.0131f
C2412 a_63204_9476# a_62844_9432# 0.08717f
C2413 _424_.A2 _421_.B 0.00212f
C2414 a_14596_1256# a_15044_1256# 0.01328f
C2415 a_4156_7864# a_4604_7864# 0.01222f
C2416 a_64772_4772# a_65220_4772# 0.01328f
C2417 a_65668_3204# a_66116_3204# 0.01328f
C2418 _330_.A1 a_37964_18191# 0.03524f
C2419 _243_.ZN a_58140_26680# 0.00316f
C2420 a_4156_13703# a_4940_13703# 0.00443f
C2421 a_5276_29383# a_5724_29383# 0.0131f
C2422 _351_.A2 a_26160_27165# 0.00318f
C2423 a_6172_30951# a_6084_31048# 0.28563f
C2424 _409_.ZN _397_.A4 0.0159f
C2425 a_12356_1636# VPWR 0.20348f
C2426 _459_.CLK a_22996_25156# 0.00676f
C2427 a_61972_13800# a_62060_12135# 0.00151f
C2428 _384_.ZN _284_.A2 0.0316f
C2429 _284_.ZN _402_.A1 2.07421f
C2430 a_59396_12612# a_59036_12568# 0.08707f
C2431 a_51240_20452# a_51912_20452# 0.00488f
C2432 _243_.B2 VPWR 0.59125f
C2433 _325_.A2 a_42896_18504# 0.02199f
C2434 a_63616_31128# vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN 0.01578f
C2435 a_49764_31048# _392_.A2 0.00245f
C2436 a_61276_1159# VPWR 0.32517f
C2437 a_45696_20072# a_46084_19759# 0.00393f
C2438 a_64636_1159# a_64996_1256# 0.08717f
C2439 _350_.A2 _294_.A2 0.04091f
C2440 _395_.A1 a_48308_23588# 0.01078f
C2441 a_1020_19975# VPWR 0.30073f
C2442 a_47076_11044# a_47524_11044# 0.01328f
C2443 _474_.CLK a_55252_20072# 0.03113f
C2444 _435_.A3 a_37472_24419# 0.00129f
C2445 a_37444_25156# a_37084_25112# 0.08663f
C2446 a_2364_18407# VPWR 0.30029f
C2447 a_4964_1636# a_4828_1159# 0.00168f
C2448 a_1020_1592# a_1020_1159# 0.05841f
C2449 a_32828_1592# a_33276_1592# 0.01288f
C2450 a_36772_1636# a_36860_1592# 0.28563f
C2451 a_34716_20937# a_34732_19975# 0.0019f
C2452 _371_.A2 _371_.A3 0.72293f
C2453 _281_.ZN _427_.B2 0.03268f
C2454 a_43492_27912# a_43940_27912# 0.01328f
C2455 a_42596_27912# _330_.A1 0.00863f
C2456 _336_.A1 _336_.Z 0.71514f
C2457 a_27228_26247# VPWR 0.3279f
C2458 _412_.A1 a_52988_26680# 0.00495f
C2459 a_61276_1592# a_61276_1159# 0.05841f
C2460 a_22212_2824# a_22076_1592# 0.00154f
C2461 _284_.B hold2.I 1.76928f
C2462 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I a_61388_16839# 0.00118f
C2463 a_23980_21976# VPWR 0.31436f
C2464 hold1.Z _447_.Q 0.02456f
C2465 _337_.A3 a_26468_27912# 0.01304f
C2466 a_33948_18840# a_34396_18840# 0.012f
C2467 _433_.ZN a_42168_22504# 0.01478f
C2468 a_41340_2727# VPWR 0.3153f
C2469 a_62420_13800# VPWR 0.20622f
C2470 a_17036_26247# a_17484_26247# 0.0131f
C2471 a_2812_26247# a_3172_26344# 0.08717f
C2472 _412_.A1 _398_.C 0.27785f
C2473 a_44028_22020# VPWR 0.00979f
C2474 _474_.CLK a_54332_20408# 0.01193f
C2475 a_10204_29816# VPWR 0.33263f
C2476 a_62644_16936# a_62620_15704# 0.0016f
C2477 a_2812_10567# VPWR 0.30213f
C2478 vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN _245_.I1 0.13577f
C2479 a_9084_30951# uio_oe[6] 0.00293f
C2480 a_30812_15271# a_31172_15368# 0.08717f
C2481 _452_.CLK a_45732_18884# 0.04086f
C2482 a_28796_23111# VPWR 0.31467f
C2483 _439_.ZN a_41440_23208# 0.00872f
C2484 _424_.A2 _384_.A3 0.12841f
C2485 _441_.ZN _430_.ZN 0.0102f
C2486 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN 0.22738f
C2487 a_59172_26724# VPWR 0.20895f
C2488 hold2.I a_43245_24373# 0.00198f
C2489 a_44700_2727# a_45060_2824# 0.08717f
C2490 _397_.A2 _397_.A1 1.23083f
C2491 a_42392_19243# VPWR 0.75468f
C2492 a_66988_16839# a_66900_16936# 0.28563f
C2493 vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN a_59260_23111# 0.00699f
C2494 a_64412_9432# a_64412_8999# 0.05841f
C2495 a_21428_23588# a_21068_23544# 0.08707f
C2496 a_64860_18407# a_65308_18407# 0.012f
C2497 _355_.C a_22964_27967# 0.00121f
C2498 a_3708_25112# a_4156_25112# 0.0131f
C2499 _416_.A3 a_47552_19715# 0.00111f
C2500 a_1468_13703# a_1380_13800# 0.28563f
C2501 a_27924_20452# a_28372_20452# 0.01328f
C2502 a_26580_20452# a_26220_20408# 0.08717f
C2503 _359_.B _352_.A2 0.00244f
C2504 _395_.A1 _330_.A1 0.32497f
C2505 _319_.A3 a_35504_18955# 0.00319f
C2506 a_62532_18504# a_62532_17316# 0.05841f
C2507 a_36212_23588# VPWR 0.13018f
C2508 _359_.B _284_.ZN 0.32396f
C2509 a_2812_16839# a_2724_16936# 0.28563f
C2510 a_35068_1592# a_35204_1256# 0.00168f
C2511 a_18492_1592# VPWR 0.30281f
C2512 a_62756_12612# a_62396_12568# 0.08707f
C2513 a_65892_12612# a_66340_12612# 0.01328f
C2514 _304_.B a_42236_27815# 0.00379f
C2515 _325_.B a_43400_18909# 0.00736f
C2516 _325_.A1 a_41188_18840# 0.22886f
C2517 _398_.C a_51968_26724# 0.00979f
C2518 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN rst_n 0.15659f
C2519 a_37291_29535# uo_out[7] 0.00547f
C2520 _371_.A2 a_27868_28776# 0.00371f
C2521 a_65532_15271# a_65892_15368# 0.0869f
C2522 _218_.ZN _417_.Z 0.69427f
C2523 _417_.A2 a_47776_20893# 0.00173f
C2524 a_49204_12232# a_49292_10567# 0.00151f
C2525 _304_.A1 a_39178_23208# 0.01452f
C2526 a_62868_12232# a_62844_11000# 0.0016f
C2527 a_11908_1636# a_11772_1159# 0.00168f
C2528 a_39548_1592# a_40220_1592# 0.00544f
C2529 _474_.CLK a_54088_22895# 0.00224f
C2530 a_3620_26724# a_3708_26680# 0.28563f
C2531 _304_.B _284_.B 0.19303f
C2532 _400_.ZN _281_.ZN 0.00105f
C2533 a_66676_10664# a_67124_10664# 0.01328f
C2534 _435_.ZN _441_.A3 0.15459f
C2535 a_36188_1159# a_36636_1159# 0.0131f
C2536 _452_.CLK a_35492_20072# 0.01135f
C2537 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN 0.12396f
C2538 _237_.A1 _258_.I 0.02326f
C2539 _371_.ZN a_28556_29167# 0.00837f
C2540 a_4068_20452# VPWR 0.2157f
C2541 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN 0.03577f
C2542 _360_.ZN _460_.D 0.52973f
C2543 _388_.B a_43716_31048# 0.02058f
C2544 a_63740_2727# VPWR 0.31143f
C2545 a_51556_12612# VPWR 0.20622f
C2546 _330_.A1 _442_.ZN 0.02812f
C2547 a_66116_2824# a_66204_1159# 0.0027f
C2548 _417_.A2 _395_.A3 0.0207f
C2549 _452_.Q a_40332_21543# 0.01921f
C2550 a_3708_29383# a_3620_29480# 0.28563f
C2551 a_32516_20072# VPWR 0.20348f
C2552 a_40132_15368# a_40580_15368# 0.01328f
C2553 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN a_66764_20408# 0.00218f
C2554 a_65644_23544# vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I 0.00329f
C2555 a_3708_15704# a_3708_15271# 0.05841f
C2556 _319_.A2 _448_.D 0.0095f
C2557 a_64300_10567# VPWR 0.34599f
C2558 a_42236_15271# a_42148_15368# 0.28563f
C2559 a_64412_17272# a_64436_16936# 0.00172f
C2560 a_36636_21543# a_36996_21640# 0.08674f
C2561 a_26468_23208# VPWR 0.23302f
C2562 a_43580_15271# a_44028_15271# 0.0131f
C2563 uio_in[1] uio_in[0] 0.03809f
C2564 a_52512_19715# a_52408_19759# 0.10745f
C2565 a_34708_29860# uo_out[4] 0.01602f
C2566 _336_.A2 VPWR 2.02131f
C2567 _451_.Q a_38644_19368# 0.06672f
C2568 a_56124_2727# a_56036_2824# 0.28563f
C2569 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I a_57244_27815# 0.03106f
C2570 a_15156_22020# a_15604_22020# 0.01328f
C2571 _327_.Z a_38788_20072# 0.00172f
C2572 a_39772_19975# a_40132_20072# 0.0869f
C2573 a_67548_17272# a_67996_17272# 0.01222f
C2574 a_62084_15748# VPWR 0.22733f
C2575 _284_.ZN _495_.I 0.00476f
C2576 _311_.Z a_36860_23111# 0.0045f
C2577 _416_.A1 _324_.B 0.0389f
C2578 a_21764_23208# a_21852_21543# 0.00151f
C2579 a_6084_1256# VPWR 0.20348f
C2580 a_7092_31048# VPWR 0.22417f
C2581 a_25236_23588# a_24876_23544# 0.08717f
C2582 a_27924_23588# a_28372_23588# 0.01328f
C2583 a_36996_1256# a_37444_1256# 0.01328f
C2584 a_2276_4772# VPWR 0.20634f
C2585 a_20084_25156# a_19724_25112# 0.08707f
C2586 a_58252_16839# a_58612_16936# 0.08674f
C2587 a_65868_13703# a_66316_13703# 0.0131f
C2588 a_16252_2727# a_16700_2727# 0.0131f
C2589 _268_.A1 a_52640_29860# 0.00494f
C2590 a_51980_13703# a_52340_13800# 0.08707f
C2591 _349_.A4 a_26970_29480# 0.00264f
C2592 a_36548_26344# _444_.D 0.00481f
C2593 a_38764_16839# a_39124_16936# 0.08707f
C2594 a_56012_10567# a_56036_9476# 0.0016f
C2595 a_45732_10664# a_45732_9476# 0.05841f
C2596 _327_.A2 a_41188_18840# 0.16047f
C2597 a_32292_1636# VPWR 0.22423f
C2598 a_42012_1592# a_42148_1256# 0.00168f
C2599 a_64076_16839# VPWR 0.31594f
C2600 a_3172_1636# a_2812_1592# 0.08707f
C2601 _447_.Q _301_.A1 0.97762f
C2602 _260_.A1 _304_.ZN 0.06907f
C2603 a_42236_27815# VPWR 0.31133f
C2604 _450_.D a_43328_18559# 0.00205f
C2605 a_1380_29860# a_1828_29860# 0.01328f
C2606 a_61860_27912# a_61948_26247# 0.00151f
C2607 a_54916_21640# VPWR 0.20897f
C2608 _447_.Q a_39236_20072# 0.00228f
C2609 a_1380_17316# a_1020_17272# 0.08717f
C2610 a_3172_17316# a_3620_17316# 0.01328f
C2611 a_55252_23588# clk 0.00645f
C2612 a_35204_31048# uo_out[4] 0.00178f
C2613 a_46492_1592# a_46940_1592# 0.01288f
C2614 a_53212_11000# a_53660_11000# 0.01288f
C2615 a_52116_16936# a_52564_16936# 0.01328f
C2616 a_57156_11044# a_57244_11000# 0.28563f
C2617 _330_.A1 a_36636_17272# 0.00453f
C2618 _459_.Q _363_.Z 0.29129f
C2619 a_31484_30951# _223_.I 0.03694f
C2620 _294_.A2 _334_.A1 0.26148f
C2621 _230_.I ui_in[3] 0.00176f
C2622 a_52228_19368# a_53100_18407# 0.00107f
C2623 _284_.B VPWR 1.93674f
C2624 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN 0.61336f
C2625 _346_.A2 VPWR 1.32167f
C2626 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN a_65072_29860# 0.04776f
C2627 a_66787_30600# vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN 0.00292f
C2628 a_14796_27815# a_15244_27815# 0.0131f
C2629 _336_.A2 a_28903_24776# 0.00435f
C2630 a_23220_20452# VPWR 0.20692f
C2631 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I 0.00693f
C2632 a_37444_25156# _444_.D 0.01303f
C2633 a_2276_15748# a_2364_15704# 0.28563f
C2634 _268_.A1 _274_.A3 0.842f
C2635 _276_.A2 _274_.A1 0.00976f
C2636 a_48172_18840# a_48196_17316# 0.00131f
C2637 a_57692_12568# VPWR 0.32364f
C2638 a_17060_2824# a_17508_2824# 0.01328f
C2639 a_14684_29383# a_15044_29480# 0.08717f
C2640 a_54556_21543# a_54468_21640# 0.28563f
C2641 a_58388_10664# VPWR 0.23601f
C2642 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I 0.6482f
C2643 a_3260_8999# a_3172_9096# 0.28563f
C2644 a_4156_7431# a_4068_7528# 0.28563f
C2645 a_57244_27815# vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.00306f
C2646 a_43750_23544# a_44162_24120# 0.4995f
C2647 a_5388_5863# a_5300_5960# 0.28563f
C2648 a_52988_15271# a_53572_15368# 0.01675f
C2649 a_61836_25515# vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I 0.00847f
C2650 a_64860_4295# a_64772_4392# 0.28563f
C2651 _452_.CLK a_43664_17317# 0.00387f
C2652 _402_.A1 a_46356_24072# 0.30697f
C2653 _430_.ZN _437_.ZN 0.13624f
C2654 a_31620_15368# VPWR 0.20348f
C2655 vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I 0.07284f
C2656 vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I 0.02911f
C2657 _397_.A1 _330_.A1 0.03775f
C2658 a_21876_22020# a_22548_22020# 0.00347f
C2659 _268_.A2 _258_.ZN 0.00469f
C2660 a_67100_2727# a_67460_2824# 0.08674f
C2661 a_35068_15271# VPWR 0.3552f
C2662 a_1380_14180# a_1020_14136# 0.08717f
C2663 a_3172_14180# a_3620_14180# 0.01328f
C2664 _363_.Z _461_.D 0.13147f
C2665 a_62196_26724# VPWR 0.20665f
C2666 a_32476_29167# VPWR 0.396f
C2667 a_67460_17316# VPWR 0.20622f
C2668 a_31284_23588# a_30924_23544# 0.0869f
C2669 a_4940_7431# VPWR 0.31945f
C2670 a_28484_1256# VPWR 0.20348f
C2671 a_65308_4295# VPWR 0.30378f
C2672 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN a_58588_21543# 0.00639f
C2673 a_62956_13703# a_62868_13800# 0.28563f
C2674 a_59397_26344# VPWR 0.58279f
C2675 _441_.ZN _441_.A3 0.13938f
C2676 _459_.CLK _294_.ZN 0.34608f
C2677 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN 0.0354f
C2678 a_31708_17272# a_31708_16839# 0.05841f
C2679 a_11091_30644# VPWR 0.18981f
C2680 a_35652_17316# a_35628_16839# 0.00172f
C2681 a_49740_16839# a_49652_16936# 0.28563f
C2682 a_62084_18504# VPWR 0.20348f
C2683 a_24316_26247# a_24228_26344# 0.28563f
C2684 _337_.ZN a_30388_28776# 0.10995f
C2685 a_1828_23208# a_1828_22020# 0.05841f
C2686 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_56124_27815# 0.00109f
C2687 a_8636_1159# a_8996_1256# 0.08717f
C2688 a_52876_12135# a_53324_12135# 0.01288f
C2689 a_66876_12568# a_66764_12135# 0.02634f
C2690 a_45956_1636# VPWR 0.20348f
C2691 a_43828_16936# VPWR 0.20665f
C2692 _442_.ZN a_39860_25156# 0.00621f
C2693 _452_.CLK a_37444_26724# 0.01904f
C2694 _294_.A2 a_35652_31048# 0.00118f
C2695 a_1828_29480# a_2276_29480# 0.01328f
C2696 a_9668_1636# a_10116_1636# 0.01328f
C2697 a_23980_23544# a_24092_23111# 0.02634f
C2698 _427_.ZN a_53884_20408# 0.00393f
C2699 _265_.ZN a_43296_28733# 0.00122f
C2700 a_41440_28363# a_43003_28409# 0.41635f
C2701 a_8100_29860# a_8772_29860# 0.00347f
C2702 a_31172_17316# a_30812_17272# 0.08707f
C2703 a_8548_2824# VPWR 0.22888f
C2704 a_50748_11000# a_50636_10567# 0.02634f
C2705 a_53796_1636# a_53436_1592# 0.08707f
C2706 _359_.B _223_.ZN 0.00154f
C2707 _474_.D VPWR 0.55868f
C2708 _434_.ZN a_38131_22804# 0.00201f
C2709 a_15244_24679# a_15692_24679# 0.0131f
C2710 a_17472_28363# a_18028_28777# 0.8399f
C2711 _378_.ZN a_18400_28733# 0.01625f
C2712 a_58588_1159# a_59036_1159# 0.0131f
C2713 a_66676_20452# a_66764_20408# 0.28563f
C2714 a_53548_18407# a_53460_18504# 0.28563f
C2715 a_62084_15368# VPWR 0.20897f
C2716 a_49056_29977# VPWR 0.00217f
C2717 a_67100_18840# a_67548_18840# 0.01222f
C2718 a_54356_18504# VPWR 0.20789f
C2719 a_18380_25112# VPWR 0.3356f
C2720 _304_.B a_52360_26355# 0.04875f
C2721 a_34160_20523# VPWR 1.14106f
C2722 a_28124_30600# VPWR 0.37039f
C2723 a_4940_12135# VPWR 0.31945f
C2724 _378_.I a_17932_27815# 0.00169f
C2725 a_35652_15748# a_36100_15748# 0.01328f
C2726 a_32068_15748# a_32156_15704# 0.28563f
C2727 a_20060_2727# a_20196_1636# 0.00154f
C2728 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN a_56796_15271# 0.01919f
C2729 _397_.A1 a_48988_26369# 0.00186f
C2730 _379_.A2 uio_out[5] 0.58739f
C2731 _427_.A2 a_52920_22760# 0.06045f
C2732 _474_.CLK a_55744_22505# 0.00134f
C2733 clkbuf_1_0__f_clk.I _447_.Q 0.00114f
C2734 _459_.CLK a_22636_29383# 0.00421f
C2735 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN 0.00107f
C2736 a_29244_21543# a_29268_20452# 0.0016f
C2737 _452_.CLK a_41004_16839# 0.00239f
C2738 a_2364_15704# VPWR 0.30029f
C2739 _250_.B a_62396_27815# 0.03177f
C2740 a_40668_20408# _327_.Z 0.00237f
C2741 a_54020_15368# VPWR 0.20348f
C2742 VPWR ui_in[6] 0.00108f
C2743 a_42896_18504# a_43824_18147# 1.16391f
C2744 _432_.ZN a_40973_24776# 0.00406f
C2745 a_54192_22851# _427_.ZN 0.0032f
C2746 a_25236_22020# a_25324_21976# 0.28563f
C2747 a_53076_24776# clk 0.00108f
C2748 a_28820_22020# a_29268_22020# 0.01328f
C2749 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN VPWR 0.81567f
C2750 a_47052_16839# a_47500_16839# 0.01288f
C2751 a_45732_14180# a_45372_14136# 0.08707f
C2752 _237_.A1 _255_.ZN 0.05658f
C2753 a_38764_16839# VPWR 0.31547f
C2754 a_50884_1256# VPWR 0.20981f
C2755 a_36300_23544# a_36748_23544# 0.01255f
C2756 a_26556_30951# a_26468_31048# 0.28563f
C2757 vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I 0.01427f
C2758 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN 0.00168f
C2759 a_59396_1256# a_59844_1256# 0.01328f
C2760 a_59732_13800# a_60180_13800# 0.01328f
C2761 a_38428_2727# a_39100_2727# 0.00544f
C2762 _359_.ZN a_33148_25641# 0.00385f
C2763 a_41048_17341# a_42572_16839# 0.0011f
C2764 a_19716_29977# VPWR 0.00272f
C2765 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN 0.0216f
C2766 _230_.I _267_.A2 0.01908f
C2767 a_36996_17316# VPWR 0.20578f
C2768 a_19524_23208# a_19636_22020# 0.02666f
C2769 _268_.A1 _324_.C 0.08905f
C2770 a_35088_20893# a_34716_20937# 0.10745f
C2771 a_52092_1592# VPWR 0.3289f
C2772 a_20060_1159# a_19972_1256# 0.28563f
C2773 a_50188_12135# a_50100_12232# 0.28563f
C2774 _313_.ZN a_33276_23111# 0.00321f
C2775 a_33376_23659# a_33724_23111# 0.0074f
C2776 _229_.I a_60059_28776# 0.00928f
C2777 a_63740_12568# a_63764_12232# 0.00172f
C2778 a_23084_25112# a_23108_24776# 0.00172f
C2779 a_11460_29860# a_11548_29816# 0.28563f
C2780 a_15044_29860# a_15492_29860# 0.01328f
C2781 a_37532_17272# a_37980_17272# 0.012f
C2782 _402_.A1 a_46620_22504# 0.00142f
C2783 _358_.A3 a_33164_24679# 0.00393f
C2784 _474_.CLK _381_.Z 0.05184f
C2785 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_57604_14180# 0.00516f
C2786 a_67324_11000# a_67772_11000# 0.01288f
C2787 a_57692_11000# a_57580_10567# 0.02634f
C2788 a_45088_29123# VPWR 0.5078f
C2789 a_56708_1636# a_56796_1592# 0.28563f
C2790 a_60292_1636# a_60740_1636# 0.01328f
C2791 a_30724_2824# VPWR 0.20968f
C2792 _304_.B _474_.Q 0.03434f
C2793 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN 1.25018f
C2794 a_25884_23111# a_26556_23111# 0.00544f
C2795 a_4940_23111# a_5300_23208# 0.08674f
C2796 a_67741_30600# _249_.A2 0.00145f
C2797 a_17484_24679# a_17844_24776# 0.08717f
C2798 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_56964_26724# 0.58563f
C2799 a_2724_9476# VPWR 0.20782f
C2800 a_54244_2824# a_54244_1636# 0.05841f
C2801 a_50436_2824# a_50300_1592# 0.00154f
C2802 a_9892_2824# a_9980_1159# 0.0027f
C2803 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN _248_.B1 0.13937f
C2804 a_51556_14180# VPWR 0.20348f
C2805 a_5388_18407# a_5300_18504# 0.28563f
C2806 a_37532_26680# a_37532_26247# 0.05841f
C2807 a_52360_26355# VPWR 1.10758f
C2808 a_29351_28293# _371_.A3 0.00117f
C2809 _397_.A2 _389_.ZN 0.53584f
C2810 a_2724_31048# a_2724_29860# 0.05841f
C2811 a_32292_26344# VPWR 0.20688f
C2812 a_26916_31048# a_26427_29977# 0.03071f
C2813 a_15492_29480# VPWR 0.21284f
C2814 a_66316_12135# VPWR 0.32291f
C2815 _351_.ZN _457_.D 0.0066f
C2816 a_61940_29076# VPWR 0.00417f
C2817 a_39460_2824# a_39908_2824# 0.01328f
C2818 a_27004_2727# a_27140_1636# 0.00154f
C2819 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN 0.10101f
C2820 a_2276_24776# VPWR 0.20634f
C2821 _454_.Q _351_.ZN 0.00639f
C2822 a_67012_7528# VPWR 0.20348f
C2823 _281_.A1 _427_.ZN 0.14733f
C2824 a_18760_29032# a_19140_29612# 0.00257f
C2825 a_27812_21640# a_27924_20452# 0.02666f
C2826 a_1468_19975# a_1828_20072# 0.08717f
C2827 a_41252_15748# VPWR 0.20909f
C2828 _424_.B1 _424_.ZN 0.07915f
C2829 _255_.I a_59348_29076# 0.00281f
C2830 a_56684_23544# a_56572_23111# 0.02634f
C2831 _294_.ZN uo_out[7] 0.625f
C2832 _362_.ZN uo_out[6] 0.15188f
C2833 a_54444_18407# vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN 0.00894f
C2834 a_46180_9476# a_46628_9476# 0.01328f
C2835 _311_.A2 a_34980_22895# 0.50183f
C2836 a_31284_22020# a_30924_21976# 0.0869f
C2837 _260_.ZN a_44028_22020# 0.00159f
C2838 a_52092_14136# a_52540_14136# 0.012f
C2839 _474_.D _424_.B2 0.02652f
C2840 _337_.A3 _457_.D 0.00166f
C2841 a_64884_26724# a_64972_26680# 0.28563f
C2842 a_932_12612# a_1020_12568# 0.28563f
C2843 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I VPWR 0.87358f
C2844 a_50860_18407# a_50884_17316# 0.0016f
C2845 _435_.ZN _300_.ZN 0.00194f
C2846 _459_.CLK a_22548_28292# 0.00213f
C2847 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I a_61076_23208# 0.00172f
C2848 _399_.A2 _384_.A1 0.01875f
C2849 _447_.Q a_37296_22020# 0.00303f
C2850 _454_.Q _337_.A3 0.00798f
C2851 a_22660_23208# a_22636_21976# 0.0016f
C2852 a_67572_10664# a_67548_9432# 0.0016f
C2853 a_33724_23111# a_33152_22091# 0.00105f
C2854 _340_.ZN a_23627_27967# 0.00185f
C2855 a_26468_23208# a_26580_22020# 0.02666f
C2856 a_49092_17316# VPWR 0.21245f
C2857 _358_.A3 a_31348_25156# 0.01909f
C2858 a_65892_1636# VPWR 0.24003f
C2859 a_30812_1159# a_31396_1256# 0.01675f
C2860 a_46628_12232# a_47076_12232# 0.01328f
C2861 a_58140_12568# a_58052_11044# 0.00151f
C2862 a_31088_30301# _371_.A1 0.00208f
C2863 a_60716_12135# a_61076_12232# 0.08707f
C2864 a_19748_1636# a_19836_1592# 0.28563f
C2865 a_23332_1636# a_23780_1636# 0.01328f
C2866 a_32268_23544# a_32292_23208# 0.00172f
C2867 a_21852_21543# VPWR 0.31389f
C2868 a_17508_29860# a_17596_29816# 0.28563f
C2869 _474_.CLK a_52640_29860# 0.01003f
C2870 a_44744_26355# _284_.B 0.01302f
C2871 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN a_52316_27815# 0.00759f
C2872 _231_.ZN vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN 0.22913f
C2873 a_54556_11000# a_54580_10664# 0.00172f
C2874 a_53124_2824# VPWR 0.20815f
C2875 a_40132_1636# a_39996_1159# 0.00168f
C2876 _474_.Q VPWR 3.57489f
C2877 _427_.B1 _417_.A2 0.00145f
C2878 a_24988_23111# a_24900_23208# 0.28563f
C2879 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I a_61972_20452# 0.00412f
C2880 a_19972_24776# a_20420_24776# 0.01328f
C2881 a_52316_9432# VPWR 0.33981f
C2882 a_61188_2824# a_61188_1636# 0.05841f
C2883 a_57380_2824# a_57244_1592# 0.00154f
C2884 a_59372_14136# VPWR 0.29679f
C2885 a_35540_18504# a_35988_18504# 0.01328f
C2886 _362_.ZN uo_out[5] 0.00104f
C2887 a_60180_12232# VPWR 0.20595f
C2888 a_45732_15748# a_45820_15704# 0.28563f
C2889 a_41788_15704# a_42236_15704# 0.01288f
C2890 a_38316_20408# VPWR 0.31605f
C2891 _416_.A1 _403_.ZN 0.0171f
C2892 _474_.CLK _274_.A3 0.43226f
C2893 a_10876_2727# a_11236_2824# 0.08717f
C2894 a_47388_15704# VPWR 0.29679f
C2895 a_10092_30951# uio_oe[4] 0.00238f
C2896 a_43892_20072# VPWR 0.00407f
C2897 a_63068_19975# a_63516_19975# 0.0131f
C2898 _343_.A2 a_23834_28292# 0.00898f
C2899 _304_.B _395_.A2 0.05857f
C2900 a_34396_18840# a_34308_17316# 0.0027f
C2901 a_51780_9476# a_51868_9432# 0.28563f
C2902 a_57120_31048# ui_in[4] 0.00182f
C2903 a_60180_14180# a_60964_14180# 0.00276f
C2904 _447_.Q a_42154_21236# 0.00307f
C2905 a_1380_20452# a_1828_20452# 0.01328f
C2906 _459_.CLK a_24100_29480# 0.00149f
C2907 _324_.C a_46171_27508# 0.01007f
C2908 _452_.Q a_40108_16839# 0.00558f
C2909 a_63616_31128# VPWR 0.95533f
C2910 a_45284_12612# a_45372_12568# 0.28563f
C2911 a_60828_2727# a_61276_2727# 0.0131f
C2912 a_48868_12612# a_49316_12612# 0.01328f
C2913 _474_.CLK _383_.A2 0.13559f
C2914 a_4852_24776# a_4964_23588# 0.02666f
C2915 a_32292_23208# a_32268_21976# 0.0016f
C2916 a_42236_1159# a_42148_1256# 0.28563f
C2917 a_66204_18840# a_66116_17316# 0.00151f
C2918 a_16252_1159# VPWR 0.33444f
C2919 a_4852_20072# a_5300_20072# 0.01328f
C2920 a_61500_12568# a_61412_11044# 0.00151f
C2921 a_64324_7528# a_64324_6340# 0.05841f
C2922 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN a_61276_19975# 0.00647f
C2923 a_4068_12232# a_4068_11044# 0.05841f
C2924 _300_.A2 a_38340_21327# 0.13878f
C2925 a_65220_5960# a_65220_4772# 0.05841f
C2926 a_66116_4392# a_66116_3204# 0.05841f
C2927 a_19076_21640# VPWR 0.21908f
C2928 a_22352_25987# a_22996_25156# 0.01381f
C2929 _441_.A2 _304_.A1 0.33604f
C2930 _381_.Z _398_.C 0.00511f
C2931 a_53572_17316# a_53660_17272# 0.28563f
C2932 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN 0.01578f
C2933 a_49628_17272# a_50076_17272# 0.01288f
C2934 a_47612_10567# a_47972_10664# 0.08717f
C2935 a_45732_18884# a_45820_18840# 0.28563f
C2936 a_61612_10567# a_62060_10567# 0.01288f
C2937 _370_.B a_32476_29167# 0.00951f
C2938 a_2364_1159# a_2812_1159# 0.0131f
C2939 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN a_64100_27912# 0.00369f
C2940 a_7876_2824# a_7740_1592# 0.00154f
C2941 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I 0.00514f
C2942 _452_.CLK a_42168_22504# 0.02803f
C2943 a_23556_23208# a_24004_23208# 0.01328f
C2944 _424_.A2 _402_.B 0.00273f
C2945 _384_.A1 _424_.A1 0.00243f
C2946 a_63292_9432# VPWR 0.31143f
C2947 a_30140_21543# a_30588_21543# 0.01288f
C2948 a_16500_23588# VPWR 0.20348f
C2949 a_66116_6340# VPWR 0.23643f
C2950 a_17932_21543# a_17844_21640# 0.28563f
C2951 a_51968_20127# VPWR 0.00204f
C2952 a_67908_3204# VPWR 0.21437f
C2953 _388_.B _459_.CLK 0.01379f
C2954 a_66116_2824# a_65980_1592# 0.00154f
C2955 a_46268_13703# VPWR 0.29679f
C2956 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN 0.06803f
C2957 _287_.A2 uo_out[6] 1.90152f
C2958 a_30778_31048# uo_out[7] 0.00119f
C2959 _419_.A4 a_49068_20408# 0.49786f
C2960 a_25232_27165# a_25867_26841# 0.02112f
C2961 a_37084_25112# VPWR 0.31233f
C2962 a_49316_11044# VPWR 0.21035f
C2963 a_49092_15748# a_48732_15704# 0.08707f
C2964 a_61860_2824# a_62308_2824# 0.01328f
C2965 _230_.I vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN 0.00244f
C2966 _245_.Z a_60740_26724# 0.00753f
C2967 _451_.Q _301_.A1 0.09086f
C2968 _441_.ZN _300_.ZN 0.03665f
C2969 _324_.C a_41564_26247# 0.00255f
C2970 a_36060_19369# VPWR 0.39698f
C2971 _451_.Q a_39236_20072# 0.00102f
C2972 a_19612_26247# VPWR 0.3491f
C2973 _284_.B _260_.ZN 0.00412f
C2974 _441_.ZN a_39860_25156# 0.01128f
C2975 a_22300_2727# a_22212_2824# 0.28563f
C2976 a_60740_26724# a_60604_26247# 0.00168f
C2977 _438_.A2 a_35616_24776# 0.00116f
C2978 _267_.A2 a_52068_29480# 0.00246f
C2979 _395_.A2 VPWR 1.31935f
C2980 a_57156_9476# a_57604_9476# 0.01328f
C2981 a_3172_1256# a_3620_1256# 0.01328f
C2982 a_37516_27599# a_37860_27967# 0.00275f
C2983 a_1380_28292# VPWR 0.20348f
C2984 a_3620_31048# a_4068_31048# 0.01328f
C2985 a_64548_14180# a_64188_14136# 0.08707f
C2986 a_15156_20452# a_15244_20408# 0.28563f
C2987 _342_.ZN _454_.Q 0.00341f
C2988 _459_.CLK a_26954_28776# 0.00101f
C2989 a_46984_23588# VPWR 0.52142f
C2990 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I 0.80408f
C2991 a_20732_1592# a_20868_1256# 0.00168f
C2992 a_50996_13800# a_51084_12135# 0.00151f
C2993 _352_.A2 a_24228_26344# 0.00163f
C2994 a_58228_27912# _243_.ZN 0.01269f
C2995 vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN VPWR 0.8951f
C2996 _478_.D a_54824_22045# 0.0026f
C2997 _424_.B1 a_52436_18884# 0.00367f
C2998 a_20379_29977# a_19744_30301# 0.02112f
C2999 a_20672_30301# a_18816_29931# 0.02366f
C3000 _260_.ZN a_43245_24373# 0.00142f
C3001 a_38428_1159# VPWR 0.35728f
C3002 _252_.ZN a_61500_27815# 0.00429f
C3003 a_53212_1159# a_53572_1256# 0.08717f
C3004 _330_.A1 _437_.ZN 0.09768f
C3005 a_52340_12232# a_52452_11044# 0.02666f
C3006 a_932_11044# a_1380_11044# 0.01328f
C3007 _384_.A1 a_54804_23588# 0.00187f
C3008 a_29468_1592# a_29916_1592# 0.01288f
C3009 _336_.Z a_29244_23111# 0.01195f
C3010 a_61388_16839# a_61836_16839# 0.0131f
C3011 a_47972_31048# a_48104_30219# 0.03633f
C3012 _260_.A1 _328_.A2 0.12671f
C3013 a_46848_20893# a_46476_20937# 0.10745f
C3014 a_45920_20523# a_47776_20893# 0.02307f
C3015 _419_.A4 a_48776_20204# 0.02867f
C3016 a_36212_23588# _311_.Z 0.00305f
C3017 _474_.CLK _324_.C 0.21213f
C3018 a_58924_10567# a_58836_10664# 0.28563f
C3019 a_1380_18504# a_1380_17316# 0.05841f
C3020 _459_.CLK a_36284_29167# 0.01775f
C3021 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN VPWR 0.68524f
C3022 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN a_62060_23111# 0.0023f
C3023 a_17396_22020# VPWR 0.20348f
C3024 a_36548_21640# VPWR 0.13849f
C3025 _393_.A3 _381_.Z 0.66856f
C3026 _390_.ZN _397_.A4 0.00265f
C3027 _402_.A1 _470_.D 0.10777f
C3028 a_1916_18840# a_2364_18840# 0.0131f
C3029 a_23980_23544# VPWR 0.31389f
C3030 a_28796_21543# a_29156_21640# 0.08707f
C3031 a_4516_18884# a_4156_18840# 0.08674f
C3032 _467_.D a_17472_28363# 0.00775f
C3033 a_50196_22805# VPWR 0.00723f
C3034 a_68108_13703# VPWR 0.35601f
C3035 a_18492_2727# VPWR 0.31745f
C3036 _399_.A1 a_49405_22805# 0.00352f
C3037 a_40244_21640# a_40132_20452# 0.02666f
C3038 _459_.CLK _362_.B 0.0241f
C3039 a_58116_30344# ui_in[4] 0.00318f
C3040 a_3620_29860# VPWR 0.22347f
C3041 a_48104_30219# VPWR 0.70467f
C3042 _287_.A1 a_33776_29123# 0.00939f
C3043 a_55452_11000# VPWR 0.31436f
C3044 _330_.ZN a_37840_18559# 0.00159f
C3045 a_62172_15704# a_62172_15271# 0.05841f
C3046 a_39324_26247# a_39684_26344# 0.0869f
C3047 _455_.D VPWR 0.37155f
C3048 _355_.C a_17596_29816# 0.03117f
C3049 _452_.Q a_39772_20408# 0.01836f
C3050 _355_.C a_24392_28248# 0.02181f
C3051 a_42778_21812# _325_.B 0.00144f
C3052 a_17036_27815# VPWR 0.32271f
C3053 a_67012_15748# a_67100_15704# 0.28563f
C3054 a_33276_2727# a_33636_2824# 0.08717f
C3055 _457_.D a_27328_25227# 0.00127f
C3056 a_63764_23588# a_64212_23588# 0.01328f
C3057 _397_.A1 _393_.A1 0.03502f
C3058 a_49492_18840# a_49896_18909# 0.41635f
C3059 input9.Z vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.01838f
C3060 a_62756_9476# a_62844_9432# 0.28563f
C3061 _330_.A1 a_38336_18147# 0.06416f
C3062 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN 0.00554f
C3063 a_20396_20408# a_20844_20408# 0.0131f
C3064 a_5724_30951# a_6084_31048# 0.0869f
C3065 _351_.A2 a_24860_27209# 0.06785f
C3066 _324_.C _247_.ZN 0.00292f
C3067 a_11908_1636# VPWR 0.21814f
C3068 a_55004_12568# a_55452_12568# 0.01288f
C3069 a_51240_20452# a_51428_20452# 0.00257f
C3070 a_58948_12612# a_59036_12568# 0.28563f
C3071 _459_.CLK a_22548_25156# 0.00201f
C3072 clkbuf_1_0__f_clk.I _421_.B 0.01418f
C3073 _399_.A2 clk 0.00543f
C3074 _304_.B _427_.A2 0.14071f
C3075 _388_.B a_45596_30951# 0.00199f
C3076 a_45060_31048# a_44632_30206# 0.00638f
C3077 _424_.A2 a_52884_18884# 0.00217f
C3078 a_50068_27508# _395_.A2 0.00289f
C3079 a_25867_26841# a_26152_26841# 0.00277f
C3080 a_10204_29816# a_10340_29480# 0.00168f
C3081 a_64636_1159# a_64548_1256# 0.28563f
C3082 a_49316_31048# _392_.A2 0.00245f
C3083 a_35988_18504# a_36076_16839# 0.00151f
C3084 a_60828_1159# VPWR 0.29679f
C3085 a_55476_12232# a_55452_11000# 0.0016f
C3086 a_68108_20408# VPWR 0.36354f
C3087 a_59284_12232# a_59396_11044# 0.02666f
C3088 a_36996_25156# a_37084_25112# 0.28563f
C3089 _474_.CLK a_54804_20072# 0.02087f
C3090 _390_.ZN a_51956_26183# 0.00155f
C3091 a_1916_18407# VPWR 0.297f
C3092 a_36772_1636# a_36412_1592# 0.08707f
C3093 _371_.A2 a_27004_27815# 0.00383f
C3094 a_42148_27912# _330_.A1 0.00712f
C3095 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_56484_29480# 0.01551f
C3096 clkload0.Z _284_.A2 0.01143f
C3097 a_24764_1159# a_25212_1159# 0.0131f
C3098 a_55476_10664# a_55924_10664# 0.01328f
C3099 a_35092_18504# a_35204_17316# 0.02666f
C3100 _324_.C _265_.ZN 0.36666f
C3101 _230_.I _256_.A2 0.06621f
C3102 a_23532_21976# VPWR 0.31436f
C3103 hold1.Z a_42161_24776# 0.03531f
C3104 _455_.Q a_26916_27912# 0.00353f
C3105 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN 0.85211f
C3106 _251_.ZN a_58276_25156# 0.00495f
C3107 a_27364_21640# a_27812_21640# 0.01328f
C3108 a_40892_2727# VPWR 0.31261f
C3109 a_61972_13800# VPWR 0.20622f
C3110 a_2812_26247# a_2724_26344# 0.28563f
C3111 _474_.CLK a_54692_26344# 0.04648f
C3112 _424_.A2 _417_.Z 0.0344f
C3113 _474_.CLK a_53884_20408# 0.00977f
C3114 a_3620_15368# a_4068_15368# 0.01328f
C3115 a_9756_29816# VPWR 0.32966f
C3116 a_2364_10567# VPWR 0.30029f
C3117 a_30812_15271# a_30724_15368# 0.28563f
C3118 a_8627_30644# uio_oe[6] 0.0422f
C3119 a_28348_23111# VPWR 0.31431f
C3120 _452_.CLK a_42996_18840# 0.00557f
C3121 _439_.ZN a_41216_23208# 0.00692f
C3122 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN 0.03584f
C3123 a_32156_15271# a_32604_15271# 0.0131f
C3124 _439_.ZN _325_.A1 0.53994f
C3125 _397_.A4 a_48580_27508# 0.00164f
C3126 _459_.Q _294_.ZN 0.00481f
C3127 a_58052_26724# VPWR 0.21768f
C3128 a_44700_2727# a_44612_2824# 0.28563f
C3129 hold2.I a_42853_24373# 0.00634f
C3130 _442_.ZN _264_.B 0.00755f
C3131 vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN _231_.I 0.02333f
C3132 _272_.A2 _228_.ZN 0.56971f
C3133 a_48104_30219# _383_.ZN 0.00766f
C3134 a_64772_17316# a_65220_17316# 0.01328f
C3135 a_41188_18840# VPWR 0.79509f
C3136 _267_.ZN a_52756_29076# 0.04951f
C3137 a_66540_16839# a_66900_16936# 0.0869f
C3138 _444_.D VPWR 0.70731f
C3139 a_1916_7431# a_2364_7431# 0.0131f
C3140 a_65308_7864# a_65308_7431# 0.05841f
C3141 a_20980_23588# a_21068_23544# 0.28563f
C3142 a_1020_8999# a_1468_8999# 0.0131f
C3143 a_25572_1256# a_26020_1256# 0.01328f
C3144 a_17036_23544# a_17484_23544# 0.01288f
C3145 a_2812_5863# a_3260_5863# 0.0131f
C3146 a_66204_6296# a_66204_5863# 0.05841f
C3147 _416_.A3 a_47259_20127# 0.00235f
C3148 a_1020_13703# a_1380_13800# 0.08717f
C3149 a_3708_4295# a_4156_4295# 0.0131f
C3150 a_67100_4728# a_67100_4295# 0.05841f
C3151 a_4828_2727# a_5276_2727# 0.0131f
C3152 a_54668_13703# a_55116_13703# 0.01288f
C3153 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _409_.ZN 0.00625f
C3154 _452_.CLK _475_.D 0.00869f
C3155 a_36884_16936# a_36860_15271# 0.00134f
C3156 a_26132_20452# a_26220_20408# 0.28563f
C3157 a_16252_29383# a_16700_29383# 0.01222f
C3158 hold2.Z _435_.A3 0.04195f
C3159 a_34939_23705# VPWR 0.38699f
C3160 a_2364_16839# a_2724_16936# 0.08717f
C3161 a_18044_1592# VPWR 0.30075f
C3162 a_52540_12568# a_52428_12135# 0.02634f
C3163 a_7628_30951# a_8627_30644# 0.00646f
C3164 a_62308_12612# a_62396_12568# 0.28563f
C3165 _427_.A2 VPWR 0.89196f
C3166 _304_.B a_41228_27815# 0.03324f
C3167 a_36284_29167# uo_out[7] 0.00525f
C3168 _371_.A2 a_27460_28776# 0.00371f
C3169 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN a_51084_28248# 0.00165f
C3170 a_51196_21543# VPWR 0.32261f
C3171 a_66228_12232# a_66340_11044# 0.02666f
C3172 _252_.ZN a_59036_26247# 0.01009f
C3173 a_65532_15271# a_65444_15368# 0.28563f
C3174 a_49852_11000# a_50300_11000# 0.01288f
C3175 a_40916_16936# a_41364_16936# 0.01328f
C3176 _474_.CLK a_54192_22851# 0.00326f
C3177 a_43268_1636# a_43716_1636# 0.01328f
C3178 _383_.A2 _393_.A3 0.0094f
C3179 _252_.ZN a_61860_27912# 0.00211f
C3180 a_67100_15704# a_67236_15368# 0.00168f
C3181 _454_.D VPWR 0.41688f
C3182 a_3620_26724# a_3260_26680# 0.08717f
C3183 a_1020_26680# a_1468_26680# 0.0131f
C3184 _384_.ZN _381_.A2 0.12084f
C3185 _443_.D a_37980_26247# 0.0023f
C3186 _362_.ZN _460_.Q 0.28878f
C3187 _400_.ZN a_46156_25112# 0.00145f
C3188 _362_.B uo_out[7] 0.04333f
C3189 _324_.C _398_.C 0.18626f
C3190 _294_.ZN _461_.D 0.01052f
C3191 _304_.B a_43253_25940# 0.00927f
C3192 _452_.CLK a_34644_20072# 0.00524f
C3193 a_56572_29383# _258_.ZN 0.00519f
C3194 _360_.ZN a_32292_26344# 0.00942f
C3195 _371_.ZN a_28928_29123# 0.00202f
C3196 a_3620_20452# VPWR 0.22347f
C3197 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I 0.59821f
C3198 a_24900_27912# _351_.A2 0.0896f
C3199 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN a_64412_29816# 0.00887f
C3200 _388_.B a_43268_31048# 0.01831f
C3201 _330_.A1 a_39536_26795# 0.03793f
C3202 a_51108_12612# VPWR 0.20627f
C3203 a_63292_2727# VPWR 0.31143f
C3204 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I a_63404_20408# 0.00399f
C3205 vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I 0.01711f
C3206 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I 0.06254f
C3207 a_17396_26344# a_17844_26344# 0.01328f
C3208 _452_.Q _432_.ZN 0.02226f
C3209 a_5636_2824# a_6084_2824# 0.01328f
C3210 a_5724_2727# a_5860_1636# 0.00154f
C3211 a_3260_29383# a_3620_29480# 0.08717f
C3212 a_67884_18407# a_67796_18504# 0.28563f
C3213 a_65196_23544# vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I 0.00163f
C3214 a_32068_20072# VPWR 0.20348f
C3215 a_58476_17272# a_58924_17272# 0.01222f
C3216 a_63852_10567# VPWR 0.31547f
C3217 a_41564_15271# a_42148_15368# 0.01675f
C3218 a_25884_27815# a_25796_27912# 0.28563f
C3219 _319_.A2 a_35716_20072# 0.00716f
C3220 a_25796_23208# VPWR 0.21584f
C3221 a_36636_21543# a_36548_21640# 0.28563f
C3222 _238_.I a_59572_29076# 0.26177f
C3223 a_54356_16936# a_54332_15704# 0.0016f
C3224 a_40244_18180# a_40636_18180# 0.00705f
C3225 a_52024_20083# a_52408_19759# 1.16391f
C3226 a_28036_26724# VPWR 0.20768f
C3227 a_34260_29860# uo_out[4] 0.01727f
C3228 a_52764_27815# a_52900_26724# 0.00154f
C3229 _452_.CLK _317_.A2 0.03872f
C3230 _451_.Q a_39268_18840# 0.3988f
C3231 a_61388_15704# VPWR 0.33694f
C3232 a_39772_19975# a_39684_20072# 0.28563f
C3233 a_55676_2727# a_56036_2824# 0.08717f
C3234 vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I 0.11745f
C3235 a_21516_23544# a_21428_22020# 0.00151f
C3236 a_32964_16936# a_32964_15748# 0.05841f
C3237 a_51668_18504# a_52116_18504# 0.01328f
C3238 a_24788_23588# a_24876_23544# 0.28563f
C3239 a_5636_1256# VPWR 0.20348f
C3240 a_15692_25112# a_16140_25112# 0.01288f
C3241 a_1828_4772# VPWR 0.20348f
C3242 a_19636_25156# a_19724_25112# 0.28563f
C3243 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I 0.86437f
C3244 a_6084_31048# VPWR 0.20996f
C3245 _281_.A1 a_51240_20452# 0.02696f
C3246 a_51980_13703# a_51892_13800# 0.28563f
C3247 _251_.A1 a_59260_26680# 0.00283f
C3248 a_34715_22137# VPWR 0.39703f
C3249 a_58252_16839# a_58164_16936# 0.28563f
C3250 _268_.A1 a_51457_29861# 0.00271f
C3251 a_31372_20408# a_31820_20408# 0.0131f
C3252 vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN VPWR 0.76442f
C3253 a_25100_30951# a_25652_31048# 0.01375f
C3254 a_36100_26344# _444_.D 0.00464f
C3255 _416_.A3 _419_.Z 0.2792f
C3256 _465_.D _379_.A2 0.06246f
C3257 a_38764_16839# a_38676_16936# 0.28563f
C3258 a_31708_1592# VPWR 0.35728f
C3259 a_63628_16839# VPWR 0.31594f
C3260 a_2724_1636# a_2812_1592# 0.28563f
C3261 a_6308_1636# a_6756_1636# 0.01328f
C3262 a_1916_12135# a_2364_12135# 0.0131f
C3263 a_59484_12568# a_59372_12135# 0.02634f
C3264 a_16140_23544# a_16140_23111# 0.05841f
C3265 _447_.Q a_37408_23208# 0.00899f
C3266 a_41228_27815# VPWR 0.34512f
C3267 a_5052_25112# a_4940_24679# 0.02634f
C3268 a_20084_23588# a_20060_23111# 0.00172f
C3269 a_932_17316# a_1020_17272# 0.28563f
C3270 a_54468_21640# VPWR 0.20897f
C3271 a_59732_12232# a_59820_10567# 0.00151f
C3272 a_57156_11044# a_56796_11000# 0.08707f
C3273 a_3708_11000# a_3708_10567# 0.05841f
C3274 _304_.ZN a_43646_21236# 0.00129f
C3275 a_54804_23588# clk 0.00645f
C3276 _352_.ZN a_26668_23544# 0.00135f
C3277 _265_.ZN a_42340_28409# 0.00139f
C3278 a_31484_30951# a_31396_31048# 0.28563f
C3279 a_52228_19368# a_52652_18407# 0.00118f
C3280 a_47164_1159# a_47612_1159# 0.0131f
C3281 a_36100_2824# a_35964_1592# 0.00154f
C3282 a_52228_19368# VPWR 0.82545f
C3283 _257_.B _238_.I 0.18689f
C3284 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I a_57468_16839# 0.00662f
C3285 a_64772_18884# a_65220_18884# 0.01328f
C3286 _336_.A2 a_28679_24776# 0.00549f
C3287 a_22772_20452# VPWR 0.20692f
C3288 _324_.C _393_.A3 0.41272f
C3289 a_36996_25156# _444_.D 0.01306f
C3290 vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I 0.62563f
C3291 a_2276_15748# a_1916_15704# 0.08717f
C3292 a_4068_15748# a_4516_15748# 0.01328f
C3293 a_57244_12568# VPWR 0.32088f
C3294 a_51108_15368# a_51556_15368# 0.01328f
C3295 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I 0.00924f
C3296 a_14684_29383# a_14596_29480# 0.28563f
C3297 a_54108_21543# a_54468_21640# 0.0869f
C3298 a_2812_8999# a_3172_9096# 0.08717f
C3299 a_57940_10664# VPWR 0.21742f
C3300 a_3708_7431# a_4068_7528# 0.08717f
C3301 a_43126_24119# a_44162_24120# 0.00389f
C3302 a_41488_24072# _226_.ZN 0.22827f
C3303 a_52988_15271# a_52900_15368# 0.28563f
C3304 a_4940_5863# a_5300_5960# 0.08674f
C3305 _267_.A1 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.03053f
C3306 a_56124_27815# vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.09918f
C3307 a_64412_4295# a_64772_4392# 0.08717f
C3308 a_61836_25515# a_62560_25112# 0.3026f
C3309 a_38616_24328# _437_.ZN 0.02847f
C3310 a_54556_15271# a_55004_15271# 0.0131f
C3311 a_42853_24373# VPWR 0.00186f
C3312 _399_.ZN _384_.A1 0.01821f
C3313 a_31172_15368# VPWR 0.20348f
C3314 _424_.B1 _412_.B2 0.05999f
C3315 _264_.B _435_.ZN 0.00162f
C3316 a_17932_21976# a_18380_21976# 0.01288f
C3317 a_21876_22020# a_21964_21976# 0.28563f
C3318 _243_.A1 a_59172_27912# 0.00191f
C3319 a_34620_15271# VPWR 0.34708f
C3320 a_67100_2727# a_67012_2824# 0.28563f
C3321 _268_.A2 a_56572_29383# 0.00529f
C3322 a_36076_16839# a_36524_16839# 0.01288f
C3323 a_932_14180# a_1020_14136# 0.28563f
C3324 a_40020_16936# a_39908_15748# 0.02666f
C3325 a_25324_23544# a_25236_22020# 0.00151f
C3326 a_61748_26724# VPWR 0.22884f
C3327 a_67012_17316# VPWR 0.20622f
C3328 a_32848_29123# VPWR 0.18788f
C3329 a_30836_23588# a_30924_23544# 0.28563f
C3330 a_31732_23588# a_32180_23588# 0.01328f
C3331 _251_.A1 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I 0.58811f
C3332 a_32292_23208# a_32380_21543# 0.00151f
C3333 a_4156_7431# VPWR 0.3269f
C3334 a_28036_1256# VPWR 0.20348f
C3335 a_64860_4295# VPWR 0.30145f
C3336 a_47972_1256# a_48420_1256# 0.01328f
C3337 a_48420_13800# a_49204_13800# 0.00276f
C3338 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN clk 0.57734f
C3339 a_27004_2727# a_27676_2727# 0.00544f
C3340 vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN a_56596_18504# 0.00618f
C3341 a_62508_13703# a_62868_13800# 0.08707f
C3342 _371_.ZN uio_out[0] 0.04511f
C3343 a_10540_30951# VPWR 0.32672f
C3344 a_61636_18504# VPWR 0.15208f
C3345 a_20508_23111# a_20532_22020# 0.0016f
C3346 a_49292_16839# a_49652_16936# 0.08663f
C3347 _287_.A2 _460_.Q 0.05126f
C3348 a_8636_1159# a_8548_1256# 0.28563f
C3349 a_52788_10664# a_52900_9476# 0.02666f
C3350 a_23868_26247# a_24228_26344# 0.08663f
C3351 a_43380_16936# VPWR 0.20665f
C3352 a_45508_1636# VPWR 0.20348f
C3353 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_55676_27815# 0.00212f
C3354 vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I 0.01558f
C3355 a_56348_12568# a_56372_12232# 0.00172f
C3356 _355_.C _379_.A2 0.08946f
C3357 vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN a_57492_18884# 0.00164f
C3358 a_27028_23588# a_27004_23111# 0.00172f
C3359 _452_.CLK a_36996_26724# 0.02568f
C3360 a_21068_25112# a_20956_24679# 0.02634f
C3361 a_4156_29816# a_4604_29816# 0.01288f
C3362 _260_.A1 _452_.Q 0.6696f
C3363 a_8100_29860# a_8188_29816# 0.28563f
C3364 a_25792_30301# a_26427_29977# 0.02112f
C3365 a_41440_28363# a_43296_28733# 0.02307f
C3366 _265_.ZN a_41996_28777# 0.28841f
C3367 a_34308_17316# a_34756_17316# 0.01328f
C3368 a_30724_17316# a_30812_17272# 0.28563f
C3369 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN 0.04795f
C3370 a_46404_15368# a_46268_14136# 0.00154f
C3371 a_63964_15271# a_64100_14180# 0.00154f
C3372 a_50212_15368# a_50212_14180# 0.05841f
C3373 _416_.ZN a_47636_18884# 0.00367f
C3374 a_25796_1636# a_25660_1159# 0.00168f
C3375 a_49404_1592# a_49852_1592# 0.01288f
C3376 a_53348_1636# a_53436_1592# 0.28563f
C3377 a_63652_11044# a_64100_11044# 0.01328f
C3378 a_7876_2824# VPWR 0.21435f
C3379 a_50196_21640# VPWR 0.00706f
C3380 a_33860_20072# a_33860_18884# 0.05841f
C3381 a_14796_23111# a_15244_23111# 0.0131f
C3382 a_19035_28409# a_19280_28777# 0.00232f
C3383 a_17472_28363# a_18400_28733# 1.16391f
C3384 a_53100_18407# a_53460_18504# 0.08717f
C3385 a_66676_20452# a_66316_20408# 0.08674f
C3386 a_61636_15368# VPWR 0.20897f
C3387 a_53908_18504# VPWR 0.20862f
C3388 _461_.D a_33140_29860# 0.0018f
C3389 a_17932_25112# VPWR 0.30035f
C3390 _475_.Q _427_.B2 0.00887f
C3391 a_15156_27912# a_15604_27912# 0.01328f
C3392 _325_.A1 _303_.ZN 0.48322f
C3393 a_27668_31048# VPWR 0.39857f
C3394 _393_.A1 _389_.ZN 0.19378f
C3395 a_4156_12135# VPWR 0.3269f
C3396 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN 0.00703f
C3397 a_32068_15748# a_31708_15704# 0.08707f
C3398 _275_.A2 a_52756_29076# 0.01296f
C3399 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN a_56348_15271# 0.00195f
C3400 a_28036_2824# a_28484_2824# 0.01328f
C3401 a_40892_15704# a_41028_15368# 0.00168f
C3402 _397_.A1 a_48560_26369# 0.00142f
C3403 _427_.A2 a_51240_23340# 0.00219f
C3404 a_42684_15704# a_42684_15271# 0.05841f
C3405 _251_.A1 a_63336_29480# 0.1835f
C3406 a_23108_29860# a_23084_29383# 0.00172f
C3407 a_20420_21640# a_20308_20452# 0.02666f
C3408 a_18628_21640# a_18604_20408# 0.0016f
C3409 _275_.ZN _274_.ZN 0.18419f
C3410 _452_.CLK a_40556_16839# 0.00239f
C3411 a_40668_20408# a_40668_19975# 0.05841f
C3412 a_1916_15704# VPWR 0.297f
C3413 a_53572_15368# VPWR 0.22423f
C3414 a_25236_22020# a_24876_21976# 0.08707f
C3415 a_53704_23219# _427_.ZN 0.00624f
C3416 a_45284_14180# a_45372_14136# 0.28563f
C3417 a_56796_15271# VPWR 0.3504f
C3418 a_48868_14180# a_49316_14180# 0.01328f
C3419 a_36636_17272# a_36548_15748# 0.00151f
C3420 a_30924_23544# a_30836_22020# 0.00151f
C3421 a_46964_16936# a_46852_15748# 0.02666f
C3422 a_38316_16839# VPWR 0.33043f
C3423 a_48104_30219# a_49112_29885# 0.02307f
C3424 _328_.A2 a_44276_20072# 0.09445f
C3425 a_26108_30951# a_26468_31048# 0.08674f
C3426 a_50436_1256# VPWR 0.26343f
C3427 a_63292_14136# a_63204_12612# 0.00151f
C3428 _284_.A2 a_50120_26476# 0.00343f
C3429 _359_.ZN a_33520_25597# 0.00207f
C3430 a_56516_26344# a_56828_25940# 0.00685f
C3431 _424_.B2 a_52228_19368# 0.4024f
C3432 a_36548_17316# VPWR 0.20622f
C3433 _301_.Z VPWR 0.5536f
C3434 a_27452_23111# a_27476_22020# 0.0016f
C3435 a_63404_12135# a_63852_12135# 0.01288f
C3436 a_51644_1592# VPWR 0.3289f
C3437 a_19388_1159# a_19972_1256# 0.01675f
C3438 a_55900_1592# a_56036_1256# 0.00168f
C3439 a_49740_12135# a_50100_12232# 0.08707f
C3440 a_12444_1592# a_12892_1592# 0.01288f
C3441 a_22636_23544# a_22660_23208# 0.00172f
C3442 a_12804_29480# a_13252_29480# 0.01328f
C3443 a_62756_27912# a_62644_26724# 0.02666f
C3444 _362_.ZN a_32836_27208# 0.00932f
C3445 a_11460_29860# a_11100_29816# 0.08707f
C3446 _311_.A2 _441_.B 0.09259f
C3447 _325_.A2 _323_.A3 0.60718f
C3448 _436_.B _432_.ZN 0.1972f
C3449 a_21652_29480# a_21540_28292# 0.02666f
C3450 a_49764_31048# _268_.A2 0.00157f
C3451 a_30276_2824# VPWR 0.20348f
C3452 a_56708_1636# a_56348_1592# 0.08707f
C3453 a_44795_29535# VPWR 0.36908f
C3454 _416_.A3 _416_.A2 1.01315f
C3455 a_4940_23111# a_4852_23208# 0.28563f
C3456 a_56404_27208# a_56964_26724# 0.3026f
C3457 a_17484_24679# a_17396_24776# 0.28563f
C3458 a_4940_8999# a_4964_7908# 0.0016f
C3459 a_4852_9096# a_5300_9096# 0.01328f
C3460 a_64324_7528# a_64772_7528# 0.01328f
C3461 a_2276_9476# VPWR 0.20634f
C3462 a_33948_19975# a_34732_19975# 0.00443f
C3463 _441_.ZN _264_.B 0.00825f
C3464 _294_.A2 _296_.ZN 0.00107f
C3465 a_65220_5960# a_65668_5960# 0.01328f
C3466 a_51108_14180# VPWR 0.20353f
C3467 a_35628_18407# a_36076_18407# 0.01255f
C3468 a_66116_4392# a_66564_4392# 0.01328f
C3469 a_4940_18407# a_5300_18504# 0.08674f
C3470 a_35140_26680# a_35204_26344# 0.00102f
C3471 _303_.ZN _327_.A2 0.09069f
C3472 a_31844_26344# VPWR 0.12482f
C3473 a_26916_31048# a_26720_30301# 0.0017f
C3474 a_15044_29480# VPWR 0.20665f
C3475 a_59572_29076# VPWR 1.38216f
C3476 a_65868_12135# VPWR 0.34668f
C3477 a_38564_15748# a_39012_15748# 0.01328f
C3478 _416_.A1 _421_.A1 0.09208f
C3479 a_1828_24776# VPWR 0.20348f
C3480 _454_.Q a_24304_26795# 0.00317f
C3481 a_18760_29032# a_18264_29480# 0.00488f
C3482 a_66564_7528# VPWR 0.20631f
C3483 _438_.A2 _438_.ZN 0.38162f
C3484 a_40804_15748# VPWR 0.20663f
C3485 a_1468_19975# a_1380_20072# 0.28563f
C3486 _395_.A1 _395_.A3 0.00991f
C3487 a_54444_18407# a_54892_18407# 0.012f
C3488 a_53996_18407# vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN 0.00207f
C3489 _409_.ZN _392_.A2 0.08881f
C3490 _311_.A2 a_34586_23208# 0.0113f
C3491 a_30836_22020# a_30924_21976# 0.28563f
C3492 a_31732_22020# a_32180_22020# 0.01328f
C3493 a_44571_26841# VPWR 0.35681f
C3494 _265_.ZN a_43580_27815# 0.00143f
C3495 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN 0.00253f
C3496 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I 0.68481f
C3497 a_6396_1592# a_6532_1256# 0.00168f
C3498 _285_.Z _288_.ZN 0.01524f
C3499 a_2724_12612# a_3172_12612# 0.01328f
C3500 a_49404_2727# a_49852_2727# 0.0131f
C3501 _459_.CLK a_21628_28248# 0.00832f
C3502 a_35914_28776# uo_out[7] 0.00134f
C3503 a_28256_25597# a_27884_25641# 0.10745f
C3504 a_48284_17272# a_48396_16839# 0.02634f
C3505 a_52228_17316# a_52204_16839# 0.00172f
C3506 _447_.Q a_42168_22504# 0.02356f
C3507 a_4604_26680# a_4516_25156# 0.0027f
C3508 a_48644_17316# VPWR 0.21036f
C3509 a_30812_1159# a_30724_1256# 0.28563f
C3510 a_60716_12135# a_60628_12232# 0.28563f
C3511 a_65444_1636# VPWR 0.21633f
C3512 a_19748_1636# a_19388_1592# 0.08707f
C3513 a_17508_29860# a_17148_29816# 0.0869f
C3514 _474_.CLK a_51457_29861# 0.01468f
C3515 _250_.C a_62279_28293# 0.00557f
C3516 a_21404_21543# VPWR 0.31389f
C3517 a_15156_26344# a_15156_25156# 0.05841f
C3518 a_46404_17316# a_46852_17316# 0.01328f
C3519 a_52676_2824# VPWR 0.20815f
C3520 a_50636_10567# a_51084_10567# 0.01288f
C3521 a_63068_1592# a_63652_1636# 0.01675f
C3522 _459_.Q _362_.B 0.88131f
C3523 _257_.B VPWR 0.45209f
C3524 _311_.A2 _300_.A2 0.35275f
C3525 a_52228_27912# a_52676_27912# 0.01328f
C3526 _324_.C _452_.CLK 0.44011f
C3527 a_3172_23208# a_3620_23208# 0.01328f
C3528 a_24540_23111# a_24900_23208# 0.08707f
C3529 a_51868_9432# VPWR 0.31143f
C3530 a_19164_21543# a_19612_21543# 0.01288f
C3531 a_58924_14136# VPWR 0.2963f
C3532 a_20868_2824# a_20956_1159# 0.0027f
C3533 _260_.A2 _452_.Q 0.16127f
C3534 _260_.A1 a_40357_24776# 0.00141f
C3535 a_10452_31048# a_10564_29860# 0.02666f
C3536 a_59332_29816# _257_.B 0.00348f
C3537 a_45732_15748# a_45372_15704# 0.08663f
C3538 a_59732_12232# VPWR 0.20595f
C3539 _452_.CLK _416_.ZN 0.02836f
C3540 a_50436_2824# a_50884_2824# 0.01328f
C3541 a_34844_24679# VPWR 0.37833f
C3542 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_58588_26247# 0.00471f
C3543 a_52744_26031# _412_.ZN 0.02534f
C3544 _412_.B2 a_51016_25940# 0.00815f
C3545 _459_.Q a_32628_26725# 0.03304f
C3546 a_65220_20072# VPWR 0.21513f
C3547 a_10876_2727# a_10788_2824# 0.28563f
C3548 a_46940_15704# VPWR 0.29679f
C3549 _399_.ZN clk 0.00398f
C3550 _424_.A2 _424_.ZN 0.4651f
C3551 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN 0.07726f
C3552 _417_.Z a_49988_21236# 0.39288f
C3553 _436_.B _260_.A1 0.10419f
C3554 a_49628_9432# a_50076_9432# 0.0131f
C3555 a_51780_9476# a_51420_9432# 0.08717f
C3556 _459_.CLK _402_.A1 0.05138f
C3557 a_56260_31048# ui_in[4] 0.0014f
C3558 a_55900_14136# a_56348_14136# 0.0131f
C3559 a_62532_15368# a_62508_13703# 0.00131f
C3560 a_60180_14180# a_60268_14136# 0.28563f
C3561 _459_.CLK a_22996_29480# 0.00728f
C3562 a_62532_30736# VPWR 0.45088f
C3563 _416_.A1 _409_.ZN 0.09844f
C3564 _381_.Z a_50176_26724# 0.00269f
C3565 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I VPWR 0.6969f
C3566 a_20060_24679# a_20084_23588# 0.0016f
C3567 _455_.D a_20980_25156# 0.00198f
C3568 a_15580_1159# VPWR 0.32517f
C3569 a_41788_1159# a_42148_1256# 0.08717f
C3570 a_26244_1636# a_26692_1636# 0.01328f
C3571 _300_.A2 a_37444_21640# 0.00103f
C3572 _378_.I _346_.A2 0.00193f
C3573 a_57492_12232# a_57940_12232# 0.01328f
C3574 _474_.CLK a_54780_26247# 0.01977f
C3575 a_18628_21640# VPWR 0.23378f
C3576 a_54824_22045# a_56236_22505# 0.00393f
C3577 a_53572_17316# a_53212_17272# 0.08663f
C3578 a_22352_25987# a_22548_25156# 0.0017f
C3579 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN 0.7119f
C3580 a_43400_18909# a_44320_19369# 0.00306f
C3581 a_47612_10567# a_47524_10664# 0.28563f
C3582 a_61500_11000# a_61524_10664# 0.00172f
C3583 _370_.B a_32848_29123# 0.00281f
C3584 _424_.A2 a_46356_24072# 0.00117f
C3585 a_62508_21976# vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I 0.00729f
C3586 _400_.ZN _402_.ZN 0.02005f
C3587 a_54604_23263# VPWR 0.00246f
C3588 vgaringosc.workerclkbuff_notouch_.I a_52073_30344# 0.00106f
C3589 _436_.ZN VPWR 0.31733f
C3590 a_31803_24831# a_32096_24419# 0.49319f
C3591 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN rst_n 0.0083f
C3592 vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN VPWR 0.80284f
C3593 a_62844_9432# VPWR 0.31143f
C3594 a_16052_23588# VPWR 0.20348f
C3595 a_65668_6340# VPWR 0.21209f
C3596 a_45820_13703# VPWR 0.29679f
C3597 a_54356_20072# VPWR 0.13219f
C3598 a_17484_21543# a_17844_21640# 0.08717f
C3599 a_65556_23588# clk 0.00657f
C3600 a_62980_20072# a_63428_20072# 0.01328f
C3601 a_67460_3204# VPWR 0.20348f
C3602 _294_.A2 a_29232_29931# 0.02256f
C3603 _276_.A2 vgaringosc.workerclkbuff_notouch_.I 0.10901f
C3604 _355_.C a_30476_23544# 0.00189f
C3605 a_48868_11044# VPWR 0.21134f
C3606 a_48644_15748# a_48732_15704# 0.28563f
C3607 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN a_63105_28293# 0.05851f
C3608 clkbuf_1_0__f_clk.I _402_.B 0.26847f
C3609 a_52228_15748# a_52676_15748# 0.01328f
C3610 a_36636_25112# VPWR 0.29679f
C3611 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I 0.01698f
C3612 vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN a_67996_21976# 0.0053f
C3613 a_40892_2727# a_41028_1636# 0.00154f
C3614 _294_.A2 _335_.ZN 0.08015f
C3615 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN 0.59516f
C3616 _460_.Q a_35008_27533# 0.06158f
C3617 a_36432_19325# VPWR 0.18721f
C3618 a_19164_26247# VPWR 0.33815f
C3619 _451_.Q a_38788_20072# 0.00935f
C3620 a_21852_2727# a_22212_2824# 0.08717f
C3621 a_47802_26724# VPWR 0.01471f
C3622 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I a_61188_20072# 0.00138f
C3623 _359_.B _459_.CLK 6.77688f
C3624 a_932_28292# VPWR 0.22176f
C3625 a_3708_9432# a_3708_8999# 0.05841f
C3626 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I a_67436_19975# 0.00285f
C3627 a_64100_14180# a_64188_14136# 0.28563f
C3628 a_15156_20452# a_14796_20408# 0.08717f
C3629 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN 0.78191f
C3630 a_16500_20452# a_16948_20452# 0.01328f
C3631 _279_.Z _397_.Z 0.09167f
C3632 a_24864_29931# _454_.Q 0.00155f
C3633 _327_.Z a_38852_18884# 0.01334f
C3634 a_51644_12568# a_52092_12568# 0.01288f
C3635 _276_.A2 a_52068_29480# 0.00101f
C3636 _223_.I _358_.A2 0.00267f
C3637 a_20379_29977# a_18816_29931# 0.41622f
C3638 _252_.ZN a_61052_27815# 0.0101f
C3639 hold1.Z _441_.A2 0.05571f
C3640 _260_.ZN a_42853_24373# 0.00114f
C3641 a_53212_1159# a_53124_1256# 0.28563f
C3642 a_37980_1159# VPWR 0.3289f
C3643 _384_.A1 a_54356_23588# 0.05887f
C3644 a_46628_31048# _393_.ZN 0.01245f
C3645 a_45920_20523# a_46476_20937# 0.8399f
C3646 _407_.ZN _395_.A2 0.00718f
C3647 _419_.A4 a_47552_19715# 0.00666f
C3648 a_4852_10664# a_5300_10664# 0.01328f
C3649 _284_.ZN a_40264_30320# 0.04393f
C3650 a_58476_10567# a_58836_10664# 0.08707f
C3651 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I VPWR 0.92085f
C3652 a_13340_1159# a_13788_1159# 0.0131f
C3653 _459_.CLK a_36656_29123# 0.01533f
C3654 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN a_61612_23111# 0.00177f
C3655 a_55340_19975# VPWR 0.31992f
C3656 a_16948_22020# VPWR 0.20348f
C3657 a_37472_24419# a_38616_24328# 0.00981f
C3658 _417_.A2 a_51108_21640# 0.00903f
C3659 a_23532_23544# VPWR 0.31389f
C3660 a_28796_21543# a_28708_21640# 0.28563f
C3661 a_16052_21640# a_16500_21640# 0.01328f
C3662 a_4068_18884# a_4156_18840# 0.28563f
C3663 a_67660_13703# VPWR 0.31431f
C3664 a_18044_2727# VPWR 0.31539f
C3665 _408_.ZN _384_.A3 0.00349f
C3666 vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN a_57940_20452# 0.00631f
C3667 a_3172_29860# VPWR 0.20993f
C3668 a_45904_30180# VPWR 0.39827f
C3669 a_38971_18559# a_39264_18147# 0.49319f
C3670 a_39324_26247# a_39236_26344# 0.28563f
C3671 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN _267_.A2 0.0237f
C3672 a_55004_11000# VPWR 0.31436f
C3673 _287_.A1 a_33483_29535# 0.00978f
C3674 a_65220_15748# a_65084_15271# 0.00168f
C3675 a_20844_26680# VPWR 0.32748f
C3676 _495_.I _459_.CLK 0.15223f
C3677 a_63516_15704# a_63964_15704# 0.0131f
C3678 a_67012_15748# a_66652_15704# 0.0869f
C3679 _402_.A1 uo_out[7] 0.28267f
C3680 a_16588_27815# VPWR 0.29679f
C3681 _260_.A2 a_40357_24776# 0.00214f
C3682 a_53212_29816# vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN 0.0011f
C3683 a_33276_2727# a_33188_2824# 0.28563f
C3684 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I _251_.ZN 0.00435f
C3685 _399_.ZN _416_.A3 0.00124f
C3686 a_60604_9432# a_61052_9432# 0.0131f
C3687 a_62756_9476# a_62396_9432# 0.08717f
C3688 a_4604_23544# a_5052_23544# 0.01222f
C3689 a_3708_7864# a_4156_7864# 0.0131f
C3690 a_14148_1256# a_14596_1256# 0.01328f
C3691 a_4604_6296# a_5052_6296# 0.01222f
C3692 a_64324_4772# a_64772_4772# 0.01328f
C3693 a_28804_27208# _355_.B 0.0091f
C3694 _324_.C a_43668_19668# 0.39334f
C3695 a_3708_13703# a_4156_13703# 0.0131f
C3696 a_65220_3204# a_65668_3204# 0.01328f
C3697 _459_.CLK a_32144_26724# 0.00812f
C3698 a_5724_30951# a_5636_31048# 0.28563f
C3699 a_4828_29383# a_5276_29383# 0.0131f
C3700 _480_.Q _402_.A1 0.06058f
C3701 _351_.A2 a_25232_27165# 0.03071f
C3702 a_58948_12612# a_58588_12568# 0.08707f
C3703 a_61524_13800# a_61612_12135# 0.00151f
C3704 a_11460_1636# VPWR 0.23804f
C3705 _359_.B _371_.A3 0.00446f
C3706 _388_.B a_45148_30951# 0.00425f
C3707 a_44612_31048# a_44632_30206# 0.017f
C3708 _436_.B _260_.A2 0.00986f
C3709 a_48868_31048# _392_.A2 0.00246f
C3710 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _267_.ZN 0.00712f
C3711 a_68020_20452# VPWR 0.23672f
C3712 a_60380_1159# VPWR 0.29679f
C3713 a_64188_1159# a_64548_1256# 0.08717f
C3714 a_32380_1592# a_32828_1592# 0.01288f
C3715 a_36324_1636# a_36412_1592# 0.28563f
C3716 a_46628_11044# a_47076_11044# 0.01328f
C3717 a_36996_25156# a_36636_25112# 0.0869f
C3718 _350_.A1 _290_.ZN 0.08815f
C3719 a_1468_18407# VPWR 0.29679f
C3720 a_16700_29383# uio_oe[0] 0.0027f
C3721 a_4852_16936# a_5300_16936# 0.01328f
C3722 _371_.A2 a_26556_27815# 0.0013f
C3723 _311_.Z a_34715_22137# 0.00189f
C3724 _230_.I _238_.ZN 0.04335f
C3725 a_43044_27912# a_43492_27912# 0.01328f
C3726 _336_.A2 _336_.Z 0.50582f
C3727 a_48384_26724# _284_.A2 0.02165f
C3728 _330_.A1 _316_.A3 0.35385f
C3729 _452_.CLK a_45396_22020# 0.01003f
C3730 a_60828_1592# a_60828_1159# 0.05841f
C3731 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _390_.ZN 0.07465f
C3732 a_21764_2824# a_21628_1592# 0.00154f
C3733 a_23084_21976# VPWR 0.31436f
C3734 _455_.Q a_26468_27912# 0.00983f
C3735 _337_.A3 a_25796_27912# 0.06394f
C3736 a_33500_18840# a_33948_18840# 0.0131f
C3737 _447_.Q _317_.A2 0.97462f
C3738 a_51620_19911# a_52016_19759# 0.00232f
C3739 _439_.ZN VPWR 0.57915f
C3740 a_40444_2727# VPWR 0.31143f
C3741 _412_.A1 _384_.A3 0.90799f
C3742 a_61524_13800# VPWR 0.20622f
C3743 a_2364_26247# a_2724_26344# 0.08717f
C3744 a_16588_26247# a_17036_26247# 0.0131f
C3745 _337_.ZN _336_.A1 0.57733f
C3746 a_9308_29816# VPWR 0.3289f
C3747 _388_.B a_43232_29480# 0.03473f
C3748 a_1916_10567# VPWR 0.297f
C3749 a_62196_16936# a_62172_15704# 0.0016f
C3750 a_65332_16936# a_65220_15748# 0.02666f
C3751 uio_in[1] uio_in[2] 0.01021f
C3752 a_7628_30951# uio_oe[6] 0.00315f
C3753 _451_.Q a_40668_20408# 0.01696f
C3754 _359_.B uo_out[7] 0.07385f
C3755 a_27900_23111# VPWR 0.31431f
C3756 _439_.ZN a_41012_23208# 0.00183f
C3757 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I a_65756_23111# 0.01035f
C3758 _311_.A2 _452_.Q 0.03488f
C3759 _397_.A2 clk 0.07005f
C3760 _230_.I a_63721_28776# 0.00288f
C3761 _284_.ZN hold1.Z 0.00136f
C3762 a_56964_26724# VPWR 0.6314f
C3763 a_44252_2727# a_44612_2824# 0.08717f
C3764 _264_.B a_41488_24072# 0.02462f
C3765 _441_.A2 _301_.A1 0.00937f
C3766 a_66540_16839# a_66452_16936# 0.28563f
C3767 a_64412_18407# a_64860_18407# 0.0131f
C3768 a_20980_23588# a_20620_23544# 0.08707f
C3769 a_3260_25112# a_3708_25112# 0.0131f
C3770 a_1020_13703# a_932_13800# 0.28563f
C3771 _416_.A3 a_46252_19759# 0.00248f
C3772 _359_.B _480_.Q 0.03595f
C3773 a_25548_20408# a_26220_20408# 0.00544f
C3774 a_27476_20452# a_27924_20452# 0.01328f
C3775 _325_.ZN a_44724_17316# 0.00175f
C3776 a_41476_26344# _435_.A3 0.01196f
C3777 a_35232_24029# VPWR 0.51773f
C3778 a_62084_18504# a_62084_17316# 0.05841f
C3779 _246_.B2 _243_.A1 0.0011f
C3780 a_2364_16839# a_2276_16936# 0.28563f
C3781 _284_.ZN a_45396_25156# 0.00948f
C3782 a_65444_12612# a_65892_12612# 0.01328f
C3783 a_17596_1592# VPWR 0.29825f
C3784 a_62308_12612# a_61948_12568# 0.08707f
C3785 _304_.B a_40780_27815# 0.00582f
C3786 a_51332_24072# VPWR 1.32324f
C3787 _251_.A1 _243_.ZN 0.00461f
C3788 _384_.A3 a_51968_26724# 0.00296f
C3789 a_34756_24776# a_33376_23659# 0.00999f
C3790 a_36656_29123# uo_out[7] 0.00716f
C3791 a_65084_15271# a_65444_15368# 0.0869f
C3792 vgaringosc.workerclkbuff_notouch_.I _397_.A1 0.00107f
C3793 _363_.Z uo_out[4] 0.00501f
C3794 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN a_59172_23588# 0.03831f
C3795 a_11460_1636# a_11324_1159# 0.00168f
C3796 a_62420_12232# a_62396_11000# 0.0016f
C3797 _330_.ZN VPWR 0.4182f
C3798 _474_.CLK a_53704_23219# 0.01923f
C3799 _252_.ZN a_61412_27912# 0.00427f
C3800 _441_.A3 a_40656_23588# 0.00196f
C3801 a_22064_27912# VPWR 1.11159f
C3802 _459_.CLK uio_out[4] 0.07387f
C3803 a_3172_26724# a_3260_26680# 0.28563f
C3804 _443_.D a_37532_26247# 0.00227f
C3805 a_66228_10664# a_66676_10664# 0.01328f
C3806 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I a_55956_25940# 0.0021f
C3807 _267_.A2 _228_.ZN 0.0022f
C3808 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I 0.65437f
C3809 _433_.ZN _432_.ZN 0.21632f
C3810 a_35740_1159# a_36188_1159# 0.0131f
C3811 _400_.ZN a_46068_25156# 0.00338f
C3812 a_30795_29977# a_31080_29977# 0.00277f
C3813 _452_.CLK a_33860_20072# 0.00785f
C3814 a_32380_26247# a_32292_26344# 0.28563f
C3815 _371_.ZN a_28000_29480# 0.06669f
C3816 a_3172_20452# VPWR 0.20993f
C3817 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN a_64324_29860# 0.00591f
C3818 a_41922_31073# uo_out[3] 0.00223f
C3819 a_37291_29535# a_37536_29167# 0.00232f
C3820 _388_.B a_42820_31048# 0.01897f
C3821 a_62844_2727# VPWR 0.31143f
C3822 a_50660_12612# VPWR 0.22943f
C3823 a_65668_2824# a_65756_1159# 0.0027f
C3824 a_67436_18407# a_67796_18504# 0.08663f
C3825 _427_.A2 a_53660_21543# 0.00695f
C3826 clkload0.Z _381_.A2 0.00345f
C3827 a_39684_15368# a_40132_15368# 0.01328f
C3828 a_31620_20072# VPWR 0.20348f
C3829 _304_.ZN a_44028_22020# 0.00173f
C3830 a_3260_29383# a_3172_29480# 0.28563f
C3831 a_65196_23544# a_65644_23544# 0.01222f
C3832 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN a_67124_20452# 0.00189f
C3833 a_63404_10567# VPWR 0.31547f
C3834 a_3260_15704# a_3260_15271# 0.05841f
C3835 a_41564_15271# a_41476_15368# 0.28563f
C3836 _447_.Q _434_.ZN 0.06582f
C3837 _319_.A2 a_35492_20072# 0.01363f
C3838 a_35816_21192# a_36548_21640# 0.02091f
C3839 a_63964_17272# a_63988_16936# 0.00172f
C3840 a_25348_23208# VPWR 0.20728f
C3841 _238_.I a_59348_29076# 0.00197f
C3842 a_40244_18180# a_40452_18180# 0.00478f
C3843 a_60828_26680# a_60212_25156# 0.00235f
C3844 a_43132_15271# a_43580_15271# 0.0131f
C3845 a_52024_20083# a_52512_19715# 0.8399f
C3846 a_27588_26724# VPWR 0.21161f
C3847 a_33812_29860# uo_out[4] 0.00223f
C3848 a_14708_22020# a_15156_22020# 0.01328f
C3849 a_55676_2727# a_55588_2824# 0.28563f
C3850 a_60940_15704# VPWR 0.33181f
C3851 a_39324_19975# a_39684_20072# 0.0869f
C3852 a_67100_17272# a_67548_17272# 0.01222f
C3853 a_21316_23208# a_21404_21543# 0.00151f
C3854 _274_.A1 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.05533f
C3855 a_5188_1256# VPWR 0.20348f
C3856 a_5636_31048# VPWR 0.20815f
C3857 a_24788_23588# a_24428_23544# 0.08717f
C3858 a_27476_23588# a_27924_23588# 0.01328f
C3859 a_36548_1256# a_36996_1256# 0.01328f
C3860 a_19636_25156# a_19276_25112# 0.08707f
C3861 a_1380_4772# VPWR 0.20348f
C3862 a_51532_13703# a_51892_13800# 0.08707f
C3863 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I 0.68625f
C3864 a_57468_16839# a_58164_16936# 0.01227f
C3865 a_65420_13703# a_65868_13703# 0.0131f
C3866 a_35008_22461# VPWR 0.55267f
C3867 _281_.ZN a_52081_21236# 0.00192f
C3868 a_15580_2727# a_16252_2727# 0.00544f
C3869 a_33076_20452# a_33164_20408# 0.28563f
C3870 _370_.B a_32476_28776# 0.0012f
C3871 a_38316_16839# a_38676_16936# 0.08707f
C3872 a_55564_10567# a_55588_9476# 0.0016f
C3873 a_45284_10664# a_45284_9476# 0.05841f
C3874 a_63180_16839# VPWR 0.31594f
C3875 a_41564_1592# a_41700_1256# 0.00168f
C3876 a_31260_1592# VPWR 0.32824f
C3877 _447_.Q a_36772_23208# 0.01314f
C3878 a_40780_27815# VPWR 0.31508f
C3879 a_2724_1636# a_2364_1592# 0.08707f
C3880 a_61412_27912# a_61500_26247# 0.0027f
C3881 a_932_29860# a_1380_29860# 0.01328f
C3882 a_2724_17316# a_3172_17316# 0.01328f
C3883 a_54020_21640# VPWR 0.20911f
C3884 a_54356_23588# clk 0.00645f
C3885 a_56708_11044# a_56796_11000# 0.28563f
C3886 _304_.B _303_.ZN 1.22055f
C3887 a_51668_16936# a_52116_16936# 0.01328f
C3888 a_46044_1592# a_46492_1592# 0.01288f
C3889 _251_.A1 _258_.ZN 0.08143f
C3890 _265_.ZN a_41872_28409# 0.00207f
C3891 _284_.B _279_.Z 0.00997f
C3892 a_20756_26724# _455_.D 0.03559f
C3893 _294_.A2 _223_.I 1.31658f
C3894 clkbuf_1_0__f_clk.I _441_.A2 0.00188f
C3895 uio_in[5] uio_in[4] 0.01021f
C3896 a_50280_19369# VPWR 0.21462f
C3897 _247_.ZN a_60276_29032# 0.01366f
C3898 _451_.Q a_40780_21543# 0.02074f
C3899 a_22324_20452# VPWR 0.22767f
C3900 _336_.A1 a_27924_24776# 0.002f
C3901 a_36548_25156# _444_.D 0.01357f
C3902 a_1828_15748# a_1916_15704# 0.28563f
C3903 a_56796_12568# VPWR 0.3337f
C3904 a_16612_2824# a_17060_2824# 0.01328f
C3905 a_47724_18840# a_47748_17316# 0.00131f
C3906 a_48888_19243# a_49540_17316# 0.00107f
C3907 a_14236_29383# a_14596_29480# 0.08717f
C3908 a_25652_31048# a_25792_30301# 0.00585f
C3909 _379_.A2 a_19372_30345# 0.00317f
C3910 a_54108_21543# a_54020_21640# 0.28563f
C3911 a_2812_8999# a_2724_9096# 0.28563f
C3912 a_57492_10664# VPWR 0.2121f
C3913 a_58252_18407# a_58164_18504# 0.28563f
C3914 _378_.ZN a_17932_27815# 0.0245f
C3915 a_52540_15271# a_52900_15368# 0.08717f
C3916 a_56124_27815# a_56036_27912# 0.28563f
C3917 a_55676_27815# vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.00718f
C3918 _304_.B _397_.A4 0.80434f
C3919 a_3708_7431# a_3620_7528# 0.28563f
C3920 a_43126_24119# a_43750_23544# 0.10659f
C3921 a_4940_5863# a_4852_5960# 0.28563f
C3922 a_64412_4295# a_64324_4392# 0.28563f
C3923 _495_.I a_43268_31048# 0.00189f
C3924 a_4068_21640# a_4068_20452# 0.05841f
C3925 a_30724_15368# VPWR 0.22176f
C3926 a_66652_2727# a_67012_2824# 0.0869f
C3927 a_21876_22020# a_21516_21976# 0.08663f
C3928 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN 0.21302f
C3929 a_33948_15271# VPWR 0.33071f
C3930 a_2724_14180# a_3172_14180# 0.01328f
C3931 a_60828_26680# VPWR 0.35008f
C3932 _275_.A2 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I 0.49226f
C3933 a_66564_17316# VPWR 0.20904f
C3934 a_31920_29480# VPWR 1.10462f
C3935 _251_.A1 a_62560_25112# 0.77089f
C3936 a_50996_28292# _408_.ZN 0.00615f
C3937 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I 0.00393f
C3938 a_27588_1256# VPWR 0.2304f
C3939 a_3708_7431# VPWR 0.33374f
C3940 _474_.CLK _428_.Z 0.00286f
C3941 a_30836_23588# a_30476_23544# 0.0869f
C3942 a_25936_25597# a_25643_25273# 0.49319f
C3943 a_64412_4295# VPWR 0.3038f
C3944 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I 0.00586f
C3945 a_62508_13703# a_62420_13800# 0.28563f
C3946 _260_.A1 _433_.ZN 0.42328f
C3947 _261_.ZN _432_.ZN 0.00918f
C3948 vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN a_54804_18504# 0.00359f
C3949 a_10092_30951# VPWR 0.31381f
C3950 a_31260_17272# a_31260_16839# 0.05841f
C3951 a_35204_17316# a_35180_16839# 0.00172f
C3952 a_28124_30600# uio_out[0] 0.09659f
C3953 a_49292_16839# a_49204_16936# 0.28563f
C3954 a_1380_23208# a_1380_22020# 0.05841f
C3955 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_55228_27815# 0.01967f
C3956 a_23868_26247# a_23780_26344# 0.28563f
C3957 a_42932_16936# VPWR 0.21984f
C3958 a_45060_1636# VPWR 0.20348f
C3959 a_7964_1159# a_8548_1256# 0.01675f
C3960 a_1380_29480# a_1828_29480# 0.01328f
C3961 a_9220_1636# a_9668_1636# 0.01328f
C3962 uo_out[4] uo_out[3] 0.03336f
C3963 a_52428_12135# a_52876_12135# 0.01288f
C3964 a_66428_12568# a_66316_12135# 0.02634f
C3965 uo_out[2] uo_out[1] 0.08493f
C3966 a_23532_23544# a_23644_23111# 0.02634f
C3967 _452_.CLK a_36548_26724# 0.05188f
C3968 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I 0.00292f
C3969 _325_.B a_43664_17317# 0.01027f
C3970 a_8100_29860# a_7740_29816# 0.08663f
C3971 a_41440_28363# a_41996_28777# 0.8399f
C3972 _265_.ZN a_42368_28733# 0.01755f
C3973 _416_.ZN a_45820_18840# 0.00952f
C3974 _303_.ZN VPWR 1.71865f
C3975 a_50300_11000# a_50188_10567# 0.02634f
C3976 _398_.C a_53704_23219# 0.00194f
C3977 a_7428_2824# VPWR 0.20815f
C3978 a_53348_1636# a_52988_1592# 0.08707f
C3979 _249_.A2 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I 0.69155f
C3980 _243_.ZN a_58020_27508# 0.44493f
C3981 _252_.ZN _251_.ZN 0.27514f
C3982 a_14796_24679# a_15244_24679# 0.0131f
C3983 a_53100_18407# a_53012_18504# 0.28563f
C3984 a_58140_1159# a_58588_1159# 0.0131f
C3985 a_66228_20452# a_66316_20408# 0.28563f
C3986 a_66676_20452# a_67124_20452# 0.01328f
C3987 a_61188_15368# VPWR 0.23106f
C3988 _304_.B a_51956_26183# 0.01032f
C3989 a_66652_18840# a_67100_18840# 0.01255f
C3990 a_53460_18504# VPWR 0.20595f
C3991 a_17484_25112# VPWR 0.29719f
C3992 _461_.D a_32916_29860# 0.00621f
C3993 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I a_63964_19975# 0.00286f
C3994 _324_.B a_45156_21236# 0.00439f
C3995 a_27004_30951# VPWR 0.37312f
C3996 a_16028_29816# a_16052_28292# 0.00134f
C3997 _421_.B _473_.Q 0.00551f
C3998 a_33164_20408# VPWR 0.34815f
C3999 a_31620_15748# a_31708_15704# 0.28563f
C4000 a_35204_15748# a_35652_15748# 0.01328f
C4001 a_3708_12135# VPWR 0.33374f
C4002 _393_.A1 a_45484_28248# 0.00508f
C4003 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN a_67772_21543# 0.00306f
C4004 _397_.A1 a_48292_26369# 0.00116f
C4005 _325_.A1 _452_.D 0.00138f
C4006 vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN 0.00999f
C4007 a_51332_24072# a_51240_23340# 0.00205f
C4008 _379_.A2 a_20003_29611# 0.03277f
C4009 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN VPWR 0.76452f
C4010 _424_.B1 _281_.ZN 0.59502f
C4011 _397_.A4 VPWR 1.35334f
C4012 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN VPWR 1.36116f
C4013 _268_.A2 _251_.A1 0.09456f
C4014 _452_.CLK a_40108_16839# 0.00239f
C4015 a_28796_21543# a_28820_20452# 0.0016f
C4016 a_1468_15704# VPWR 0.29679f
C4017 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN 0.03839f
C4018 a_52900_15368# VPWR 0.21513f
C4019 a_24788_22020# a_24876_21976# 0.28563f
C4020 a_28372_22020# a_28820_22020# 0.01328f
C4021 a_56348_15271# VPWR 0.31569f
C4022 a_46604_16839# a_47052_16839# 0.01288f
C4023 a_37868_16839# VPWR 0.31389f
C4024 _395_.A1 a_49764_26724# 0.0296f
C4025 a_49764_1256# VPWR 0.21599f
C4026 a_58948_1256# a_59396_1256# 0.01328f
C4027 a_26108_30951# a_26020_31048# 0.28563f
C4028 a_59284_13800# a_59732_13800# 0.01328f
C4029 a_37980_2727# a_38428_2727# 0.0131f
C4030 a_56516_26344# a_56388_25940# 0.00284f
C4031 _359_.ZN a_32592_25227# 0.0034f
C4032 a_19076_23208# a_19188_22020# 0.02666f
C4033 _231_.ZN a_59172_23588# 0.13441f
C4034 a_36100_17316# VPWR 0.20639f
C4035 a_19388_1159# a_19300_1256# 0.28563f
C4036 a_51196_1592# VPWR 0.3289f
C4037 a_49740_12135# a_49652_12232# 0.28563f
C4038 a_63292_12568# a_63316_12232# 0.00172f
C4039 a_15940_1636# a_16612_1636# 0.00347f
C4040 a_22636_25112# a_22660_24776# 0.00172f
C4041 a_39268_18840# a_40416_18885# 0.00291f
C4042 _421_.B _475_.D 0.08581f
C4043 a_14596_29860# a_15044_29860# 0.01328f
C4044 a_11012_29860# a_11100_29816# 0.28563f
C4045 _474_.CLK _470_.Q 0.30493f
C4046 a_37084_17272# a_37532_17272# 0.01288f
C4047 a_57244_11000# a_57132_10567# 0.02634f
C4048 a_66876_11000# a_67324_11000# 0.01288f
C4049 _390_.ZN _392_.A2 0.08497f
C4050 a_29828_2824# VPWR 0.20348f
C4051 a_56260_1636# a_56348_1592# 0.28563f
C4052 a_59844_1636# a_60292_1636# 0.01328f
C4053 _384_.A3 _473_.Q 0.41908f
C4054 a_43788_29167# VPWR 0.39596f
C4055 a_4156_23111# a_4852_23208# 0.01227f
C4056 _300_.A2 a_38764_20408# 0.07671f
C4057 _416_.A3 a_47860_21640# 0.01723f
C4058 a_25436_23111# a_25884_23111# 0.012f
C4059 a_17036_24679# a_17396_24776# 0.08717f
C4060 a_1828_9476# VPWR 0.20348f
C4061 _340_.A2 _359_.B 0.03135f
C4062 a_50660_14180# VPWR 0.2267f
C4063 a_9444_2824# a_9532_1159# 0.0027f
C4064 a_4940_18407# a_4852_18504# 0.28563f
C4065 a_51956_26183# VPWR 0.36905f
C4066 a_37084_26680# a_37084_26247# 0.05841f
C4067 a_26468_31048# a_26720_30301# 0.0031f
C4068 a_2276_31048# a_2276_29860# 0.05841f
C4069 a_65420_12135# VPWR 0.32173f
C4070 a_14596_29480# VPWR 0.20665f
C4071 a_26556_2727# a_26692_1636# 0.00154f
C4072 a_39012_2824# a_39460_2824# 0.01328f
C4073 _416_.A1 a_45128_26031# 0.00913f
C4074 a_43750_23544# a_44282_24164# 0.0013f
C4075 _459_.Q _359_.B 0.10193f
C4076 _261_.ZN _260_.A1 0.06424f
C4077 a_1380_24776# VPWR 0.20348f
C4078 _476_.Q _427_.ZN 0.02442f
C4079 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I VPWR 0.84781f
C4080 a_66116_7528# VPWR 0.23643f
C4081 a_932_3204# VPWR 0.22176f
C4082 a_27364_21640# a_27476_20452# 0.02666f
C4083 a_40356_15748# VPWR 0.20671f
C4084 a_1020_19975# a_1380_20072# 0.08717f
C4085 _324_.C vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.00427f
C4086 a_52024_20083# a_53348_18884# 0.00179f
C4087 a_56236_23544# a_56124_23111# 0.02634f
C4088 a_30836_22020# a_30476_21976# 0.0869f
C4089 a_45732_9476# a_46180_9476# 0.01328f
C4090 _285_.Z a_39480_28776# 0.00891f
C4091 a_49496_30345# _392_.A2 0.01005f
C4092 a_51644_14136# a_52092_14136# 0.01288f
C4093 a_44864_27165# VPWR 0.50827f
C4094 _265_.ZN a_43132_27815# 0.0052f
C4095 _459_.CLK a_24228_26344# 0.01229f
C4096 a_26427_29977# a_26712_29977# 0.00277f
C4097 _294_.A2 a_37584_29123# 0.00648f
C4098 _398_.C _428_.Z 0.14479f
C4099 _397_.A4 a_50068_27508# 0.04011f
C4100 _300_.ZN a_40656_23588# 0.01541f
C4101 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN a_55140_15748# 0.00471f
C4102 a_35710_28776# uo_out[7] 0.00171f
C4103 a_50412_18407# a_50436_17316# 0.0016f
C4104 a_48196_17316# VPWR 0.20897f
C4105 _454_.Q _455_.Q 0.16831f
C4106 a_64996_1636# VPWR 0.20816f
C4107 a_67124_10664# a_67100_9432# 0.0016f
C4108 a_30364_1159# a_30724_1256# 0.08717f
C4109 a_46180_12232# a_46628_12232# 0.01328f
C4110 a_60268_12135# a_60628_12232# 0.08707f
C4111 a_57692_12568# a_57604_11044# 0.00151f
C4112 a_57044_23588# a_57020_23111# 0.00172f
C4113 a_31820_23544# a_31844_23208# 0.00172f
C4114 a_19300_1636# a_19388_1592# 0.28563f
C4115 a_22884_1636# a_23332_1636# 0.01328f
C4116 _359_.B _461_.D 0.6237f
C4117 a_17060_29860# a_17148_29816# 0.28563f
C4118 _365_.ZN _460_.Q 0.0205f
C4119 a_44340_26183# _284_.B 0.00619f
C4120 _381_.A2 a_50120_26476# 0.0375f
C4121 a_20956_21543# VPWR 0.31389f
C4122 _397_.A2 a_49652_29480# 0.02474f
C4123 _416_.A1 _267_.ZN 0.00121f
C4124 _279_.Z _474_.Q 0.63344f
C4125 _260_.A2 _433_.ZN 0.05849f
C4126 a_54108_11000# a_54132_10664# 0.00172f
C4127 a_39548_1592# a_39548_1159# 0.05841f
C4128 a_64188_11000# a_64300_10567# 0.02634f
C4129 a_52228_2824# VPWR 0.20815f
C4130 a_52756_29076# VPWR 0.58765f
C4131 a_24540_23111# a_24452_23208# 0.28563f
C4132 a_19524_24776# a_19972_24776# 0.01328f
C4133 a_56124_28248# _241_.I0 0.02344f
C4134 a_51420_9432# VPWR 0.31143f
C4135 _416_.A1 _390_.ZN 0.9319f
C4136 a_60740_2824# a_60740_1636# 0.05841f
C4137 a_56932_2824# a_56796_1592# 0.00154f
C4138 a_57692_14136# VPWR 0.33325f
C4139 a_35092_18504# a_35540_18504# 0.01328f
C4140 a_45284_15748# a_45372_15704# 0.28563f
C4141 a_59284_12232# VPWR 0.20595f
C4142 a_41340_15704# a_41788_15704# 0.01288f
C4143 _342_.ZN _343_.A2 0.21315f
C4144 _452_.CLK a_45696_20072# 0.01964f
C4145 a_62532_30736# vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN 0.00486f
C4146 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I clk 0.03622f
C4147 a_34396_24679# VPWR 0.33297f
C4148 a_52848_25987# _412_.ZN 0.23238f
C4149 _245_.I1 vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN 0.00474f
C4150 a_64772_20072# VPWR 0.20727f
C4151 _459_.Q a_32144_26724# 0.00122f
C4152 a_10428_2727# a_10788_2824# 0.08717f
C4153 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN a_63316_20452# 0.05209f
C4154 _397_.A1 a_49764_26724# 0.00136f
C4155 _441_.A3 _448_.Q 0.0158f
C4156 a_62620_19975# a_63068_19975# 0.0131f
C4157 a_46492_15704# VPWR 0.30141f
C4158 a_57156_27912# a_56964_26724# 0.00181f
C4159 a_51332_9476# a_51420_9432# 0.28563f
C4160 a_26556_30951# uio_out[2] 0.00333f
C4161 a_60180_14180# a_59820_14136# 0.0869f
C4162 a_932_20452# a_1380_20452# 0.01328f
C4163 a_61860_30736# VPWR 0.55097f
C4164 _324_.C a_45169_27509# 0.0013f
C4165 _419_.A4 a_48384_26724# 0.00232f
C4166 a_60380_2727# a_60828_2727# 0.0131f
C4167 a_48420_12612# a_48868_12612# 0.01328f
C4168 _381_.Z a_49952_26724# 0.00236f
C4169 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN 0.06536f
C4170 a_15132_1159# VPWR 0.29679f
C4171 a_41788_1159# a_41700_1256# 0.28563f
C4172 a_31844_23208# a_31820_21976# 0.0016f
C4173 a_65756_18840# a_65668_17316# 0.0027f
C4174 a_61052_12568# a_60964_11044# 0.00151f
C4175 a_932_6340# a_1020_6296# 0.28563f
C4176 a_4068_20072# a_4852_20072# 0.00276f
C4177 a_3620_12232# a_3620_11044# 0.05841f
C4178 a_64772_5960# a_64772_4772# 0.05841f
C4179 a_65668_4392# a_65668_3204# 0.05841f
C4180 _474_.CLK a_52744_26031# 0.003f
C4181 a_60285_30600# _255_.I 0.0029f
C4182 _237_.A1 _324_.C 0.56008f
C4183 a_17844_21640# VPWR 0.21215f
C4184 a_49180_17272# a_49628_17272# 0.01288f
C4185 a_54824_22045# a_55744_22505# 0.00306f
C4186 a_53124_17316# a_53212_17272# 0.28563f
C4187 a_22059_26399# a_22548_25156# 0.03071f
C4188 _470_.Q _398_.C 0.00183f
C4189 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_59372_13703# 0.00283f
C4190 _355_.C _340_.ZN 0.17836f
C4191 a_47164_10567# a_47524_10664# 0.08717f
C4192 a_1916_1159# a_2364_1159# 0.0131f
C4193 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I VPWR 0.88326f
C4194 a_61164_10567# a_61612_10567# 0.01288f
C4195 a_7428_2824# a_7292_1592# 0.00154f
C4196 _370_.B a_31920_29480# 0.06575f
C4197 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN 0.00361f
C4198 a_53648_23263# VPWR 0.00204f
C4199 a_23108_23208# a_23556_23208# 0.01328f
C4200 a_65108_23588# clk 0.00647f
C4201 a_62396_9432# VPWR 0.31143f
C4202 a_15604_23588# VPWR 0.20348f
C4203 a_65220_6340# VPWR 0.20921f
C4204 a_45372_13703# VPWR 0.30073f
C4205 a_17484_21543# a_17396_21640# 0.28563f
C4206 a_29692_21543# a_30140_21543# 0.01288f
C4207 a_67012_3204# VPWR 0.20348f
C4208 a_65668_2824# a_65532_1592# 0.00154f
C4209 a_31844_2824# a_31932_1159# 0.0027f
C4210 a_45036_28248# _330_.A1 0.03157f
C4211 _384_.A3 a_51540_24776# 0.00228f
C4212 a_18180_31048# a_18044_29816# 0.00154f
C4213 _427_.ZN a_55364_21640# 0.00684f
C4214 a_25232_27165# a_24860_27209# 0.10745f
C4215 a_36188_25112# VPWR 0.32608f
C4216 a_48420_11044# VPWR 0.20348f
C4217 clkbuf_1_0__f_clk.I a_46356_24072# 0.03126f
C4218 a_48644_15748# a_48284_15704# 0.08707f
C4219 a_61188_2824# a_61860_2824# 0.00347f
C4220 _455_.Q a_23284_26724# 0.00204f
C4221 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I _248_.B1 0.00144f
C4222 a_35504_18955# VPWR 1.10973f
C4223 a_18716_26247# VPWR 0.32987f
C4224 a_21852_2727# a_21764_2824# 0.28563f
C4225 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I 0.10617f
C4226 a_56708_9476# a_57156_9476# 0.01328f
C4227 a_2724_1256# a_3172_1256# 0.01328f
C4228 a_3172_31048# a_3620_31048# 0.01328f
C4229 a_64100_14180# a_63740_14136# 0.08707f
C4230 _261_.ZN _260_.A2 0.15945f
C4231 a_67236_14180# a_67684_14180# 0.01328f
C4232 a_14708_20452# a_14796_20408# 0.28563f
C4233 _279_.Z a_46984_23588# 0.0241f
C4234 a_20284_1592# a_20420_1256# 0.00168f
C4235 _242_.Z vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I 0.05929f
C4236 a_64212_13800# a_64188_12568# 0.0016f
C4237 a_50548_13800# a_50636_12135# 0.00151f
C4238 _241_.I0 a_56836_27208# 0.01094f
C4239 _337_.ZN a_27676_26247# 0.00149f
C4240 _300_.ZN a_39475_21236# 0.00467f
C4241 _284_.ZN a_43003_28409# 0.03277f
C4242 a_27172_24328# a_27028_23588# 0.03517f
C4243 _252_.ZN a_60604_27815# 0.04048f
C4244 a_37532_1159# VPWR 0.3289f
C4245 a_51892_12232# a_52004_11044# 0.02666f
C4246 a_52764_1159# a_53124_1256# 0.08717f
C4247 a_29020_1592# a_29468_1592# 0.01288f
C4248 _260_.A1 _327_.Z 0.00685f
C4249 a_45920_20523# a_46848_20893# 1.16391f
C4250 a_35232_24029# _311_.Z 0.0011f
C4251 a_34939_23705# a_34980_22895# 0.02615f
C4252 _419_.A4 a_47259_20127# 0.0026f
C4253 a_58476_10567# a_58388_10664# 0.28563f
C4254 a_64324_29860# VPWR 0.14875f
C4255 a_932_18504# a_932_17316# 0.05841f
C4256 _381_.A2 a_50308_26476# 0.00216f
C4257 _459_.CLK a_35728_29480# 0.04746f
C4258 _330_.ZN a_38676_16936# 0.00388f
C4259 a_54892_19975# VPWR 0.31556f
C4260 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN a_61164_23111# 0.00471f
C4261 a_16500_22020# VPWR 0.20348f
C4262 _393_.A3 _470_.Q 0.022f
C4263 _417_.A2 a_50644_21640# 0.00168f
C4264 a_23084_23544# VPWR 0.31389f
C4265 a_67212_13703# VPWR 0.31431f
C4266 a_17596_2727# VPWR 0.31289f
C4267 a_1468_18840# a_1916_18840# 0.0131f
C4268 a_4068_18884# a_3708_18840# 0.08717f
C4269 a_28348_21543# a_28708_21640# 0.08707f
C4270 _411_.A2 _284_.A2 1.12853f
C4271 a_2724_29860# VPWR 0.20782f
C4272 a_45416_29885# VPWR 1.1029f
C4273 _287_.A1 a_32476_29167# 0.02295f
C4274 a_53212_29816# _267_.A2 0.51515f
C4275 a_55140_15748# vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I 0.00242f
C4276 a_54556_11000# VPWR 0.31436f
C4277 a_20396_26680# VPWR 0.31993f
C4278 _294_.ZN uo_out[4] 1.89789f
C4279 _452_.Q a_38764_20408# 0.00167f
C4280 a_22992_27555# a_23627_27967# 0.02112f
C4281 a_66564_15748# a_66652_15704# 0.28563f
C4282 a_16140_27815# VPWR 0.29679f
C4283 a_32828_2727# a_33188_2824# 0.08717f
C4284 a_63316_23588# a_63764_23588# 0.01328f
C4285 _276_.A2 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN 0.00127f
C4286 _342_.ZN a_24952_29032# 0.02541f
C4287 _330_.A1 _448_.Q 0.01713f
C4288 a_62308_9476# a_62396_9432# 0.28563f
C4289 a_61500_27815# _245_.Z 0.00277f
C4290 a_28124_26680# _355_.B 0.00993f
C4291 a_21652_20452# a_22324_20452# 0.00347f
C4292 a_19948_20408# a_20396_20408# 0.0131f
C4293 _437_.A1 _435_.ZN 0.11842f
C4294 _275_.A2 _416_.A1 0.47377f
C4295 _324_.C a_43444_19668# 0.00379f
C4296 a_58924_18840# a_58836_17316# 0.00251f
C4297 a_5276_30951# a_5636_31048# 0.0869f
C4298 a_25796_27912# a_24304_26795# 0.00103f
C4299 a_11012_1636# VPWR 0.21526f
C4300 _459_.CLK a_21516_25112# 0.00593f
C4301 a_54556_12568# a_55004_12568# 0.01288f
C4302 a_58500_12612# a_58588_12568# 0.28563f
C4303 vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I 0.06742f
C4304 a_37516_27599# a_37444_26724# 0.00175f
C4305 _388_.B a_44700_30951# 0.01415f
C4306 _474_.CLK a_56932_23208# 0.00279f
C4307 a_35540_18504# a_35628_16839# 0.00151f
C4308 a_25796_24776# a_25772_23544# 0.0016f
C4309 a_9756_29816# a_9892_29480# 0.00168f
C4310 _369_.ZN _355_.B 0.00238f
C4311 _375_.Z a_22188_29383# 0.00135f
C4312 a_59932_1159# VPWR 0.29679f
C4313 a_58836_12232# a_58948_11044# 0.02666f
C4314 a_64188_1159# a_64100_1256# 0.28563f
C4315 _402_.A1 a_47636_25940# 0.00696f
C4316 a_67212_20408# VPWR 0.34932f
C4317 a_55028_12232# a_55004_11000# 0.0016f
C4318 a_36324_1636# a_35964_1592# 0.08707f
C4319 a_36548_25156# a_36636_25112# 0.28563f
C4320 a_1020_18407# VPWR 0.30073f
C4321 _416_.A3 a_47483_20569# 0.02887f
C4322 _311_.Z a_35008_22461# 0.00817f
C4323 _251_.A1 _241_.I0 1.33355f
C4324 a_41140_27912# _330_.A1 0.00866f
C4325 _452_.CLK a_44948_22020# 0.00134f
C4326 a_55028_10664# a_55476_10664# 0.01328f
C4327 a_24316_1159# a_24764_1159# 0.0131f
C4328 a_34644_18504# a_34756_17316# 0.02666f
C4329 _419_.A4 _419_.Z 0.61291f
C4330 a_22636_21976# VPWR 0.31898f
C4331 a_37644_23544# VPWR 0.35878f
C4332 a_61076_13800# VPWR 0.20622f
C4333 a_26916_21640# a_27364_21640# 0.01328f
C4334 _447_.Q a_36148_21976# 0.00374f
C4335 a_39996_2727# VPWR 0.31143f
C4336 _412_.A1 a_52900_26724# 0.00235f
C4337 a_2364_26247# a_2276_26344# 0.28563f
C4338 a_3172_15368# a_3620_15368# 0.01328f
C4339 a_8860_29816# VPWR 0.33352f
C4340 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN 0.01395f
C4341 _250_.C a_60940_28248# 0.00362f
C4342 a_1468_10567# VPWR 0.29679f
C4343 _324_.C _451_.Q 0.0202f
C4344 a_7180_30951# uio_oe[6] 0.00214f
C4345 a_5388_15271# a_5300_15368# 0.28563f
C4346 a_27452_23111# VPWR 0.3229f
C4347 _451_.Q a_40220_20408# 0.04206f
C4348 a_65644_23544# a_65756_23111# 0.02634f
C4349 a_31708_15271# a_32156_15271# 0.0131f
C4350 a_34939_23705# a_35224_23705# 0.00277f
C4351 _230_.I a_63313_28776# 0.00182f
C4352 a_60740_26724# a_61748_26724# 0.00196f
C4353 a_44252_2727# a_44164_2824# 0.28563f
C4354 _285_.Z _284_.ZN 0.29464f
C4355 a_64324_17316# a_64772_17316# 0.01328f
C4356 a_66092_16839# a_66452_16936# 0.0869f
C4357 _452_.CLK _260_.A1 0.00697f
C4358 a_16588_23544# a_17036_23544# 0.01288f
C4359 a_20532_23588# a_20620_23544# 0.28563f
C4360 a_25124_1256# a_25572_1256# 0.01328f
C4361 a_2364_5863# a_2812_5863# 0.0131f
C4362 a_65756_6296# a_65756_5863# 0.05841f
C4363 a_64860_7864# a_64860_7431# 0.05841f
C4364 a_1468_7431# a_1916_7431# 0.0131f
C4365 a_66652_4728# a_66652_4295# 0.05841f
C4366 a_3260_4295# a_3708_4295# 0.0131f
C4367 a_54220_13703# a_54668_13703# 0.01288f
C4368 _416_.A3 a_46624_19715# 0.04652f
C4369 _325_.ZN a_44276_17316# 0.01587f
C4370 a_4156_2727# a_4828_2727# 0.00544f
C4371 a_36436_16936# a_36412_15271# 0.00134f
C4372 _268_.A2 _409_.ZN 0.02601f
C4373 a_41028_26344# _435_.A3 0.02259f
C4374 _359_.B a_43232_29480# 0.04829f
C4375 _355_.C _355_.B 0.19443f
C4376 a_15580_29383# a_16252_29383# 0.00544f
C4377 a_33932_24073# VPWR 0.40749f
C4378 _402_.A1 a_46156_25112# 0.0133f
C4379 a_1916_16839# a_2276_16936# 0.08717f
C4380 a_17148_1592# VPWR 0.29679f
C4381 a_61860_12612# a_61948_12568# 0.28563f
C4382 _448_.Q _226_.ZN 0.02791f
C4383 a_52092_12568# a_51980_12135# 0.02634f
C4384 _284_.ZN a_44948_25156# 0.02777f
C4385 a_7180_30951# a_7628_30951# 0.01222f
C4386 _325_.B a_42996_18840# 0.04427f
C4387 a_20664_29977# uio_out[6] 0.00118f
C4388 a_35728_29480# uo_out[7] 0.0124f
C4389 a_65084_15271# a_64996_15368# 0.28563f
C4390 a_49404_11000# a_49852_11000# 0.01288f
C4391 a_40468_16936# a_40916_16936# 0.01328f
C4392 a_65780_12232# a_65892_11044# 0.02666f
C4393 a_42820_1636# a_43268_1636# 0.01328f
C4394 a_37408_18504# VPWR 1.10974f
C4395 _252_.ZN a_60964_27912# 0.01229f
C4396 _441_.A3 a_40452_23588# 0.02154f
C4397 a_21268_27912# VPWR 0.00405f
C4398 a_66652_15704# a_66788_15368# 0.00168f
C4399 a_3172_26724# a_2812_26680# 0.08717f
C4400 a_23556_29860# uio_out[4] 0.00308f
C4401 _474_.CLK _393_.ZN 0.00673f
C4402 _397_.A1 a_52676_27912# 0.00132f
C4403 _324_.C _384_.A3 0.07258f
C4404 a_16240_26795# a_17932_26247# 0.01084f
C4405 _448_.Q _300_.ZN 0.44148f
C4406 a_2724_20452# VPWR 0.20782f
C4407 a_31932_26247# a_32292_26344# 0.08674f
C4408 a_62396_2727# VPWR 0.31143f
C4409 a_50212_12612# VPWR 0.22223f
C4410 _388_.B a_41922_31073# 0.01658f
C4411 a_16948_26344# a_17396_26344# 0.01328f
C4412 a_48384_26724# _381_.A2 0.02124f
C4413 a_5052_28248# a_4964_26724# 0.00151f
C4414 a_5276_2727# a_5412_1636# 0.00154f
C4415 a_5188_2824# a_5636_2824# 0.01328f
C4416 a_67436_18407# a_67348_18504# 0.28563f
C4417 a_58028_17272# a_58476_17272# 0.01222f
C4418 a_2812_29383# a_3172_29480# 0.08717f
C4419 _351_.A2 a_25204_26841# 0.00135f
C4420 a_31172_20072# VPWR 0.20348f
C4421 _437_.A1 _441_.ZN 0.21925f
C4422 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN a_66676_20452# 0.0013f
C4423 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I 0.03176f
C4424 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.74677f
C4425 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN a_57132_18407# 0.00102f
C4426 a_62956_10567# VPWR 0.31547f
C4427 _459_.CLK _459_.D 0.03277f
C4428 a_41116_15271# a_41476_15368# 0.08717f
C4429 a_24900_23208# VPWR 0.20622f
C4430 a_51620_19911# a_52408_19759# 0.02112f
C4431 a_27140_26724# VPWR 0.17561f
C4432 a_4604_28248# a_5052_28248# 0.01222f
C4433 a_55228_2727# a_55588_2824# 0.08717f
C4434 _495_.I a_43232_29480# 0.00179f
C4435 a_39324_19975# a_39236_20072# 0.28563f
C4436 a_59172_23588# clk 0.00549f
C4437 _359_.B a_42820_31048# 0.0016f
C4438 a_21068_23544# a_20980_22020# 0.00151f
C4439 a_32516_16936# a_32516_15748# 0.05841f
C4440 a_51220_18504# a_51668_18504# 0.01328f
C4441 a_19188_25156# a_19276_25112# 0.28563f
C4442 a_4740_1256# VPWR 0.22423f
C4443 a_5188_31048# VPWR 0.20815f
C4444 a_24340_23588# a_24428_23544# 0.28563f
C4445 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I _250_.ZN 0.02715f
C4446 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN a_61412_17316# 0.00636f
C4447 a_15244_25112# a_15692_25112# 0.01288f
C4448 a_57468_16839# a_57380_16936# 0.28563f
C4449 _476_.Q a_51240_20452# 0.08134f
C4450 _256_.A2 ui_in[3] 0.00238f
C4451 _281_.ZN a_51877_21236# 0.00435f
C4452 a_30924_20408# a_31372_20408# 0.0131f
C4453 a_33076_20452# a_32716_20408# 0.08717f
C4454 a_33708_22505# VPWR 0.40534f
C4455 a_51532_13703# a_51444_13800# 0.28563f
C4456 a_24652_30951# a_25100_30951# 0.01222f
C4457 a_41228_27815# a_41392_27165# 0.00105f
C4458 _317_.A2 _319_.A2 0.85546f
C4459 a_61860_27912# _245_.Z 0.00165f
C4460 a_39268_18840# _331_.ZN 0.00882f
C4461 a_38316_16839# a_38228_16936# 0.28563f
C4462 a_31484_26680# _358_.A3 0.00707f
C4463 _281_.ZN a_46794_25156# 0.01244f
C4464 _474_.CLK _476_.Q 0.00235f
C4465 a_1468_12135# a_1916_12135# 0.0131f
C4466 a_59036_12568# a_58924_12135# 0.02634f
C4467 a_30812_1592# VPWR 0.29679f
C4468 a_62732_16839# VPWR 0.31594f
C4469 a_19636_23588# a_19612_23111# 0.00172f
C4470 a_2276_1636# a_2364_1592# 0.28563f
C4471 a_5860_1636# a_6308_1636# 0.01328f
C4472 a_15692_23544# a_15692_23111# 0.05841f
C4473 _294_.A2 _363_.Z 0.18943f
C4474 a_53572_21640# VPWR 0.1475f
C4475 a_34404_31048# uo_out[4] 0.00185f
C4476 a_41116_26247# _260_.A1 0.00127f
C4477 a_56708_11044# a_56348_11000# 0.08707f
C4478 a_59284_12232# a_59372_10567# 0.00151f
C4479 a_3260_11000# a_3260_10567# 0.05841f
C4480 _255_.I _243_.ZN 0.04607f
C4481 _251_.A1 a_56572_29383# 0.00383f
C4482 _350_.A1 _369_.ZN 0.04829f
C4483 _324_.B a_49604_22020# 0.00141f
C4484 _284_.B a_47297_25596# 0.01674f
C4485 _294_.A2 a_31396_31048# 0.02102f
C4486 a_20308_26724# _455_.D 0.00608f
C4487 a_20756_26724# a_20844_26680# 0.28563f
C4488 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I a_60416_25156# 0.00131f
C4489 a_46716_1159# a_47164_1159# 0.0131f
C4490 a_39460_2824# a_39460_1636# 0.05841f
C4491 a_35652_2824# a_35516_1592# 0.00154f
C4492 _294_.A2 a_36960_27912# 0.00117f
C4493 a_17932_27815# a_18096_27165# 0.00105f
C4494 a_64324_18884# a_64772_18884# 0.01328f
C4495 a_50384_19204# VPWR 0.42821f
C4496 a_21740_20408# VPWR 0.33981f
C4497 _336_.A2 a_26548_24372# 0.07315f
C4498 _451_.Q a_40332_21543# 0.04664f
C4499 _397_.A2 a_49044_28292# 0.00106f
C4500 a_36100_25156# _444_.D 0.02427f
C4501 _355_.C a_25643_25273# 0.01312f
C4502 a_56348_12568# VPWR 0.31423f
C4503 a_3620_15748# a_4068_15748# 0.01328f
C4504 a_1828_15748# a_1468_15704# 0.08717f
C4505 a_50660_15368# a_51108_15368# 0.01328f
C4506 a_14236_29383# a_14148_29480# 0.28563f
C4507 _252_.B a_59036_26247# 0.00195f
C4508 a_53660_21543# a_54020_21640# 0.0869f
C4509 _379_.A2 a_19744_30301# 0.00202f
C4510 a_19328_28733# a_20396_27815# 0.03096f
C4511 a_57044_10664# VPWR 0.23085f
C4512 a_57580_18407# a_58164_18504# 0.01675f
C4513 _419_.A4 _416_.A2 0.43889f
C4514 a_2364_8999# a_2724_9096# 0.08717f
C4515 a_55676_27815# a_56036_27912# 0.08663f
C4516 a_3260_7431# a_3620_7528# 0.08717f
C4517 a_55228_27815# vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.00123f
C4518 a_42796_23981# a_43750_23544# 0.00231f
C4519 a_4156_5863# a_4852_5960# 0.01227f
C4520 a_52540_15271# a_52452_15368# 0.28563f
C4521 _495_.I a_42820_31048# 0.01411f
C4522 a_932_4392# a_1380_4392# 0.01328f
C4523 _421_.A1 _282_.ZN 0.06528f
C4524 _474_.Q a_48888_19243# 0.30559f
C4525 _388_.B _384_.ZN 0.15205f
C4526 a_54108_15271# a_54556_15271# 0.0131f
C4527 a_5300_15368# VPWR 0.21406f
C4528 _424_.B1 a_47636_25940# 0.00197f
C4529 _436_.ZN a_41476_24776# 0.00168f
C4530 a_21428_22020# a_21516_21976# 0.28563f
C4531 a_17484_21976# a_17932_21976# 0.01288f
C4532 a_66652_2727# a_66564_2824# 0.28563f
C4533 a_35628_16839# a_36076_16839# 0.01288f
C4534 a_33500_15271# VPWR 0.30042f
C4535 a_24876_23544# a_24788_22020# 0.00151f
C4536 a_59620_27208# VPWR 0.82545f
C4537 _250_.ZN a_62763_28776# 0.00603f
C4538 a_66116_17316# VPWR 0.23915f
C4539 a_39572_16936# a_39460_15748# 0.02666f
C4540 _371_.A3 _459_.D 0.00184f
C4541 _251_.A1 a_61836_25515# 0.30428f
C4542 a_31844_23208# a_31932_21543# 0.00151f
C4543 a_47524_1256# a_47972_1256# 0.01328f
C4544 a_30388_23588# a_30476_23544# 0.28563f
C4545 _474_.CLK a_50084_24328# 0.00127f
C4546 _452_.Q a_42392_19243# 0.00164f
C4547 a_3260_7431# VPWR 0.30487f
C4548 a_24080_25227# a_24960_25641# 0.00306f
C4549 a_31284_23588# a_31732_23588# 0.01328f
C4550 a_26916_1256# VPWR 0.22634f
C4551 a_5388_4295# VPWR 0.35526f
C4552 _379_.Z VPWR 0.48929f
C4553 a_26556_2727# a_27004_2727# 0.0131f
C4554 a_62060_13703# a_62420_13800# 0.08707f
C4555 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN VPWR 0.76601f
C4556 a_47972_13800# a_48420_13800# 0.01328f
C4557 a_9635_30644# VPWR 0.18285f
C4558 a_27668_31048# uio_out[0] 0.00268f
C4559 _267_.A2 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.05276f
C4560 a_48844_16839# a_49204_16936# 0.08707f
C4561 _352_.A2 _371_.A1 0.73072f
C4562 _248_.B1 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN 0.06222f
C4563 a_20060_23111# a_20084_22020# 0.0016f
C4564 a_52340_10664# a_52316_9432# 0.0016f
C4565 a_20496_26344# a_21376_26031# 0.00306f
C4566 a_23420_26247# a_23780_26344# 0.08674f
C4567 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_53660_27815# 0.02334f
C4568 a_44612_1636# VPWR 0.20348f
C4569 a_60909_30600# _238_.I 0.0016f
C4570 a_55900_12568# a_55924_12232# 0.00172f
C4571 a_7964_1159# a_7876_1256# 0.28563f
C4572 a_42484_16936# VPWR 0.24746f
C4573 a_26580_23588# a_26556_23111# 0.00172f
C4574 _452_.CLK a_36100_26724# 0.02206f
C4575 a_20620_25112# a_20508_24679# 0.02634f
C4576 a_41440_28363# a_42368_28733# 1.16391f
C4577 _452_.CLK _260_.A2 0.13753f
C4578 a_7652_29860# a_7740_29816# 0.28563f
C4579 a_25792_30301# a_25420_30345# 0.10745f
C4580 a_3708_29816# a_4156_29816# 0.01288f
C4581 a_33860_17316# a_34308_17316# 0.01328f
C4582 a_45956_15368# a_45820_14136# 0.00154f
C4583 a_63516_15271# a_63652_14180# 0.00154f
C4584 a_49764_15368# a_49764_14180# 0.05841f
C4585 a_59172_23588# a_59260_23544# 0.28563f
C4586 a_6980_2824# VPWR 0.20815f
C4587 a_63204_11044# a_63652_11044# 0.01328f
C4588 a_52900_1636# a_52988_1592# 0.28563f
C4589 a_48956_1592# a_49404_1592# 0.01288f
C4590 a_25348_1636# a_25212_1159# 0.00168f
C4591 _287_.A1 a_32904_28776# 0.00179f
C4592 a_33412_20072# a_33412_18884# 0.05841f
C4593 a_58228_27912# a_58020_27508# 0.01565f
C4594 _416_.A1 a_37444_25156# 0.003f
C4595 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN 0.05372f
C4596 _434_.ZN a_39178_23208# 0.0022f
C4597 _452_.D VPWR 0.49824f
C4598 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN a_55228_15704# 0.00103f
C4599 _397_.A2 _284_.A2 0.04436f
C4600 a_52652_18407# a_53012_18504# 0.08717f
C4601 a_54356_18504# a_54444_16839# 0.0027f
C4602 a_53012_18504# VPWR 0.20595f
C4603 _384_.A1 _395_.A3 0.07134f
C4604 a_17036_25112# VPWR 0.29679f
C4605 _303_.ZN a_39780_22805# 0.09748f
C4606 _260_.A1 a_43668_19668# 0.00257f
C4607 _288_.ZN a_38472_30169# 0.00827f
C4608 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I a_63516_19975# 0.00348f
C4609 a_32716_20408# VPWR 0.31594f
C4610 a_14708_27912# a_15156_27912# 0.01328f
C4611 a_26556_30951# VPWR 0.31248f
C4612 _340_.ZN uio_out[3] 0.00265f
C4613 a_3260_12135# VPWR 0.30487f
C4614 a_31620_15748# a_31260_15704# 0.08707f
C4615 _393_.A1 a_45036_28248# 0.00142f
C4616 a_40444_15704# a_40580_15368# 0.00168f
C4617 a_27588_2824# a_28036_2824# 0.01328f
C4618 _304_.B vgaringosc.ro_inv1.inv_array_notouch_\[1\].I 0.00426f
C4619 a_65668_26344# vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN 0.03524f
C4620 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN 0.00353f
C4621 _325_.A1 a_41776_18504# 0.0015f
C4622 _379_.A2 a_18760_29032# 0.41309f
C4623 a_22560_30288# a_22636_29383# 0.01356f
C4624 a_42236_15704# a_42236_15271# 0.05841f
C4625 _437_.A1 _437_.ZN 1.37888f
C4626 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN VPWR 0.84065f
C4627 _304_.B a_52852_24372# 0.03742f
C4628 a_19972_21640# a_19860_20452# 0.02666f
C4629 _256_.A2 _267_.A2 0.00107f
C4630 _452_.CLK a_39660_16839# 0.00245f
C4631 vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I clk 0.00556f
C4632 a_1020_15704# VPWR 0.30073f
C4633 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I a_65072_29860# 0.00568f
C4634 a_40220_20408# a_40220_19975# 0.05841f
C4635 a_52452_15368# VPWR 0.20348f
C4636 _441_.A2 a_42168_22504# 0.0031f
C4637 _247_.ZN _252_.B 0.60367f
C4638 a_24788_22020# a_24428_21976# 0.08707f
C4639 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN 0.64338f
C4640 vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN 0.00647f
C4641 a_55900_15271# VPWR 0.32709f
C4642 _452_.CLK a_37892_17316# 0.00158f
C4643 a_30476_23544# a_30388_22020# 0.00151f
C4644 a_48420_14180# a_48868_14180# 0.01328f
C4645 a_36188_17272# a_36100_15748# 0.00151f
C4646 _304_.B a_43564_27209# 0.00338f
C4647 a_46516_16936# a_46404_15748# 0.02666f
C4648 a_37420_16839# VPWR 0.31389f
C4649 _474_.CLK a_55364_21640# 0.05896f
C4650 a_25652_31048# a_26020_31048# 0.02601f
C4651 hold2.Z _264_.B 0.02787f
C4652 a_49316_1256# VPWR 0.20761f
C4653 a_59172_22020# vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I 0.00318f
C4654 VPWR uo_out[6] 0.97315f
C4655 _328_.A2 a_43892_20072# 0.00145f
C4656 a_62844_14136# a_62756_12612# 0.00151f
C4657 _421_.A1 a_47412_23588# 0.00142f
C4658 a_41048_17341# a_41004_16839# 0.01084f
C4659 _294_.A2 uo_out[3] 0.00189f
C4660 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN a_59172_23208# 0.07148f
C4661 a_28054_30196# VPWR 0.60228f
C4662 a_49740_29383# _392_.A2 0.05465f
C4663 a_35652_17316# VPWR 0.2065f
C4664 a_27004_23111# a_27028_22020# 0.0016f
C4665 _384_.A3 _281_.A1 0.17793f
C4666 _447_.Q a_39772_20408# 0.01451f
C4667 a_50748_1592# VPWR 0.33825f
C4668 a_18940_1159# a_19300_1256# 0.08717f
C4669 a_62956_12135# a_63404_12135# 0.01288f
C4670 _421_.B a_47271_21640# 0.11777f
C4671 a_12356_29480# a_12804_29480# 0.01328f
C4672 a_49292_12135# a_49652_12232# 0.08707f
C4673 a_11996_1592# a_12444_1592# 0.01288f
C4674 a_15940_1636# a_16028_1592# 0.28563f
C4675 _397_.A4 _407_.ZN 0.0398f
C4676 _473_.Q _417_.Z 0.00216f
C4677 a_62308_27912# a_62196_26724# 0.02666f
C4678 _311_.A2 a_38575_24072# 0.0024f
C4679 a_11012_29860# a_10652_29816# 0.08707f
C4680 a_35616_24776# a_36496_24463# 0.00306f
C4681 _358_.A3 a_30796_24463# 0.00125f
C4682 a_56708_15368# a_56708_14180# 0.05841f
C4683 _416_.ZN a_46628_18504# 0.00153f
C4684 a_49316_31048# a_49764_31048# 0.01328f
C4685 a_56260_1636# a_55900_1592# 0.08707f
C4686 a_44160_29123# VPWR 0.18819f
C4687 a_29380_2824# VPWR 0.20348f
C4688 _294_.A2 a_35660_27508# 0.00486f
C4689 _300_.A2 a_38316_20408# 0.0097f
C4690 a_4156_23111# a_4068_23208# 0.28563f
C4691 _362_.ZN _358_.A3 0.26652f
C4692 a_17036_24679# a_16948_24776# 0.28563f
C4693 a_25436_24679# a_25884_24679# 0.012f
C4694 a_33500_19975# a_33948_19975# 0.0131f
C4695 a_1380_9476# VPWR 0.20348f
C4696 a_4068_9096# a_4852_9096# 0.00276f
C4697 _234_.ZN _330_.A1 0.00191f
C4698 a_50212_14180# VPWR 0.2189f
C4699 a_64772_5960# a_65220_5960# 0.01328f
C4700 a_65668_4392# a_66116_4392# 0.01328f
C4701 a_67996_4728# a_67908_3204# 0.0027f
C4702 _303_.ZN a_39796_22504# 0.04265f
C4703 a_4156_18407# a_4852_18504# 0.01227f
C4704 a_35180_18407# a_35628_18407# 0.01255f
C4705 _393_.ZN _393_.A3 0.04786f
C4706 _313_.ZN _304_.A1 0.34111f
C4707 a_37980_15704# a_38564_15748# 0.01675f
C4708 a_64972_12135# VPWR 0.32368f
C4709 a_14148_29480# VPWR 0.20543f
C4710 a_57380_16936# vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN 0.00205f
C4711 _416_.A1 a_45232_25987# 0.00616f
C4712 _340_.ZN a_25962_29480# 0.02383f
C4713 a_42796_23981# a_43246_23610# 0.00209f
C4714 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I VPWR 0.46093f
C4715 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN 0.81205f
C4716 a_53124_15748# a_52988_15271# 0.00168f
C4717 _424_.A2 _281_.ZN 0.15011f
C4718 a_932_24776# VPWR 0.22176f
C4719 a_49180_15704# a_49180_15271# 0.05841f
C4720 a_65668_7528# VPWR 0.21209f
C4721 VPWR uo_out[5] 0.73266f
C4722 a_52852_24372# VPWR 0.79206f
C4723 _281_.A1 a_54824_22045# 0.00108f
C4724 a_67460_4392# VPWR 0.20924f
C4725 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN 0.03848f
C4726 a_1020_19975# a_932_20072# 0.28563f
C4727 a_39908_15748# VPWR 0.20658f
C4728 a_53996_18407# a_54444_18407# 0.01222f
C4729 a_41476_24776# _439_.ZN 0.00268f
C4730 a_31284_22020# a_31732_22020# 0.01328f
C4731 a_30388_22020# a_30476_21976# 0.28563f
C4732 a_49600_30180# _392_.A2 0.00761f
C4733 a_43564_27209# VPWR 0.39907f
C4734 _459_.CLK a_23780_26344# 0.05049f
C4735 _407_.ZN a_51956_26183# 0.00102f
C4736 _294_.A2 a_37291_29535# 0.00355f
C4737 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN a_64100_27912# 0.02176f
C4738 a_41440_28363# a_43132_27815# 0.01084f
C4739 _265_.ZN a_42684_27815# 0.01291f
C4740 _300_.ZN a_40452_23588# 0.00538f
C4741 _398_.C a_50084_24328# 0.45939f
C4742 a_5948_1592# a_6084_1256# 0.00168f
C4743 a_48956_2727# a_49404_2727# 0.0131f
C4744 a_2276_12612# a_2724_12612# 0.01328f
C4745 a_28891_25273# VPWR 0.37218f
C4746 a_47836_17272# a_47948_16839# 0.02634f
C4747 a_51780_17316# a_51756_16839# 0.00172f
C4748 _454_.Q a_24392_28248# 0.44724f
C4749 a_25796_23208# a_25684_22020# 0.02666f
C4750 a_23084_28248# _455_.Q 0.00123f
C4751 _459_.CLK a_40264_30320# 0.02576f
C4752 a_47748_17316# VPWR 0.20897f
C4753 a_64548_1636# VPWR 0.20655f
C4754 a_30364_1159# a_30276_1256# 0.28563f
C4755 a_19300_1636# a_18940_1592# 0.08707f
C4756 a_60268_12135# a_60180_12232# 0.28563f
C4757 _411_.A2 _419_.A4 0.40871f
C4758 a_20508_21543# VPWR 0.31389f
C4759 a_17060_29860# a_16700_29816# 0.0869f
C4760 a_17508_29860# a_17956_29860# 0.01328f
C4761 a_27676_26247# a_27588_26344# 0.28563f
C4762 a_45708_17272# a_46404_17316# 0.01227f
C4763 a_45232_25987# a_45644_26399# 0.00275f
C4764 a_14708_26344# a_14708_25156# 0.05841f
C4765 _416_.A1 a_49740_29383# 0.00941f
C4766 a_34160_20523# a_34308_18884# 0.00149f
C4767 a_47297_25596# _474_.Q 0.5562f
C4768 a_67684_11044# a_67660_10567# 0.00172f
C4769 a_50188_10567# a_50636_10567# 0.01288f
C4770 a_51780_2824# VPWR 0.20815f
C4771 a_62620_1592# a_63068_1592# 0.012f
C4772 clkbuf_1_0__f_clk.I a_47948_23111# 0.00705f
C4773 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN 0.00777f
C4774 _330_.A1 _284_.A2 0.02307f
C4775 a_24092_23111# a_24452_23208# 0.08707f
C4776 a_2724_23208# a_3172_23208# 0.01328f
C4777 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN clk 0.0428f
C4778 a_47860_23208# _324_.B 0.01735f
C4779 _371_.A1 _223_.ZN 0.36295f
C4780 a_55676_28248# _241_.I0 0.00195f
C4781 a_50972_9432# VPWR 0.31444f
C4782 a_20420_2824# a_20508_1159# 0.0027f
C4783 _373_.A2 VPWR 0.99431f
C4784 a_18716_21543# a_19164_21543# 0.01288f
C4785 a_57244_14136# VPWR 0.32088f
C4786 _304_.A1 _316_.ZN 0.00465f
C4787 _424_.B1 a_50212_20452# 0.03713f
C4788 a_10004_31048# a_10116_29860# 0.02666f
C4789 a_8100_29860# a_7964_29383# 0.00168f
C4790 a_58836_12232# VPWR 0.20657f
C4791 a_4156_29816# a_4156_29383# 0.05841f
C4792 a_45284_15748# a_44924_15704# 0.08707f
C4793 a_49764_2824# a_50436_2824# 0.00347f
C4794 _342_.ZN a_23084_29383# 0.00371f
C4795 _473_.Q a_46352_22021# 0.00138f
C4796 a_61860_30736# vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN 0.02628f
C4797 a_33612_24679# VPWR 0.3222f
C4798 a_52360_26355# _412_.ZN 0.27926f
C4799 a_40580_20452# a_40668_20408# 0.28563f
C4800 a_64324_20072# VPWR 0.20554f
C4801 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN a_61972_20452# 0.00558f
C4802 a_10428_2727# a_10340_2824# 0.28563f
C4803 a_53572_15748# VPWR 0.21241f
C4804 a_55452_21543# vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I 0.00608f
C4805 _324_.C _325_.B 0.34628f
C4806 a_49180_9432# a_49628_9432# 0.0131f
C4807 a_51332_9476# a_50972_9432# 0.08717f
C4808 a_26108_30951# uio_out[2] 0.00741f
C4809 a_26468_31048# a_26916_31048# 0.01328f
C4810 a_59732_14180# a_59820_14136# 0.28563f
C4811 a_62084_15368# a_62060_13703# 0.00131f
C4812 a_55452_14136# a_55900_14136# 0.0131f
C4813 _226_.ZN a_41664_22020# 0.01833f
C4814 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN 0.00249f
C4815 a_60909_30600# VPWR 0.78119f
C4816 _402_.A1 _402_.ZN 1.57288f
C4817 _287_.A2 _358_.A3 0.02903f
C4818 a_4068_24776# a_4068_23588# 0.05841f
C4819 a_19612_24679# a_19636_23588# 0.0016f
C4820 a_41340_1159# a_41700_1256# 0.08717f
C4821 a_14684_1159# VPWR 0.29679f
C4822 a_25796_1636# a_26244_1636# 0.01328f
C4823 a_57044_12232# a_57492_12232# 0.01328f
C4824 _419_.A4 _399_.ZN 0.02531f
C4825 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.05143f
C4826 a_17396_21640# VPWR 0.20348f
C4827 a_60285_30600# a_60401_30300# 0.02282f
C4828 _474_.CLK a_52848_25987# 0.00562f
C4829 _352_.A2 a_26220_23544# 0.00277f
C4830 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.00112f
C4831 a_53124_17316# a_52764_17272# 0.08707f
C4832 a_61052_11000# a_61076_10664# 0.00172f
C4833 a_47164_10567# a_47076_10664# 0.28563f
C4834 _251_.ZN a_60516_26344# 0.02582f
C4835 a_56036_23208# VPWR 0.12973f
C4836 _452_.CLK _311_.A2 0.03853f
C4837 a_61948_9432# VPWR 0.31143f
C4838 a_15156_23588# VPWR 0.20348f
C4839 a_62532_20072# a_62980_20072# 0.01328f
C4840 a_64772_6340# VPWR 0.20727f
C4841 a_64660_23588# clk 0.00658f
C4842 a_17036_21543# a_17396_21640# 0.08717f
C4843 a_66564_3204# VPWR 0.20631f
C4844 a_5388_13703# VPWR 0.35526f
C4845 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_58140_26680# 0.0012f
C4846 _452_.CLK a_37067_19001# 0.04074f
C4847 _424_.A2 a_50660_20452# 0.03885f
C4848 _427_.ZN a_54916_21640# 0.01058f
C4849 a_51780_15748# a_52228_15748# 0.01328f
C4850 a_48196_15748# a_48284_15704# 0.28563f
C4851 a_47972_11044# VPWR 0.20348f
C4852 a_35740_25112# VPWR 0.32943f
C4853 _455_.Q a_23060_26724# 0.00909f
C4854 a_40444_2727# a_40580_1636# 0.00154f
C4855 _459_.D a_31820_25112# 0.00423f
C4856 a_67772_21543# a_67684_21640# 0.28563f
C4857 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I _267_.A1 0.06022f
C4858 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN a_63336_29480# 0.17929f
C4859 a_17932_26247# VPWR 0.34464f
C4860 a_21404_2727# a_21764_2824# 0.08717f
C4861 a_3260_9432# a_3260_8999# 0.05841f
C4862 _424_.B1 _475_.Q 0.02055f
C4863 _241_.Z vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.00475f
C4864 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN 0.00375f
C4865 a_29356_21976# a_29268_20452# 0.00151f
C4866 a_63652_14180# a_63740_14136# 0.28563f
C4867 a_16052_20452# a_16500_20452# 0.01328f
C4868 _355_.ZN a_28460_23544# 0.00233f
C4869 _251_.ZN a_59226_25156# 0.02526f
C4870 a_23644_29816# _454_.Q 0.00253f
C4871 _324_.C _402_.B 0.14342f
C4872 a_51196_12568# a_51644_12568# 0.01288f
C4873 a_67572_13800# a_67684_12612# 0.02666f
C4874 _337_.A3 _371_.A2 1.53897f
C4875 a_21764_24776# a_21876_23588# 0.02666f
C4876 _284_.ZN a_43296_28733# 0.07895f
C4877 a_37084_1159# VPWR 0.3289f
C4878 a_52764_1159# a_52676_1256# 0.28563f
C4879 _218_.ZN a_50212_20452# 0.05681f
C4880 a_54040_22366# a_54420_21976# 0.49319f
C4881 a_45956_31048# a_45800_30345# 0.00186f
C4882 _427_.B1 _384_.A1 0.20129f
C4883 a_37444_26344# a_37892_26344# 0.01328f
C4884 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I 0.02152f
C4885 a_58028_10567# a_58388_10664# 0.08707f
C4886 a_4068_10664# a_4852_10664# 0.00276f
C4887 a_12892_1159# a_13340_1159# 0.0131f
C4888 _381_.A2 a_49212_26369# 0.0333f
C4889 _330_.ZN a_38228_16936# 0.00402f
C4890 _370_.B uo_out[6] 0.04401f
C4891 a_54444_19975# VPWR 0.31753f
C4892 a_16052_22020# VPWR 0.20348f
C4893 a_58028_18840# a_58164_18504# 0.00168f
C4894 _459_.Q _459_.D 0.0703f
C4895 a_3620_18884# a_3708_18840# 0.28563f
C4896 a_22636_23544# VPWR 0.3185f
C4897 a_28348_21543# a_28260_21640# 0.28563f
C4898 a_15604_21640# a_16052_21640# 0.01328f
C4899 a_51892_23340# VPWR 0.00829f
C4900 _411_.A2 a_51048_26680# 0.08567f
C4901 a_17148_2727# VPWR 0.31143f
C4902 a_66764_13703# VPWR 0.31431f
C4903 a_47164_30951# uio_in[3] 0.00135f
C4904 a_2276_29860# VPWR 0.20634f
C4905 _260_.A1 _447_.Q 0.03028f
C4906 a_54108_11000# VPWR 0.31436f
C4907 _287_.A1 a_32848_29123# 0.02811f
C4908 _438_.A2 a_39236_26344# 0.04014f
C4909 _244_.Z vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN 0.00135f
C4910 a_19948_26680# VPWR 0.32968f
C4911 _276_.A2 _267_.A2 0.00494f
C4912 a_15692_27815# VPWR 0.29679f
C4913 a_66564_15748# a_66204_15704# 0.0869f
C4914 a_22992_27555# a_22620_27599# 0.10745f
C4915 a_63068_15704# a_63516_15704# 0.0131f
C4916 _416_.A1 hold2.I 0.28216f
C4917 _435_.A3 a_39536_23588# 0.0122f
C4918 _230_.I vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I 0.15917f
C4919 a_32828_2727# a_32740_2824# 0.28563f
C4920 _276_.A2 a_53212_29816# 0.0375f
C4921 a_13700_1256# a_14148_1256# 0.01328f
C4922 a_3260_7864# a_3708_7864# 0.0131f
C4923 a_62308_9476# a_61948_9432# 0.08717f
C4924 _342_.ZN a_24304_29480# 0.00798f
C4925 a_4156_23544# a_4604_23544# 0.01222f
C4926 a_4156_6296# a_4604_6296# 0.01222f
C4927 a_3260_13703# a_3708_13703# 0.0131f
C4928 a_64772_3204# a_65220_3204# 0.01328f
C4929 a_10452_31048# a_10428_29383# 0.00134f
C4930 a_61052_27815# _245_.Z 0.00277f
C4931 a_21652_20452# a_21740_20408# 0.28563f
C4932 a_4156_29383# a_4828_29383# 0.00544f
C4933 a_5276_30951# a_5188_31048# 0.28563f
C4934 a_10564_1636# VPWR 0.21312f
C4935 _421_.A1 _324_.B 1.10723f
C4936 _459_.CLK a_21068_25112# 0.00613f
C4937 a_61076_13800# a_61164_12135# 0.00151f
C4938 _459_.Q a_33524_24776# 0.00152f
C4939 a_58500_12612# a_58140_12568# 0.08707f
C4940 _388_.B a_44252_30951# 0.03716f
C4941 _370_.B uo_out[5] 0.02378f
C4942 _474_.CLK a_56484_23208# 0.0128f
C4943 a_24860_27209# a_25204_26841# 0.00275f
C4944 a_63740_1159# a_64100_1256# 0.08717f
C4945 _268_.A2 _267_.ZN 0.43606f
C4946 a_59484_1159# VPWR 0.29679f
C4947 a_36548_25156# a_36188_25112# 0.0869f
C4948 a_66764_20408# VPWR 0.32938f
C4949 _402_.A1 a_47291_25940# 0.00927f
C4950 a_46180_11044# a_46628_11044# 0.01328f
C4951 a_44276_20072# a_43668_19668# 0.03202f
C4952 _375_.Z a_21740_29383# 0.00315f
C4953 a_67996_18840# VPWR 0.33674f
C4954 _416_.A3 a_47776_20893# 0.00295f
C4955 a_4068_16936# a_4852_16936# 0.00276f
C4956 a_35876_1636# a_35964_1592# 0.28563f
C4957 _258_.I _246_.B2 0.38009f
C4958 a_44476_27815# _470_.D 0.00103f
C4959 a_42596_27912# a_43044_27912# 0.01328f
C4960 _251_.A1 a_56124_28248# 0.00268f
C4961 a_40692_27912# _330_.A1 0.00417f
C4962 _437_.A1 a_37472_24419# 0.03456f
C4963 a_60380_1592# a_60380_1159# 0.05841f
C4964 _268_.A2 _390_.ZN 0.00121f
C4965 a_21316_2824# a_21180_1592# 0.00154f
C4966 a_29716_22020# VPWR 0.21241f
C4967 _455_.Q a_25796_27912# 0.01199f
C4968 a_37196_23544# VPWR 0.31544f
C4969 a_48708_29816# _384_.ZN 0.01436f
C4970 a_33052_18840# a_33500_18840# 0.0131f
C4971 _460_.Q VPWR 3.32826f
C4972 a_39548_2727# VPWR 0.31143f
C4973 a_60628_13800# VPWR 0.20862f
C4974 _218_.ZN _475_.Q 0.17428f
C4975 a_1916_26247# a_2276_26344# 0.08717f
C4976 a_16140_26247# a_16588_26247# 0.0131f
C4977 _392_.A2 VPWR 0.73074f
C4978 _337_.ZN _336_.A2 0.10692f
C4979 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN 0.83895f
C4980 vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN 0.00946f
C4981 a_15940_29860# VPWR 0.21466f
C4982 _294_.A2 _294_.ZN 0.42359f
C4983 a_64884_16936# a_64772_15748# 0.02666f
C4984 a_1020_10567# VPWR 0.30073f
C4985 a_4940_15271# a_5300_15368# 0.08674f
C4986 _237_.A1 a_60276_29032# 0.00298f
C4987 _404_.A1 _400_.ZN 0.43842f
C4988 a_27004_23111# VPWR 0.34784f
C4989 _304_.B _416_.A1 0.15753f
C4990 _411_.A2 _381_.A2 0.05529f
C4991 a_43804_2727# a_44164_2824# 0.08717f
C4992 a_60740_26724# a_60828_26680# 0.28563f
C4993 _452_.CLK a_36660_23588# 0.00154f
C4994 a_66092_16839# a_66004_16936# 0.28563f
C4995 a_63964_18407# a_64412_18407# 0.0131f
C4996 a_20532_23588# a_20172_23544# 0.08707f
C4997 _355_.C a_22620_27599# 0.03446f
C4998 a_63404_20408# a_63428_20072# 0.00172f
C4999 a_2812_25112# a_3260_25112# 0.0131f
C5000 _268_.A2 a_49496_30345# 0.00275f
C5001 a_27028_20452# a_27476_20452# 0.01328f
C5002 a_61636_18504# a_61500_17272# 0.00154f
C5003 a_40580_26344# _435_.A3 0.00116f
C5004 a_1916_16839# a_1828_16936# 0.28563f
C5005 _350_.A1 _462_.D 0.03732f
C5006 a_34304_24029# VPWR 0.19687f
C5007 _402_.A1 a_46068_25156# 0.00744f
C5008 _284_.ZN a_44500_25156# 0.02114f
C5009 _397_.A2 _419_.A4 0.06516f
C5010 a_16700_1592# VPWR 0.30141f
C5011 a_59932_11000# a_59844_9476# 0.00151f
C5012 a_64996_12612# a_65444_12612# 0.01328f
C5013 a_61860_12612# a_61500_12568# 0.08707f
C5014 _474_.CLK ui_in[4] 0.01232f
C5015 _373_.ZN a_28112_27912# 0.00118f
C5016 _230_.I a_58948_26344# 0.00564f
C5017 a_64412_15271# a_64996_15368# 0.01675f
C5018 a_61972_12232# a_61948_11000# 0.0016f
C5019 a_11012_1636# a_10876_1159# 0.00168f
C5020 a_36436_18504# VPWR 0.20757f
C5021 _252_.ZN a_60516_27912# 0.05027f
C5022 a_2724_26724# a_2812_26680# 0.28563f
C5023 a_23108_29860# uio_out[4] 0.00524f
C5024 a_35292_1159# a_35740_1159# 0.0131f
C5025 a_65780_10664# a_66228_10664# 0.01328f
C5026 _330_.ZN a_38842_17316# 0.02604f
C5027 a_31932_26247# a_31844_26344# 0.28563f
C5028 a_2276_20452# VPWR 0.20634f
C5029 _465_.D uio_out[5] 0.75839f
C5030 a_49764_12612# VPWR 0.2124f
C5031 a_61948_2727# VPWR 0.31605f
C5032 a_66988_18407# a_67348_18504# 0.0869f
C5033 a_2812_29383# a_2724_29480# 0.28563f
C5034 a_64748_23544# a_65196_23544# 0.01222f
C5035 a_59260_21976# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.00858f
C5036 a_39236_15368# a_39684_15368# 0.01328f
C5037 a_30724_20072# VPWR 0.22176f
C5038 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN a_56684_18407# 0.00606f
C5039 vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN 0.02759f
C5040 a_2812_15704# a_2812_15271# 0.05841f
C5041 a_62508_10567# VPWR 0.31547f
C5042 _459_.CLK a_31732_25156# 0.01642f
C5043 a_41116_15271# a_41028_15368# 0.28563f
C5044 vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN 0.0192f
C5045 a_60964_26344# vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I 0.00393f
C5046 a_24452_23208# VPWR 0.20622f
C5047 a_63516_17272# a_63540_16936# 0.00172f
C5048 _441_.B _301_.Z 0.00542f
C5049 _416_.A1 VPWR 3.13126f
C5050 a_42684_15271# a_43132_15271# 0.0131f
C5051 a_35008_27533# _358_.A3 0.00242f
C5052 a_25867_26841# VPWR 0.38194f
C5053 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN a_55228_15704# 0.02004f
C5054 _383_.ZN _392_.A2 0.04061f
C5055 _392_.A2 a_50068_27508# 0.00124f
C5056 a_38876_19975# a_39236_20072# 0.0869f
C5057 _330_.A1 _450_.D 1.12301f
C5058 a_55228_2727# a_55140_2824# 0.28563f
C5059 a_66652_17272# a_67100_17272# 0.01255f
C5060 _284_.ZN a_39300_31048# 0.00873f
C5061 _260_.A2 _447_.Q 0.00635f
C5062 _452_.CLK a_42684_27815# 0.00103f
C5063 a_36100_1256# a_36548_1256# 0.01328f
C5064 a_24340_23588# a_23980_23544# 0.08717f
C5065 a_20868_23208# a_20956_21543# 0.00151f
C5066 a_27028_23588# a_27476_23588# 0.01328f
C5067 a_4068_1256# VPWR 0.22181f
C5068 a_4740_31048# VPWR 0.22891f
C5069 a_19188_25156# a_18828_25112# 0.08707f
C5070 _251_.A1 a_56836_27208# 0.00164f
C5071 a_15132_2727# a_15580_2727# 0.0131f
C5072 a_34080_22461# VPWR 0.19703f
C5073 a_51084_13703# a_51444_13800# 0.08707f
C5074 a_64972_13703# a_65420_13703# 0.0131f
C5075 _476_.Q a_50748_20408# 0.01048f
C5076 a_51240_23340# a_51892_23340# 0.00195f
C5077 _250_.A2 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.03845f
C5078 a_32628_20452# a_32716_20408# 0.28563f
C5079 a_59172_26724# a_59036_26247# 0.00168f
C5080 a_18180_31048# _379_.A2 0.00149f
C5081 a_37868_16839# a_38228_16936# 0.08707f
C5082 a_61412_27912# _245_.Z 0.00308f
C5083 a_30364_1592# VPWR 0.29679f
C5084 a_62284_16839# VPWR 0.31594f
C5085 a_41116_1592# a_41252_1256# 0.00168f
C5086 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN VPWR 1.03183f
C5087 a_55116_10567# a_55140_9476# 0.0016f
C5088 a_2276_1636# a_1916_1592# 0.08707f
C5089 _478_.D a_54804_24776# 0.00202f
C5090 a_4156_25112# a_4156_24679# 0.05841f
C5091 _384_.ZN _402_.A1 0.67598f
C5092 _473_.Q a_49652_20936# 0.00456f
C5093 _438_.A2 _304_.A1 0.04454f
C5094 a_60964_27912# a_61052_26247# 0.0027f
C5095 a_40668_26247# _260_.A1 0.00149f
C5096 a_2276_17316# a_2724_17316# 0.01328f
C5097 a_53108_21640# VPWR 0.00419f
C5098 a_33956_31048# uo_out[4] 0.00135f
C5099 a_59844_11044# a_60292_11044# 0.01328f
C5100 a_56260_11044# a_56348_11000# 0.28563f
C5101 vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN 0.75747f
C5102 a_51220_16936# a_51668_16936# 0.01328f
C5103 _316_.A3 a_34716_20937# 0.00795f
C5104 a_45596_1592# a_46044_1592# 0.01288f
C5105 _324_.B a_48921_22020# 0.00271f
C5106 _427_.B1 clk 0.06089f
C5107 _294_.A2 a_30778_31048# 0.00898f
C5108 a_20756_26724# a_20396_26680# 0.08663f
C5109 a_19860_26724# _455_.D 0.00244f
C5110 a_45644_26399# VPWR 0.00246f
C5111 a_59652_25640# a_60416_25156# 0.00399f
C5112 a_64772_26344# a_65668_26344# 0.0023f
C5113 a_49896_18909# VPWR 1.13505f
C5114 _336_.A2 a_27924_24776# 0.01247f
C5115 a_21292_20408# VPWR 0.31143f
C5116 a_4940_27815# a_5388_27815# 0.01222f
C5117 a_62532_30736# ui_in[2] 0.00215f
C5118 a_35652_25156# _444_.D 0.00155f
C5119 _397_.A2 a_48820_28292# 0.01075f
C5120 _451_.Q a_38340_21327# 0.49385f
C5121 _451_.Q _432_.ZN 0.34651f
C5122 a_1380_15748# a_1468_15704# 0.28563f
C5123 a_55900_12568# VPWR 0.31389f
C5124 _355_.C a_25936_25597# 0.07595f
C5125 _247_.ZN _243_.B2 0.00595f
C5126 a_16164_2824# a_16612_2824# 0.01328f
C5127 _355_.C uio_out[5] 0.28944f
C5128 a_13788_29383# a_14148_29480# 0.08717f
C5129 _379_.A2 a_18816_29931# 0.0047f
C5130 a_53660_21543# a_53572_21640# 0.28563f
C5131 a_19328_28733# a_19948_27815# 0.02396f
C5132 _324_.C a_46352_22021# 0.00861f
C5133 a_52092_15271# a_52452_15368# 0.08717f
C5134 a_2364_8999# a_2276_9096# 0.28563f
C5135 _419_.A4 a_47860_21640# 0.13394f
C5136 a_3260_7431# a_3172_7528# 0.28563f
C5137 a_56372_10664# VPWR 0.21565f
C5138 _495_.I a_41922_31073# 0.03123f
C5139 a_55676_27815# a_55588_27912# 0.28563f
C5140 a_4156_5863# a_4068_5960# 0.28563f
C5141 a_42796_23981# a_43126_24119# 0.75472f
C5142 a_5388_4295# a_5300_4392# 0.28563f
C5143 a_3620_21640# a_3620_20452# 0.05841f
C5144 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I 0.11314f
C5145 _255_.ZN _246_.B2 0.16013f
C5146 _474_.Q a_48084_18884# 0.00699f
C5147 a_4852_15368# VPWR 0.22733f
C5148 _436_.ZN a_40973_24776# 0.00105f
C5149 _398_.C _397_.Z 0.02467f
C5150 a_21428_22020# a_21068_21976# 0.08707f
C5151 a_33052_15271# VPWR 0.29736f
C5152 a_66204_2727# a_66564_2824# 0.0869f
C5153 _300_.A2 _301_.Z 0.26714f
C5154 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN a_67684_21640# 0.02057f
C5155 _275_.A2 _268_.A2 0.20072f
C5156 a_2276_14180# a_2724_14180# 0.01328f
C5157 a_59260_26680# VPWR 0.332f
C5158 a_65668_17316# VPWR 0.21723f
C5159 a_29804_23544# a_30476_23544# 0.00544f
C5160 _416_.A1 _383_.ZN 0.0263f
C5161 a_2812_7431# VPWR 0.30213f
C5162 a_24080_25227# a_24468_25641# 0.00393f
C5163 a_26468_1256# VPWR 0.2098f
C5164 a_4940_4295# VPWR 0.31945f
C5165 a_25008_25597# a_25643_25273# 0.02112f
C5166 a_62060_13703# a_61972_13800# 0.28563f
C5167 a_65756_26247# VPWR 0.35714f
C5168 a_17148_29383# VPWR 0.30117f
C5169 a_30812_17272# a_30812_16839# 0.05841f
C5170 a_34756_17316# a_34732_16839# 0.00172f
C5171 a_41536_17636# a_41948_17433# 0.00275f
C5172 a_9084_30951# VPWR 0.32308f
C5173 _330_.A1 _419_.A4 0.00755f
C5174 _274_.A2 a_52756_29076# 0.3575f
C5175 a_48844_16839# a_48756_16936# 0.28563f
C5176 a_932_23208# a_932_22020# 0.05841f
C5177 a_7516_1159# a_7876_1256# 0.08717f
C5178 a_20496_26344# a_20884_26031# 0.00393f
C5179 a_23420_26247# a_23332_26344# 0.28563f
C5180 a_41812_16936# VPWR 0.21858f
C5181 a_44164_1636# VPWR 0.20348f
C5182 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I a_65308_19975# 0.03018f
C5183 a_65980_12568# a_65868_12135# 0.02634f
C5184 a_932_29480# a_1380_29480# 0.01328f
C5185 a_51980_12135# a_52428_12135# 0.01288f
C5186 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN a_57916_25112# 0.00204f
C5187 a_23084_23544# a_23196_23111# 0.02634f
C5188 _452_.CLK a_35140_26680# 0.04208f
C5189 a_8772_1636# a_9220_1636# 0.01328f
C5190 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN a_57940_20452# 0.00294f
C5191 a_7652_29860# a_7292_29816# 0.08707f
C5192 _247_.ZN a_59172_26724# 0.00219f
C5193 _474_.D a_50860_18407# 0.00265f
C5194 a_58252_18407# a_58388_17316# 0.00154f
C5195 a_6532_2824# VPWR 0.20815f
C5196 a_49852_11000# a_49740_10567# 0.02634f
C5197 a_52900_1636# a_52540_1592# 0.08707f
C5198 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I VPWR 0.84647f
C5199 _452_.CLK _319_.ZN 0.13308f
C5200 a_41776_18504# VPWR 0.01536f
C5201 a_52652_18407# a_52564_18504# 0.28563f
C5202 _373_.A2 a_28556_29167# 0.00874f
C5203 a_57468_1159# a_58140_1159# 0.00544f
C5204 a_66228_20452# a_66676_20452# 0.01328f
C5205 a_52564_18504# VPWR 0.20595f
C5206 a_66204_18840# a_66652_18840# 0.01255f
C5207 a_16588_25112# VPWR 0.29679f
C5208 a_32268_20408# VPWR 0.31594f
C5209 _324_.B a_49034_21640# 0.00487f
C5210 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I a_63068_19975# 0.03017f
C5211 _359_.B uo_out[4] 0.00421f
C5212 _365_.ZN uo_out[2] 0.00594f
C5213 a_26108_30951# VPWR 0.31244f
C5214 a_2812_12135# VPWR 0.30213f
C5215 a_34756_15748# a_35204_15748# 0.01328f
C5216 a_31172_15748# a_31260_15704# 0.28563f
C5217 _267_.A2 _238_.ZN 0.00192f
C5218 _397_.A4 _279_.Z 0.57671f
C5219 _412_.A1 _412_.B2 0.00127f
C5220 a_28348_21543# a_28372_20452# 0.0016f
C5221 a_65668_26344# clk 0.00125f
C5222 _452_.CLK a_39212_16839# 0.00239f
C5223 a_38764_20408# _327_.Z 0.0012f
C5224 a_64324_29860# a_65072_29860# 0.00235f
C5225 a_4964_15748# VPWR 0.21167f
C5226 a_52004_15368# VPWR 0.20348f
C5227 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN a_55900_15271# 0.00199f
C5228 a_49988_21236# a_50660_20452# 0.00171f
C5229 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I VPWR 0.97537f
C5230 a_53704_23219# a_54824_22045# 0.00136f
C5231 a_27924_22020# a_28372_22020# 0.01328f
C5232 a_24340_22020# a_24428_21976# 0.28563f
C5233 a_55452_15271# VPWR 0.32921f
C5234 a_46156_16839# a_46604_16839# 0.01288f
C5235 _452_.CLK a_37444_17316# 0.00645f
C5236 a_36972_16839# VPWR 0.31431f
C5237 _474_.CLK a_54916_21640# 0.01693f
C5238 a_48868_1256# VPWR 0.2062f
C5239 a_58500_1256# a_58948_1256# 0.01328f
C5240 _427_.B2 _419_.Z 0.01879f
C5241 a_25652_31048# a_25012_31048# 0.00782f
C5242 a_25100_30951# a_26020_31048# 0.00375f
C5243 _421_.A1 a_47172_23588# 0.00287f
C5244 a_58836_13800# a_59284_13800# 0.01328f
C5245 a_37532_2727# a_37980_2727# 0.0131f
C5246 _424_.B2 a_49896_18909# 0.00183f
C5247 a_26427_29977# VPWR 0.3827f
C5248 a_35204_17316# VPWR 0.21636f
C5249 _447_.Q a_39333_20936# 0.00929f
C5250 a_50300_1592# VPWR 0.35877f
C5251 _245_.Z _251_.ZN 0.02791f
C5252 a_18940_1159# a_18852_1256# 0.28563f
C5253 _474_.CLK _284_.B 0.00322f
C5254 a_18628_23208# a_18740_22020# 0.02666f
C5255 _451_.Q _260_.A1 1.69036f
C5256 a_62844_12568# a_62868_12232# 0.00172f
C5257 a_49292_12135# a_49204_12232# 0.28563f
C5258 a_15940_1636# a_15580_1592# 0.08663f
C5259 _421_.B a_47047_21640# 0.02811f
C5260 a_14148_29860# a_14596_29860# 0.01328f
C5261 a_10564_29860# a_10652_29816# 0.28563f
C5262 a_36636_17272# a_37084_17272# 0.01288f
C5263 _358_.A3 a_31168_24419# 0.00174f
C5264 _251_.ZN a_60604_26247# 0.00509f
C5265 _416_.ZN a_46180_18504# 0.00124f
C5266 a_66428_11000# a_66876_11000# 0.01288f
C5267 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I a_67684_24776# 0.04407f
C5268 a_28932_2824# VPWR 0.20348f
C5269 a_55812_1636# a_55900_1592# 0.28563f
C5270 a_59396_1636# a_59844_1636# 0.01328f
C5271 _303_.ZN _304_.ZN 1.04746f
C5272 a_24988_23111# a_25436_23111# 0.01288f
C5273 a_3708_23111# a_4068_23208# 0.08717f
C5274 _284_.ZN _324_.C 0.04856f
C5275 a_16588_24679# a_16948_24776# 0.08717f
C5276 _452_.CLK _460_.D 0.0023f
C5277 a_18028_28777# uio_out[7] 0.01787f
C5278 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I a_55228_15704# 0.0036f
C5279 a_40038_28720# _330_.A1 0.00145f
C5280 a_8996_2824# a_9084_1159# 0.0027f
C5281 a_49764_14180# VPWR 0.20967f
C5282 _231_.I vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN 0.0303f
C5283 a_4156_18407# a_4068_18504# 0.28563f
C5284 a_36636_26680# a_36636_26247# 0.05841f
C5285 a_33376_23659# _304_.A1 0.00728f
C5286 a_1828_31048# a_1828_29860# 0.05841f
C5287 _351_.ZN a_25524_26344# 0.0018f
C5288 a_26020_31048# a_25420_30345# 0.01033f
C5289 a_63336_29480# VPWR 0.40866f
C5290 a_13700_29480# VPWR 0.20348f
C5291 a_64300_12135# VPWR 0.34599f
C5292 _397_.A2 _381_.A2 1.25825f
C5293 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_65668_26344# 0.00354f
C5294 _416_.A1 a_44744_26355# 0.02761f
C5295 a_26108_2727# a_26244_1636# 0.00154f
C5296 a_38340_2824# a_39012_2824# 0.00347f
C5297 _229_.I ui_in[0] 0.02219f
C5298 _424_.A2 a_46156_25112# 0.0085f
C5299 a_28012_24679# VPWR 0.32279f
C5300 a_51332_24372# VPWR 0.83623f
C5301 a_67012_4392# VPWR 0.20348f
C5302 a_65220_7528# VPWR 0.20921f
C5303 _252_.B _251_.ZN 0.26408f
C5304 a_26916_21640# a_27028_20452# 0.02666f
C5305 _384_.ZN _424_.B1 0.01005f
C5306 a_39460_15748# VPWR 0.20677f
C5307 _241_.I0 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.02817f
C5308 _459_.Q _359_.ZN 0.01193f
C5309 a_45284_9476# a_45732_9476# 0.01328f
C5310 a_29804_21976# a_30476_21976# 0.00544f
C5311 a_49112_29885# _392_.A2 0.01754f
C5312 a_43936_27165# VPWR 0.18743f
C5313 _448_.D a_35936_19001# 0.00159f
C5314 _327_.Z a_37360_19325# 0.006f
C5315 a_51196_14136# a_51644_14136# 0.01288f
C5316 _281_.ZN clkbuf_1_0__f_clk.I 1.04573f
C5317 _305_.A2 _324_.B 1.33514f
C5318 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN VPWR 0.76465f
C5319 _265_.ZN a_42236_27815# 0.0522f
C5320 _294_.A2 a_36284_29167# 0.00252f
C5321 _459_.CLK a_23332_26344# 0.01108f
C5322 a_35140_26680# a_34448_25597# 0.00146f
C5323 _230_.I _247_.B 0.00653f
C5324 a_29184_25597# VPWR 0.51617f
C5325 _474_.CLK _474_.D 0.00212f
C5326 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _407_.ZN 0.01314f
C5327 _311_.A2 _447_.Q 0.03104f
C5328 a_47300_17316# VPWR 0.20909f
C5329 _294_.A2 _362_.B 0.86566f
C5330 a_66676_10664# a_66652_9432# 0.0016f
C5331 a_29916_1159# a_30276_1256# 0.08717f
C5332 a_57244_12568# a_57156_11044# 0.00151f
C5333 a_59820_12135# a_60180_12232# 0.08707f
C5334 a_45732_12232# a_46180_12232# 0.01328f
C5335 a_64100_1636# VPWR 0.20363f
C5336 _265_.ZN _284_.B 0.00114f
C5337 _386_.ZN _384_.ZN 0.09171f
C5338 a_31372_23544# a_31396_23208# 0.00172f
C5339 a_22436_1636# a_22884_1636# 0.01328f
C5340 a_18852_1636# a_18940_1592# 0.28563f
C5341 a_56596_23588# a_56572_23111# 0.00172f
C5342 a_20060_21543# VPWR 0.31389f
C5343 a_16612_29860# a_16700_29816# 0.28563f
C5344 a_27228_26247# a_27588_26344# 0.08674f
C5345 a_19612_26247# a_19636_25156# 0.0016f
C5346 a_51332_2824# VPWR 0.20815f
C5347 a_63740_11000# a_63852_10567# 0.02634f
C5348 a_53660_11000# a_53684_10664# 0.00172f
C5349 a_39100_1592# a_39100_1159# 0.05841f
C5350 _251_.A1 a_58020_27508# 0.00105f
C5351 a_24092_23111# a_24004_23208# 0.28563f
C5352 a_19076_24776# a_19524_24776# 0.01328f
C5353 a_30388_28776# _223_.ZN 0.10748f
C5354 a_56516_26344# clk 0.00276f
C5355 a_55676_28248# a_56124_28248# 0.012f
C5356 _460_.Q _360_.ZN 0.61644f
C5357 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I _243_.A1 0.00282f
C5358 _427_.B2 _424_.A1 0.26024f
C5359 a_50524_9432# VPWR 0.35477f
C5360 a_56796_14136# VPWR 0.3337f
C5361 a_28672_31048# VPWR 0.01471f
C5362 a_56484_2824# a_56348_1592# 0.00154f
C5363 a_60292_2824# a_60292_1636# 0.05841f
C5364 _304_.A1 a_33152_22091# 0.00572f
C5365 _427_.A2 _427_.ZN 0.45302f
C5366 a_34644_18504# a_35092_18504# 0.01328f
C5367 _294_.A2 a_32628_26725# 0.00162f
C5368 a_43232_29480# a_43620_29167# 0.00393f
C5369 a_58388_12232# VPWR 0.23551f
C5370 a_40892_15704# a_41340_15704# 0.01288f
C5371 a_44836_15748# a_44924_15704# 0.28563f
C5372 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I 0.66988f
C5373 a_40580_20452# a_40220_20408# 0.08663f
C5374 a_63316_23208# vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I 0.00187f
C5375 a_33164_24679# VPWR 0.32788f
C5376 a_63876_20072# VPWR 0.20348f
C5377 a_34308_21640# a_34160_20523# 0.00179f
C5378 a_9980_2727# a_10340_2824# 0.08717f
C5379 a_53124_15748# VPWR 0.20622f
C5380 a_62172_19975# a_62620_19975# 0.0131f
C5381 a_50884_9476# a_50972_9432# 0.28563f
C5382 a_25652_31048# uio_out[2] 0.09646f
C5383 a_59732_14180# a_59372_14136# 0.0869f
C5384 _447_.Q a_37444_21640# 0.02569f
C5385 _448_.Q _325_.A2 0.09536f
C5386 ui_in[0] rst_n 0.06702f
C5387 a_60285_30600# VPWR 0.57405f
C5388 a_59932_2727# a_60380_2727# 0.0131f
C5389 _416_.A1 a_49112_29885# 0.00135f
C5390 a_47972_12612# a_48420_12612# 0.01328f
C5391 _439_.ZN _441_.B 0.04008f
C5392 a_59620_23208# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.002f
C5393 _416_.A1 _260_.ZN 0.00174f
C5394 _431_.A3 VPWR 0.87254f
C5395 _398_.C _284_.B 0.02508f
C5396 a_31396_23208# a_31372_21976# 0.0016f
C5397 a_3172_12232# a_3172_11044# 0.05841f
C5398 a_3620_20072# a_4068_20072# 0.01328f
C5399 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_63404_23544# 0.01345f
C5400 a_14236_1159# VPWR 0.29679f
C5401 a_41340_1159# a_41252_1256# 0.28563f
C5402 _324_.C vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.00127f
C5403 a_24304_26795# a_25184_27209# 0.00306f
C5404 _294_.ZN a_32580_27912# 0.00322f
C5405 a_64324_5960# a_64324_4772# 0.05841f
C5406 a_65220_4392# a_65220_3204# 0.05841f
C5407 _474_.CLK a_52360_26355# 0.0291f
C5408 _352_.A2 a_25772_23544# 0.00277f
C5409 a_16948_21640# VPWR 0.20348f
C5410 a_48732_17272# a_49180_17272# 0.01288f
C5411 a_52676_17316# a_52764_17272# 0.28563f
C5412 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I 0.0051f
C5413 a_53212_15704# a_53124_14180# 0.0027f
C5414 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_58476_13703# 0.03465f
C5415 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I VPWR 0.73556f
C5416 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I 0.69814f
C5417 a_60716_10567# a_61164_10567# 0.01288f
C5418 a_46716_10567# a_47076_10664# 0.08717f
C5419 a_1468_1159# a_1916_1159# 0.0131f
C5420 a_46044_1592# a_46044_1159# 0.05841f
C5421 _454_.Q a_23920_27555# 0.17891f
C5422 a_6980_2824# a_6844_1592# 0.00154f
C5423 _443_.D _330_.A1 0.40287f
C5424 _251_.ZN a_60013_26344# 0.00765f
C5425 a_22660_23208# a_23108_23208# 0.01328f
C5426 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN a_54780_18840# 0.00769f
C5427 a_58388_18884# a_58836_18884# 0.01328f
C5428 a_31168_24419# a_31803_24831# 0.02112f
C5429 a_30240_24776# a_32096_24419# 0.02307f
C5430 _452_.CLK a_37532_25112# 0.00111f
C5431 _451_.Q _260_.A2 0.4533f
C5432 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN 0.00638f
C5433 a_61500_9432# VPWR 0.31143f
C5434 _384_.ZN _218_.ZN 0.00333f
C5435 a_14708_23588# VPWR 0.22176f
C5436 a_64324_6340# VPWR 0.22383f
C5437 a_31396_2824# a_31484_1159# 0.0027f
C5438 a_4940_13703# VPWR 0.31945f
C5439 a_17036_21543# a_16948_21640# 0.28563f
C5440 a_64212_23588# clk 0.00658f
C5441 a_66116_3204# VPWR 0.23643f
C5442 a_29244_21543# a_29692_21543# 0.01288f
C5443 _424_.A2 a_50212_20452# 0.00189f
C5444 a_17732_31048# a_17596_29816# 0.00154f
C5445 _452_.CLK a_37360_19325# 0.00721f
C5446 _427_.ZN a_54468_21640# 0.01058f
C5447 _419_.A4 a_47483_20569# 0.03107f
C5448 a_48196_15748# a_47836_15704# 0.08707f
C5449 a_31348_25156# VPWR 0.0068f
C5450 a_47524_11044# VPWR 0.20348f
C5451 a_60740_2824# a_61188_2824# 0.01328f
C5452 a_31732_25156# a_31820_25112# 0.28563f
C5453 a_11091_30644# a_11012_29860# 0.03636f
C5454 a_67884_19975# a_67796_20072# 0.28563f
C5455 _336_.A2 a_27588_26344# 0.00335f
C5456 _252_.ZN a_59652_25640# 0.00154f
C5457 _285_.Z _459_.CLK 0.0472f
C5458 _346_.B VPWR 0.76498f
C5459 a_37196_23544# _311_.Z 0.00205f
C5460 a_34396_18840# VPWR 0.3563f
C5461 a_17484_26247# VPWR 0.29719f
C5462 a_21404_2727# a_21316_2824# 0.28563f
C5463 a_49852_30951# _392_.A2 0.00208f
C5464 _379_.Z _378_.I 0.00153f
C5465 a_56124_9432# a_56708_9476# 0.01675f
C5466 _436_.B a_41228_27815# 0.00262f
C5467 a_2276_1256# a_2724_1256# 0.01328f
C5468 a_2724_31048# a_3172_31048# 0.01328f
C5469 _474_.Q a_51240_20452# 0.0038f
C5470 a_63652_14180# a_63292_14136# 0.08707f
C5471 a_66788_14180# a_67236_14180# 0.01328f
C5472 _355_.ZN a_28012_23544# 0.00715f
C5473 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN 0.96926f
C5474 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN 0.78908f
C5475 _430_.ZN a_39536_23588# 0.00113f
C5476 _337_.A3 a_26954_28776# 0.00406f
C5477 a_19836_1592# a_19972_1256# 0.00168f
C5478 _324_.C a_46356_24072# 0.39769f
C5479 a_63764_13800# a_63740_12568# 0.0016f
C5480 a_50100_13800# a_50188_12135# 0.00151f
C5481 _480_.Q a_43003_28409# 0.00376f
C5482 a_60276_29032# a_60156_27815# 0.00111f
C5483 a_52316_1159# a_52676_1256# 0.08717f
C5484 a_36636_1159# VPWR 0.3289f
C5485 _284_.ZN a_41996_28777# 0.01212f
C5486 a_51444_12232# a_51556_11044# 0.02666f
C5487 a_67572_12232# a_68020_12232# 0.01328f
C5488 a_28572_1592# a_29020_1592# 0.01288f
C5489 _467_.D a_15156_26724# 0.00137f
C5490 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.02867f
C5491 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN 0.73436f
C5492 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I VPWR 0.94475f
C5493 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I 0.07208f
C5494 _284_.ZN a_38472_30169# 0.49316f
C5495 a_58028_10567# a_57940_10664# 0.28563f
C5496 _381_.A2 a_48988_26369# 0.02338f
C5497 _330_.ZN a_37780_16936# 0.00196f
C5498 a_52408_19759# VPWR 0.1873f
C5499 a_32240_31048# uo_out[6] 0.00259f
C5500 a_15604_22020# VPWR 0.20348f
C5501 _459_.Q a_31732_25156# 0.01615f
C5502 a_28372_23588# VPWR 0.2066f
C5503 a_27900_21543# a_28260_21640# 0.08707f
C5504 a_66316_13703# VPWR 0.32333f
C5505 a_16700_2727# VPWR 0.31143f
C5506 a_3620_18884# a_3260_18840# 0.08717f
C5507 a_1020_18840# a_1468_18840# 0.0131f
C5508 a_51668_23340# VPWR 0.00743f
C5509 a_1828_29860# VPWR 0.20348f
C5510 a_61052_26247# vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I 0.00374f
C5511 a_45012_29816# VPWR 0.36854f
C5512 _287_.A1 a_31920_29480# 0.03256f
C5513 a_53660_11000# VPWR 0.31436f
C5514 a_38336_18147# a_38971_18559# 0.02112f
C5515 a_54692_15748# a_55140_15748# 0.01328f
C5516 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN a_58500_26344# 0.00636f
C5517 _384_.ZN _386_.A4 0.00898f
C5518 _324_.B a_48321_23208# 0.24512f
C5519 a_66116_15748# a_66204_15704# 0.28563f
C5520 _438_.A2 a_40004_22020# 0.00464f
C5521 _448_.D a_36836_20072# 0.0018f
C5522 a_15244_27815# VPWR 0.29679f
C5523 _435_.A3 a_39332_23588# 0.00391f
C5524 a_32380_2727# a_32740_2824# 0.08717f
C5525 _276_.A2 a_52073_30344# 0.00761f
C5526 a_61860_9476# a_61948_9432# 0.28563f
C5527 _424_.A2 _475_.Q 0.1483f
C5528 _342_.ZN a_24100_29480# 0.00223f
C5529 a_60604_27815# _245_.Z 0.00203f
C5530 a_19500_20408# a_19948_20408# 0.0131f
C5531 a_21652_20452# a_21292_20408# 0.08717f
C5532 a_58476_18840# a_58388_17316# 0.0027f
C5533 a_4828_30951# a_5188_31048# 0.0869f
C5534 a_26780_1592# a_26916_1256# 0.00168f
C5535 a_58052_12612# a_58140_12568# 0.28563f
C5536 a_54108_12568# a_54556_12568# 0.01288f
C5537 a_5052_12568# a_4940_12135# 0.02634f
C5538 a_10116_1636# VPWR 0.21153f
C5539 _478_.D a_54892_23544# 0.01674f
C5540 _459_.Q a_33076_24776# 0.12434f
C5541 _459_.CLK a_20620_25112# 0.00613f
C5542 _388_.B a_43804_30951# 0.0196f
C5543 a_32240_31048# uo_out[5] 0.02959f
C5544 a_43716_31048# a_43828_29860# 0.02666f
C5545 a_9308_29816# a_9444_29480# 0.00168f
C5546 a_25348_24776# a_25324_23544# 0.0016f
C5547 a_66316_20408# VPWR 0.33818f
C5548 a_59036_1159# VPWR 0.29679f
C5549 a_35092_18504# a_35180_16839# 0.00151f
C5550 a_63740_1159# a_63652_1256# 0.28563f
C5551 a_36100_25156# a_36188_25112# 0.28563f
C5552 a_54580_12232# a_54556_11000# 0.0016f
C5553 a_35876_1636# a_35516_1592# 0.08707f
C5554 a_67548_18840# VPWR 0.31547f
C5555 a_58388_12232# a_58500_11044# 0.02666f
C5556 _416_.A3 a_46476_20937# 0.03587f
C5557 _398_.C a_52360_26355# 0.00914f
C5558 _258_.I a_57220_29861# 0.00185f
C5559 a_39796_27912# _330_.A1 0.00865f
C5560 a_54580_10664# a_55028_10664# 0.01328f
C5561 a_23868_1159# a_24316_1159# 0.0131f
C5562 _437_.A1 a_37179_24831# 0.01476f
C5563 a_61300_15748# a_61276_15271# 0.00172f
C5564 _355_.C _373_.ZN 1.13669f
C5565 a_29268_22020# VPWR 0.20669f
C5566 _287_.A2 _362_.ZN 0.04393f
C5567 a_36748_23544# VPWR 0.31415f
C5568 a_26468_21640# a_26916_21640# 0.01328f
C5569 _285_.Z uo_out[7] 0.15386f
C5570 a_39100_2727# VPWR 0.31605f
C5571 a_53572_2824# a_53660_1159# 0.0027f
C5572 a_60180_13800# VPWR 0.20595f
C5573 _467_.D uio_out[7] 0.00705f
C5574 _436_.ZN _452_.Q 0.06638f
C5575 a_1916_26247# a_1828_26344# 0.28563f
C5576 a_2724_15368# a_3172_15368# 0.01328f
C5577 a_15492_29860# VPWR 0.20646f
C5578 _474_.CLK _395_.A2 0.09357f
C5579 a_67772_11000# VPWR 0.33562f
C5580 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN 0.17932f
C5581 a_4940_15271# a_4852_15368# 0.28563f
C5582 _452_.CLK a_42392_19243# 0.00703f
C5583 a_26556_23111# VPWR 0.32672f
C5584 _424_.B1 a_51576_25896# 0.00165f
C5585 a_34715_22137# a_35000_22137# 0.00277f
C5586 a_31260_15271# a_31708_15271# 0.0131f
C5587 a_67996_17272# a_67908_15748# 0.00151f
C5588 a_60740_26724# a_59620_27208# 0.07589f
C5589 _325_.ZN a_44752_18147# 0.00565f
C5590 a_43804_2727# a_43716_2824# 0.28563f
C5591 _294_.A2 a_35914_28776# 0.0019f
C5592 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I _324_.C 0.02254f
C5593 a_63876_17316# a_64324_17316# 0.01328f
C5594 _452_.CLK a_36212_23588# 0.00306f
C5595 _441_.B _303_.ZN 0.18706f
C5596 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I 0.07109f
C5597 a_29563_29535# a_29848_29535# 0.00277f
C5598 a_65420_16839# a_66004_16936# 0.01675f
C5599 a_67100_9432# a_67548_9432# 0.0131f
C5600 a_1020_7431# a_1468_7431# 0.0131f
C5601 a_64412_7864# a_64412_7431# 0.05841f
C5602 a_20084_23588# a_20172_23544# 0.28563f
C5603 _459_.CLK _371_.A1 0.07073f
C5604 a_24676_1256# a_25124_1256# 0.01328f
C5605 _355_.C a_22992_27555# 0.02838f
C5606 a_4964_25156# a_5052_25112# 0.28563f
C5607 a_16140_23544# a_16588_23544# 0.01288f
C5608 _284_.ZN a_43580_27815# 0.03914f
C5609 a_2812_4295# a_3260_4295# 0.0131f
C5610 a_66204_4728# a_66204_4295# 0.05841f
C5611 a_65308_6296# a_65308_5863# 0.05841f
C5612 a_1916_5863# a_2364_5863# 0.0131f
C5613 a_67772_14136# a_67660_13703# 0.02634f
C5614 a_49764_31048# a_49496_30345# 0.01055f
C5615 a_3708_2727# a_4156_2727# 0.0131f
C5616 a_53772_13703# a_54220_13703# 0.01288f
C5617 _268_.A2 a_49600_30180# 0.00434f
C5618 a_35988_16936# a_35964_15271# 0.00134f
C5619 _459_.Q a_35108_28776# 0.00122f
C5620 _355_.C _465_.D 0.95451f
C5621 _424_.B2 a_52408_19759# 0.02938f
C5622 a_15132_29383# a_15580_29383# 0.0131f
C5623 _350_.A1 a_36288_31048# 0.00232f
C5624 a_1468_16839# a_1828_16936# 0.08717f
C5625 _284_.ZN a_44028_25156# 0.02606f
C5626 a_23780_1636# VPWR 0.20968f
C5627 a_61412_12612# a_61500_12568# 0.28563f
C5628 a_51644_12568# a_51532_12135# 0.02634f
C5629 _398_.C _474_.Q 0.05617f
C5630 _448_.Q a_44162_24120# 0.01085f
C5631 a_6723_30644# a_7180_30951# 0.00916f
C5632 a_47636_23588# VPWR 0.00833f
C5633 _474_.CLK vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN 0.01154f
C5634 _304_.B a_52660_21640# 0.00196f
C5635 a_33524_24776# a_33376_23659# 0.00179f
C5636 vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN 0.02209f
C5637 a_64412_15271# a_64324_15368# 0.28563f
C5638 a_48956_11000# a_49404_11000# 0.01288f
C5639 a_42372_1636# a_42820_1636# 0.01328f
C5640 a_65332_12232# a_65444_11044# 0.02666f
C5641 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I 0.01626f
C5642 a_35988_18504# VPWR 0.20595f
C5643 _334_.A1 a_35292_26247# 0.00143f
C5644 a_40020_16936# a_40468_16936# 0.01328f
C5645 _270_.A2 _272_.A2 0.40625f
C5646 _447_.Q a_43819_24372# 0.00999f
C5647 a_66204_15704# a_66340_15368# 0.00168f
C5648 a_22560_30288# uio_out[4] 0.29344f
C5649 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN 0.02033f
C5650 a_2724_26724# a_2364_26680# 0.08717f
C5651 a_4516_26724# a_4964_26724# 0.01328f
C5652 _474_.CLK a_48104_30219# 0.03733f
C5653 _243_.B2 a_58588_26247# 0.00264f
C5654 _260_.A1 _325_.B 0.00298f
C5655 a_29788_30345# a_30132_29977# 0.00275f
C5656 _303_.ZN _328_.A2 0.06888f
C5657 a_18096_27165# a_19612_26247# 0.00467f
C5658 a_30724_26020# a_31844_26344# 0.006f
C5659 a_1828_20452# VPWR 0.20348f
C5660 a_19076_31048# uio_out[5] 0.00444f
C5661 _450_.D _332_.Z 0.00201f
C5662 a_49316_12612# VPWR 0.21035f
C5663 a_61276_2727# VPWR 0.33981f
C5664 a_4604_28248# a_4516_26724# 0.0027f
C5665 a_66988_18407# a_66900_18504# 0.28563f
C5666 a_4828_2727# a_4964_1636# 0.00154f
C5667 a_4740_2824# a_5188_2824# 0.01328f
C5668 a_16500_26344# a_16948_26344# 0.01328f
C5669 a_5300_20072# VPWR 0.21406f
C5670 a_57580_17272# a_58028_17272# 0.01255f
C5671 a_2364_29383# a_2724_29480# 0.08717f
C5672 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN a_61500_17272# 0.00677f
C5673 a_4964_15748# a_4940_15271# 0.00172f
C5674 a_62060_10567# VPWR 0.31547f
C5675 _460_.Q a_35652_26344# 0.00332f
C5676 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN 0.0071f
C5677 _459_.CLK a_30476_25112# 0.00323f
C5678 a_40668_15271# a_41028_15368# 0.08717f
C5679 a_4940_21543# a_4964_20452# 0.0016f
C5680 _412_.B2 a_51540_24776# 0.00386f
C5681 a_60516_26344# vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I 0.02911f
C5682 a_24004_23208# VPWR 0.20622f
C5683 _424_.A2 _402_.ZN 0.03811f
C5684 a_38971_18559# a_39216_18191# 0.00232f
C5685 _272_.B1 _258_.ZN 0.00449f
C5686 a_51620_19911# a_52024_20083# 0.41635f
C5687 a_26160_27165# VPWR 0.52906f
C5688 _397_.A1 a_46837_29076# 0.00987f
C5689 a_4156_28248# a_4604_28248# 0.01222f
C5690 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN clk 0.01187f
C5691 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN 0.04127f
C5692 a_54780_2727# a_55140_2824# 0.08717f
C5693 _330_.A1 a_41776_20072# 0.01262f
C5694 a_38876_19975# a_38788_20072# 0.28563f
C5695 a_20620_23544# a_20532_22020# 0.00151f
C5696 _244_.Z clk 0.00253f
C5697 _300_.ZN a_38576_22504# 0.07542f
C5698 a_32068_16936# a_32068_15748# 0.05841f
C5699 _260_.A2 a_42161_24776# 0.01746f
C5700 a_50772_18504# a_51220_18504# 0.01328f
C5701 a_14796_25112# a_15244_25112# 0.01288f
C5702 a_23892_23588# a_23980_23544# 0.28563f
C5703 a_18740_25156# a_18828_25112# 0.28563f
C5704 a_3620_1256# VPWR 0.22197f
C5705 a_4068_31048# VPWR 0.22189f
C5706 _246_.B2 a_60916_29612# 0.00139f
C5707 a_51084_13703# a_50996_13800# 0.28563f
C5708 a_51240_23340# a_51668_23340# 0.00223f
C5709 a_30476_20408# a_30924_20408# 0.0131f
C5710 a_32628_20452# a_32268_20408# 0.08717f
C5711 a_24196_31048# a_24652_30951# 0.0065f
C5712 a_19372_30345# uio_out[5] 0.04792f
C5713 a_60964_27912# _245_.Z 0.00308f
C5714 _243_.ZN VPWR 0.42906f
C5715 a_37868_16839# a_37780_16936# 0.28563f
C5716 a_54420_21976# VPWR 0.37255f
C5717 a_61836_16839# VPWR 0.33064f
C5718 _478_.D a_54356_24776# 0.00298f
C5719 a_29916_1592# VPWR 0.29679f
C5720 _417_.Z a_49672_19668# 0.00757f
C5721 a_19188_23588# a_19164_23111# 0.00172f
C5722 a_1020_12135# a_1468_12135# 0.0131f
C5723 a_58588_12568# a_58476_12135# 0.02634f
C5724 a_15244_23544# a_15244_23111# 0.05841f
C5725 _447_.Q a_36860_23111# 0.06066f
C5726 a_5412_1636# a_5860_1636# 0.01328f
C5727 a_1828_1636# a_1916_1592# 0.28563f
C5728 _473_.Q a_49448_20936# 0.00255f
C5729 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_57492_23588# 0.00164f
C5730 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_62796_25640# 0.00492f
C5731 _371_.A1 _371_.A3 0.61285f
C5732 a_52660_21640# VPWR 0.00636f
C5733 a_2812_11000# a_2812_10567# 0.05841f
C5734 a_56260_11044# a_55900_11000# 0.08707f
C5735 a_33508_31048# uo_out[4] 0.00112f
C5736 a_58836_12232# a_58924_10567# 0.00151f
C5737 a_16240_26795# a_17120_27209# 0.00306f
C5738 a_60405_31198# ui_in[3] 0.00102f
C5739 a_18096_27165# _455_.D 0.00158f
C5740 a_20308_26724# a_20396_26680# 0.28563f
C5741 a_59652_25640# a_60064_25156# 0.00736f
C5742 a_44688_26399# VPWR 0.00204f
C5743 a_46044_1159# a_46716_1159# 0.00544f
C5744 a_35204_2824# a_35068_1592# 0.00154f
C5745 a_39012_2824# a_39012_1636# 0.05841f
C5746 _448_.Q _302_.Z 1.20473f
C5747 a_63876_18884# a_64324_18884# 0.01328f
C5748 _336_.A2 a_26756_24801# 0.0051f
C5749 a_20844_20408# VPWR 0.31143f
C5750 a_41476_26344# a_41564_24679# 0.0014f
C5751 _397_.A2 a_48596_28292# 0.00676f
C5752 a_61860_30736# ui_in[2] 0.57278f
C5753 a_1380_15748# a_1020_15704# 0.08717f
C5754 a_3172_15748# a_3620_15748# 0.01328f
C5755 a_55452_12568# VPWR 0.31389f
C5756 _355_.C a_24636_25641# 0.00545f
C5757 a_11772_2727# a_11908_1636# 0.00154f
C5758 _452_.Q _439_.ZN 0.15586f
C5759 a_64748_23111# vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN 0.00102f
C5760 a_50212_15368# a_50660_15368# 0.01328f
C5761 _229_.I _250_.ZN 0.4771f
C5762 a_13788_29383# a_13700_29480# 0.28563f
C5763 a_19164_30951# uio_out[5] 0.01273f
C5764 _360_.ZN a_33164_24679# 0.00142f
C5765 _395_.A2 _398_.C 0.3975f
C5766 a_1916_8999# a_2276_9096# 0.08717f
C5767 a_55924_10664# VPWR 0.20614f
C5768 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_65756_26247# 0.001f
C5769 a_52092_15271# a_52004_15368# 0.28563f
C5770 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN 0.06829f
C5771 a_55228_27815# a_55588_27912# 0.08674f
C5772 a_2812_7431# a_3172_7528# 0.08717f
C5773 a_3708_5863# a_4068_5960# 0.08717f
C5774 a_4940_4295# a_5300_4392# 0.08674f
C5775 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I a_65668_27912# 0.00436f
C5776 _371_.A1 uo_out[7] 0.08272f
C5777 _474_.Q a_47636_18884# 0.00184f
C5778 a_53660_15271# a_54108_15271# 0.0131f
C5779 a_4068_15368# VPWR 0.22146f
C5780 _334_.A1 _437_.A1 0.0038f
C5781 _255_.ZN a_57220_29861# 0.13181f
C5782 _398_.C a_46984_23588# 0.02081f
C5783 _436_.ZN a_40357_24776# 0.08453f
C5784 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I a_62084_18884# 0.00731f
C5785 a_66204_2727# a_66116_2824# 0.28563f
C5786 a_17036_21976# a_17484_21976# 0.01288f
C5787 a_20980_22020# a_21068_21976# 0.28563f
C5788 a_32604_15271# VPWR 0.29679f
C5789 a_58140_26680# VPWR 0.3532f
C5790 a_50436_30689# _268_.A2 0.19678f
C5791 a_24428_23544# a_24340_22020# 0.00151f
C5792 a_35180_16839# a_35628_16839# 0.01288f
C5793 a_39124_16936# a_39012_15748# 0.02666f
C5794 a_65220_17316# VPWR 0.20921f
C5795 _251_.A1 a_60084_25640# 0.00558f
C5796 a_31396_23208# a_31484_21543# 0.00151f
C5797 a_29848_29535# VPWR 0.00204f
C5798 a_2364_7431# VPWR 0.30029f
C5799 a_26020_1256# VPWR 0.20772f
C5800 a_30836_23588# a_31284_23588# 0.01328f
C5801 a_47076_1256# a_47524_1256# 0.01328f
C5802 a_24080_25227# a_25643_25273# 0.41635f
C5803 a_4156_4295# VPWR 0.3269f
C5804 a_26108_2727# a_26556_2727# 0.0131f
C5805 a_47524_13800# a_47972_13800# 0.01328f
C5806 a_64860_26247# VPWR 0.34004f
C5807 a_16700_29383# VPWR 0.29679f
C5808 a_61612_13703# a_61972_13800# 0.08707f
C5809 a_8627_30644# VPWR 0.18927f
C5810 a_48396_16839# a_48756_16936# 0.08707f
C5811 a_20003_29611# uio_out[5] 0.552f
C5812 a_51892_10664# a_51868_9432# 0.0016f
C5813 a_19612_23111# a_19636_22020# 0.0016f
C5814 a_22352_25987# a_23332_26344# 0.00702f
C5815 a_41364_16936# VPWR 0.20986f
C5816 a_43716_1636# VPWR 0.20348f
C5817 a_7516_1159# a_7428_1256# 0.28563f
C5818 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I a_64860_19975# 0.00473f
C5819 a_55452_12568# a_55476_12232# 0.00172f
C5820 a_20172_25112# a_20060_24679# 0.02634f
C5821 _268_.A2 _272_.B1 0.13692f
C5822 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN a_55788_25112# 0.00613f
C5823 a_3260_29816# a_3708_29816# 0.01288f
C5824 a_7204_29860# a_7292_29816# 0.28563f
C5825 _436_.B _436_.ZN 0.0999f
C5826 _258_.ZN VPWR 0.69766f
C5827 a_33412_17316# a_33860_17316# 0.01328f
C5828 _351_.A2 VPWR 0.39735f
C5829 a_62756_11044# a_63204_11044# 0.01328f
C5830 a_63068_15271# a_63204_14180# 0.00154f
C5831 a_24900_1636# a_24764_1159# 0.00168f
C5832 a_48508_1592# a_48956_1592# 0.01288f
C5833 a_52452_1636# a_52540_1592# 0.28563f
C5834 a_6084_2824# VPWR 0.20815f
C5835 a_58924_17272# VPWR 0.33773f
C5836 _452_.CLK a_34160_20523# 0.07321f
C5837 a_32964_20072# a_32964_18884# 0.05841f
C5838 a_4940_23111# a_5388_23111# 0.01222f
C5839 a_29680_26724# VPWR 0.01466f
C5840 a_41572_18504# VPWR 0.00713f
C5841 a_19035_28409# a_18400_28733# 0.02112f
C5842 _373_.A2 a_28928_29123# 0.00129f
C5843 a_52204_18407# a_52564_18504# 0.08717f
C5844 a_45956_2824# a_45956_1636# 0.05841f
C5845 a_42148_2824# a_42012_1592# 0.00154f
C5846 a_53908_18504# a_53996_16839# 0.0027f
C5847 a_52116_18504# VPWR 0.20595f
C5848 a_16140_25112# VPWR 0.29679f
C5849 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I a_62620_19975# 0.00473f
C5850 a_35740_30951# uo_out[2] 0.00207f
C5851 a_48529_22460# _473_.Q 0.51759f
C5852 a_25652_31048# VPWR 0.36065f
C5853 a_31820_20408# VPWR 0.31594f
C5854 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN 0.00109f
C5855 _397_.A1 _395_.A1 0.11321f
C5856 a_31172_15748# a_30812_15704# 0.08707f
C5857 a_2364_12135# VPWR 0.30029f
C5858 a_39996_15704# a_40132_15368# 0.00168f
C5859 _336_.Z a_28891_25273# 0.01085f
C5860 a_26916_2824# a_27588_2824# 0.00347f
C5861 _450_.D a_43452_18191# 0.21205f
C5862 a_28054_30196# uio_out[0] 0.00531f
C5863 _304_.B _268_.A2 0.02974f
C5864 _397_.A4 a_47297_25596# 0.02996f
C5865 a_20672_30301# a_22188_29383# 0.00467f
C5866 a_19948_27815# uio_out[7] 0.00127f
C5867 _340_.ZN _454_.Q 0.00484f
C5868 _343_.A2 a_24392_28248# 0.5288f
C5869 _270_.A2 _228_.ZN 0.25335f
C5870 _324_.C _470_.D 0.06347f
C5871 a_19524_21640# a_19412_20452# 0.02666f
C5872 a_39772_20408# a_39772_19975# 0.05841f
C5873 a_4516_15748# VPWR 0.20862f
C5874 _274_.A1 a_56484_29480# 0.0236f
C5875 a_51556_15368# VPWR 0.20348f
C5876 _352_.A2 a_25928_25273# 0.00112f
C5877 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN a_55452_15271# 0.00171f
C5878 _251_.A1 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN 0.02636f
C5879 a_49988_21236# a_50212_20452# 0.00102f
C5880 a_62560_25112# VPWR 0.52839f
C5881 a_24340_22020# a_23980_21976# 0.08707f
C5882 a_55004_15271# VPWR 0.32938f
C5883 a_35740_17272# a_35652_15748# 0.00151f
C5884 _304_.B a_43008_26795# 0.01513f
C5885 a_47972_14180# a_48420_14180# 0.01328f
C5886 _452_.CLK a_36996_17316# 0.01602f
C5887 a_36524_16839# VPWR 0.31389f
C5888 a_25100_30951# a_25012_31048# 0.28563f
C5889 _252_.B _242_.Z 0.00509f
C5890 _474_.CLK a_54468_21640# 0.00741f
C5891 a_48420_1256# VPWR 0.20348f
C5892 a_62396_14136# a_62308_12612# 0.00151f
C5893 a_47636_25940# clkbuf_1_0__f_clk.I 0.00295f
C5894 a_34756_17316# VPWR 0.23214f
C5895 _424_.A1 a_54692_20452# 0.00112f
C5896 a_26720_30301# VPWR 0.57659f
C5897 a_26556_23111# a_26580_22020# 0.0016f
C5898 a_18492_1159# a_18852_1256# 0.08717f
C5899 a_59172_26724# _251_.ZN 0.002f
C5900 _384_.A3 _476_.Q 0.1007f
C5901 a_49852_1592# VPWR 0.30447f
C5902 _447_.Q a_38764_20408# 0.00977f
C5903 a_11684_29480# a_12356_29480# 0.00347f
C5904 a_62508_12135# a_62956_12135# 0.01288f
C5905 a_48508_12135# a_49204_12232# 0.01227f
C5906 a_15492_1636# a_15580_1592# 0.28563f
C5907 a_11548_1592# a_11996_1592# 0.01288f
C5908 _474_.CLK a_52228_19368# 0.03059f
C5909 a_61860_27912# a_61748_26724# 0.02666f
C5910 a_32268_23544# a_32380_23111# 0.02634f
C5911 a_10564_29860# a_10204_29816# 0.08707f
C5912 _358_.A3 a_30240_24776# 0.00145f
C5913 a_48868_31048# a_49316_31048# 0.01328f
C5914 a_56260_15368# a_56260_14180# 0.05841f
C5915 a_56348_11000# a_56460_10567# 0.02634f
C5916 a_60292_11044# a_60268_10567# 0.00172f
C5917 a_28484_2824# VPWR 0.20348f
C5918 _251_.A1 _255_.I 0.05246f
C5919 a_55228_1592# a_55900_1592# 0.00544f
C5920 a_3708_23111# a_3620_23208# 0.28563f
C5921 _459_.CLK a_20396_27815# 0.00158f
C5922 a_24988_24679# a_25436_24679# 0.01288f
C5923 a_16588_24679# a_16500_24776# 0.28563f
C5924 a_18400_28733# uio_out[7] 0.04109f
C5925 a_55140_15748# a_55228_15704# 0.28563f
C5926 a_3620_9096# a_4068_9096# 0.01328f
C5927 _437_.A1 _448_.Q 0.05142f
C5928 a_33052_19975# a_33500_19975# 0.0131f
C5929 a_4940_7431# a_4964_6340# 0.0016f
C5930 a_4852_7528# a_5300_7528# 0.01328f
C5931 a_64324_5960# a_64772_5960# 0.01328f
C5932 a_65220_4392# a_65668_4392# 0.01328f
C5933 _294_.A2 _359_.B 0.83325f
C5934 a_49316_14180# VPWR 0.21389f
C5935 a_34732_18407# a_35180_18407# 0.01255f
C5936 a_3708_18407# a_4068_18504# 0.08717f
C5937 a_26020_31048# a_25792_30301# 0.00186f
C5938 _351_.ZN a_25300_26344# 0.00866f
C5939 a_13252_29480# VPWR 0.20348f
C5940 a_37532_15704# a_37980_15704# 0.012f
C5941 a_63852_12135# VPWR 0.31547f
C5942 _268_.A2 VPWR 1.40185f
C5943 _334_.A1 a_37844_29860# 0.00311f
C5944 _358_.A3 a_36548_26344# 0.00178f
C5945 a_52676_15748# a_52540_15271# 0.00168f
C5946 a_48732_15704# a_48732_15271# 0.05841f
C5947 a_27172_24328# VPWR 0.51923f
C5948 _424_.A2 a_46068_25156# 0.00209f
C5949 _251_.A1 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN 0.00461f
C5950 a_64772_7528# VPWR 0.20727f
C5951 a_66564_4392# VPWR 0.20631f
C5952 _438_.A2 _301_.A1 0.07835f
C5953 a_39012_15748# VPWR 0.20676f
C5954 _241_.I0 a_56404_27208# 0.11424f
C5955 a_56124_28248# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.0017f
C5956 a_30836_22020# a_31284_22020# 0.01328f
C5957 a_53548_18407# a_53996_18407# 0.01222f
C5958 uio_in[4] uio_in[3] 0.01021f
C5959 _398_.C _427_.A2 0.13771f
C5960 a_43008_26795# VPWR 1.10464f
C5961 a_46156_25112# clkbuf_1_0__f_clk.I 0.0021f
C5962 _474_.D a_50748_20408# 0.0426f
C5963 a_54892_18407# VPWR 0.31795f
C5964 a_25420_30345# a_25764_29977# 0.00275f
C5965 _294_.A2 a_36656_29123# 0.00266f
C5966 _373_.A2 uio_out[0] 0.01078f
C5967 _424_.B1 clkload0.Z 0.00258f
C5968 a_5500_1592# a_5636_1256# 0.00168f
C5969 a_48508_2727# a_48956_2727# 0.0131f
C5970 a_27884_25641# VPWR 0.39762f
C5971 a_49404_18407# a_49540_17316# 0.00154f
C5972 a_1828_12612# a_2276_12612# 0.01328f
C5973 _459_.CLK a_18028_28777# 0.00442f
C5974 a_47388_17272# a_47500_16839# 0.02634f
C5975 a_51332_17316# a_51308_16839# 0.00172f
C5976 _417_.A2 _384_.A1 0.11729f
C5977 a_46852_17316# VPWR 0.20885f
C5978 a_25348_23208# a_25236_22020# 0.02666f
C5979 a_63652_1636# VPWR 0.22423f
C5980 a_29916_1159# a_29828_1256# 0.28563f
C5981 a_59820_12135# a_59732_12232# 0.28563f
C5982 a_18852_1636# a_18492_1592# 0.08707f
C5983 _475_.Q a_49988_21236# 0.00912f
C5984 _474_.CLK a_53908_18504# 0.00373f
C5985 a_16028_29816# a_16700_29816# 0.00544f
C5986 a_17060_29860# a_17508_29860# 0.01328f
C5987 a_19612_21543# VPWR 0.32678f
C5988 a_27228_26247# a_27140_26344# 0.28563f
C5989 a_45260_17272# a_45708_17272# 0.01255f
C5990 a_49740_10567# a_50188_10567# 0.01288f
C5991 a_62172_1592# a_62620_1592# 0.01288f
C5992 a_67236_11044# a_67212_10567# 0.00172f
C5993 a_50884_2824# VPWR 0.21449f
C5994 _452_.Q _303_.ZN 1.97258f
C5995 a_2276_23208# a_2724_23208# 0.01328f
C5996 a_23644_23111# a_24004_23208# 0.08707f
C5997 a_50076_9432# VPWR 0.32111f
C5998 a_17932_21543# a_18716_21543# 0.00443f
C5999 a_19972_2824# a_20060_1159# 0.0027f
C6000 _325_.A1 _324_.B 0.29135f
C6001 a_56348_14136# VPWR 0.31423f
C6002 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.0373f
C6003 _294_.A2 a_32144_26724# 0.00898f
C6004 a_57940_12232# VPWR 0.21723f
C6005 a_44836_15748# a_44476_15704# 0.08707f
C6006 a_3708_29816# a_3708_29383# 0.05841f
C6007 a_7652_29860# a_7516_29383# 0.00168f
C6008 a_49316_2824# a_49764_2824# 0.01328f
C6009 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I a_57132_18407# 0.02997f
C6010 _419_.Z a_52452_21236# 0.00552f
C6011 a_40132_20452# a_40220_20408# 0.28563f
C6012 a_32096_24419# VPWR 0.52133f
C6013 a_62868_23208# vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I 0.00364f
C6014 a_51956_26183# _412_.ZN 0.03083f
C6015 a_63428_20072# VPWR 0.20348f
C6016 a_9980_2727# a_9892_2824# 0.28563f
C6017 a_52676_15748# VPWR 0.20622f
C6018 a_55004_21543# a_55452_21543# 0.012f
C6019 a_50884_9476# a_50524_9432# 0.08717f
C6020 _258_.I vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.00159f
C6021 a_26020_31048# a_26468_31048# 0.01328f
C6022 a_25100_30951# uio_out[2] 0.04244f
C6023 a_55004_14136# a_55452_14136# 0.0131f
C6024 a_59284_14180# a_59372_14136# 0.28563f
C6025 a_61636_15368# a_61612_13703# 0.00131f
C6026 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I 0.02706f
C6027 _447_.Q a_36996_21640# 0.01811f
C6028 a_22560_30288# a_22548_29480# 0.00117f
C6029 _437_.A1 a_37532_26680# 0.01573f
C6030 a_60180_13800# a_60292_12612# 0.02666f
C6031 a_56372_13800# a_56348_12568# 0.0016f
C6032 _350_.A1 _350_.A2 2.18194f
C6033 a_59172_23208# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.00169f
C6034 _402_.A1 a_50120_26476# 0.00294f
C6035 _287_.A2 a_31031_27208# 0.00115f
C6036 a_38752_26344# VPWR 0.01426f
C6037 a_13788_1159# VPWR 0.29679f
C6038 a_19164_24679# a_19188_23588# 0.0016f
C6039 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_62284_23544# 0.00945f
C6040 a_40892_1159# a_41252_1256# 0.08717f
C6041 a_3620_24776# a_3620_23588# 0.05841f
C6042 a_32292_23208# a_32180_22020# 0.02666f
C6043 a_56372_12232# a_57044_12232# 0.00347f
C6044 _460_.D a_33148_25641# 0.2143f
C6045 a_24304_26795# a_24692_27209# 0.00393f
C6046 a_25348_1636# a_25796_1636# 0.01328f
C6047 _294_.ZN a_32132_27912# 0.00431f
C6048 a_16500_21640# VPWR 0.20348f
C6049 a_21052_26031# a_21516_25112# 0.00104f
C6050 a_52676_17316# a_52316_17272# 0.08707f
C6051 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN a_59260_21976# 0.00614f
C6052 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_59172_22020# 0.00193f
C6053 a_42996_18840# a_43392_19369# 0.00232f
C6054 a_65668_27912# VPWR 0.23462f
C6055 a_46716_10567# a_46628_10664# 0.28563f
C6056 _260_.A1 _441_.A2 0.05282f
C6057 _454_.Q a_23627_27967# 0.00174f
C6058 _442_.ZN _441_.ZN 0.08951f
C6059 _251_.ZN a_59397_26344# 0.04515f
C6060 a_54692_18884# a_54780_18840# 0.28563f
C6061 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN a_54332_18840# 0.00225f
C6062 a_30240_24776# a_31803_24831# 0.41635f
C6063 a_31168_24419# a_30796_24463# 0.10745f
C6064 _452_.CLK a_37084_25112# 0.00111f
C6065 _324_.B _327_.A2 0.01272f
C6066 a_63764_23588# clk 0.00127f
C6067 a_61052_9432# VPWR 0.31143f
C6068 a_5052_23544# VPWR 0.33516f
C6069 a_5052_6296# VPWR 0.33516f
C6070 a_25420_30345# uio_out[2] 0.00121f
C6071 a_4156_13703# VPWR 0.3269f
C6072 a_16588_21543# a_16948_21640# 0.08717f
C6073 a_65668_3204# VPWR 0.21209f
C6074 a_62084_20072# a_62532_20072# 0.01328f
C6075 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_56836_27208# 0.00141f
C6076 _255_.I a_58020_27508# 0.00103f
C6077 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I a_67684_24776# 0.04846f
C6078 _424_.A2 a_49068_20408# 0.00519f
C6079 _355_.C a_30836_23588# 0.00236f
C6080 _419_.A4 a_47776_20893# 0.04258f
C6081 _452_.CLK a_36060_19369# 0.02774f
C6082 _427_.ZN a_54020_21640# 0.01058f
C6083 a_47076_11044# VPWR 0.20348f
C6084 a_31124_25156# VPWR 0.0142f
C6085 a_47748_15748# a_47836_15704# 0.28563f
C6086 a_51332_15748# a_51780_15748# 0.01328f
C6087 a_39996_2727# a_40132_1636# 0.00154f
C6088 a_67436_19975# a_67796_20072# 0.08663f
C6089 _459_.Q _371_.A1 0.0719f
C6090 a_17036_26247# VPWR 0.2974f
C6091 a_33948_18840# VPWR 0.30233f
C6092 a_20956_2727# a_21316_2824# 0.08717f
C6093 a_49404_30951# _392_.A2 0.00208f
C6094 _311_.A2 a_39178_23208# 0.00461f
C6095 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN 0.00747f
C6096 VPWR uo_out[2] 0.75918f
C6097 _452_.Q a_40356_15748# 0.00186f
C6098 _304_.B _282_.ZN 0.00103f
C6099 a_2812_9432# a_2812_8999# 0.05841f
C6100 _436_.B a_40780_27815# 0.03773f
C6101 a_63204_14180# a_63292_14136# 0.28563f
C6102 a_28908_21976# a_28820_20452# 0.00151f
C6103 a_52540_14136# a_52428_13703# 0.02634f
C6104 a_15604_20452# a_16052_20452# 0.01328f
C6105 _474_.Q a_50748_20408# 0.03092f
C6106 _430_.ZN a_39332_23588# 0.00102f
C6107 _327_.Z a_41188_18840# 0.19063f
C6108 _247_.ZN a_59572_29076# 0.49455f
C6109 _337_.A3 a_26750_28776# 0.00228f
C6110 _455_.Q _371_.A2 2.42126f
C6111 a_67124_13800# a_67236_12612# 0.02666f
C6112 a_50748_12568# a_51196_12568# 0.01288f
C6113 _267_.A2 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 1.48185f
C6114 _424_.A1 a_52452_21236# 0.04585f
C6115 a_43232_29480# a_43003_28409# 0.00173f
C6116 _480_.Q a_43296_28733# 0.20236f
C6117 a_21316_24776# a_21428_23588# 0.02666f
C6118 _284_.ZN a_42368_28733# 0.01919f
C6119 a_52316_1159# a_52228_1256# 0.28563f
C6120 a_36188_1159# VPWR 0.3289f
C6121 a_46628_31048# a_45416_29885# 0.00187f
C6122 a_45956_31048# a_45904_30180# 0.00255f
C6123 a_36996_26344# a_37444_26344# 0.01328f
C6124 a_43828_29860# _480_.Q 0.00376f
C6125 vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I a_67996_21976# 0.00474f
C6126 _427_.B1 a_52452_24072# 0.26809f
C6127 a_65644_23544# VPWR 0.32804f
C6128 a_3620_10664# a_4068_10664# 0.01328f
C6129 a_12444_1159# a_12892_1159# 0.0131f
C6130 a_57580_10567# a_57940_10664# 0.08707f
C6131 _250_.B a_62503_28293# 0.09756f
C6132 _381_.A2 a_48560_26369# 0.01688f
C6133 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I 0.00559f
C6134 a_52512_19715# VPWR 0.39698f
C6135 _459_.Q a_30476_25112# 0.00971f
C6136 a_37179_24831# a_37464_24831# 0.00277f
C6137 a_15156_22020# VPWR 0.20348f
C6138 a_33188_23208# a_33636_23208# 0.01328f
C6139 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN 0.00229f
C6140 _245_.Z vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I 0.00291f
C6141 a_27924_23588# VPWR 0.20348f
C6142 a_15156_21640# a_15604_21640# 0.01328f
C6143 _467_.D a_16588_28248# 0.05186f
C6144 a_65868_13703# VPWR 0.34719f
C6145 a_16252_2727# VPWR 0.31605f
C6146 a_3172_18884# a_3260_18840# 0.28563f
C6147 a_42148_2824# a_42236_1159# 0.0027f
C6148 a_51428_23340# VPWR 0.00646f
C6149 a_27900_21543# a_27812_21640# 0.28563f
C6150 _399_.A1 a_50732_23233# 0.00436f
C6151 a_1380_29860# VPWR 0.20348f
C6152 a_60604_26247# vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I 0.00354f
C6153 a_38336_18147# a_37964_18191# 0.10745f
C6154 a_43916_29816# VPWR 0.32359f
C6155 a_53212_11000# VPWR 0.31898f
C6156 _441_.A3 _438_.ZN 0.02891f
C6157 _251_.A1 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.23728f
C6158 a_62620_15704# a_63068_15704# 0.0131f
C6159 a_66116_15748# a_65756_15704# 0.0869f
C6160 _448_.D a_36612_20072# 0.00621f
C6161 a_14796_27815# VPWR 0.30073f
C6162 _330_.A1 _400_.ZN 0.04527f
C6163 _257_.B _247_.ZN 0.0542f
C6164 a_43008_26795# a_44744_26355# 0.00569f
C6165 a_64748_23111# a_65756_23111# 0.00323f
C6166 a_32380_2727# a_32292_2824# 0.28563f
C6167 _457_.D a_25643_25273# 0.01957f
C6168 _282_.ZN VPWR 0.62603f
C6169 a_3708_23544# a_4156_23544# 0.0131f
C6170 a_13252_1256# a_13700_1256# 0.01328f
C6171 a_63204_9476# a_63652_9476# 0.01328f
C6172 a_61860_9476# a_61500_9432# 0.08717f
C6173 a_3708_6296# a_4156_6296# 0.0131f
C6174 _325_.A2 _450_.D 0.02778f
C6175 a_2812_7864# a_3260_7864# 0.0131f
C6176 a_19076_31048# _465_.D 0.01202f
C6177 a_4604_4728# a_5052_4728# 0.01222f
C6178 a_2812_13703# a_3260_13703# 0.0131f
C6179 a_64324_3204# a_64772_3204# 0.01328f
C6180 a_27676_26680# a_28124_26680# 0.012f
C6181 _247_.B _244_.Z 0.3956f
C6182 a_60268_14136# a_60268_13703# 0.05841f
C6183 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I 0.00689f
C6184 a_21204_20452# a_21292_20408# 0.28563f
C6185 a_10004_31048# a_9980_29383# 0.00134f
C6186 a_3708_29383# a_4156_29383# 0.0131f
C6187 a_4828_30951# a_4740_31048# 0.28563f
C6188 a_51791_30644# vgaringosc.ro_inv1.inv_array_notouch_\[1\].I 0.13041f
C6189 _270_.A2 ui_in[3] 0.02834f
C6190 a_9668_1636# VPWR 0.20854f
C6191 _459_.CLK a_20172_25112# 0.00383f
C6192 a_60628_13800# a_60716_12135# 0.0027f
C6193 a_58052_12612# a_57692_12568# 0.08707f
C6194 _478_.D a_54444_23544# 0.00828f
C6195 _455_.Q a_22996_25156# 0.00436f
C6196 _388_.B a_43356_30951# 0.01769f
C6197 a_67124_20452# VPWR 0.20904f
C6198 a_43892_20072# a_43668_19668# 0.01751f
C6199 a_58588_1159# VPWR 0.30504f
C6200 a_45732_11044# a_46180_11044# 0.01328f
C6201 _350_.A1 _334_.A1 0.1107f
C6202 a_63292_1159# a_63652_1256# 0.08717f
C6203 a_35428_1636# a_35516_1592# 0.28563f
C6204 a_39012_1636# a_39460_1636# 0.01328f
C6205 a_3620_16936# a_4068_16936# 0.01328f
C6206 _474_.CLK a_54356_20072# 0.05291f
C6207 a_67100_18840# VPWR 0.31547f
C6208 _416_.A3 a_46848_20893# 0.0647f
C6209 a_36100_25156# a_35740_25112# 0.0869f
C6210 _258_.I a_56596_29861# 0.07391f
C6211 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN a_62196_23588# 0.00613f
C6212 a_42148_27912# a_42596_27912# 0.01328f
C6213 a_932_10664# a_932_9476# 0.05841f
C6214 _441_.ZN _435_.ZN 0.08581f
C6215 _402_.A1 _404_.A1 0.14072f
C6216 _437_.A1 a_36172_24463# 0.00105f
C6217 a_59932_1592# a_59932_1159# 0.05841f
C6218 a_49764_26724# _284_.A2 0.01292f
C6219 _436_.ZN _433_.ZN 0.43707f
C6220 a_33860_18504# a_33860_17316# 0.05841f
C6221 a_20868_2824# a_20732_1592# 0.00154f
C6222 _230_.I _229_.I 2.31632f
C6223 a_28820_22020# VPWR 0.20684f
C6224 a_36300_23544# VPWR 0.31438f
C6225 a_59732_13800# VPWR 0.20595f
C6226 _465_.D a_19372_30345# 0.23387f
C6227 a_32604_18840# a_33052_18840# 0.0131f
C6228 a_38428_2727# VPWR 0.33981f
C6229 a_15692_26247# a_16140_26247# 0.0131f
C6230 a_1468_26247# a_1828_26344# 0.08717f
C6231 a_59708_23111# vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I 0.00311f
C6232 _352_.A2 _336_.A1 0.16601f
C6233 _252_.B a_60156_27815# 0.01148f
C6234 _474_.CLK a_47802_26724# 0.00384f
C6235 a_15044_29860# VPWR 0.2085f
C6236 a_64436_16936# a_64324_15748# 0.02666f
C6237 _260_.A2 _441_.A2 0.02011f
C6238 a_67324_11000# VPWR 0.31589f
C6239 _287_.A1 uo_out[6] 1.54368f
C6240 a_4156_15271# a_4852_15368# 0.01227f
C6241 _451_.Q a_38764_20408# 0.00195f
C6242 a_25884_23111# VPWR 0.34806f
C6243 a_64748_23544# a_64748_23111# 0.05841f
C6244 _424_.B1 a_50120_26476# 0.00817f
C6245 _452_.CLK _444_.D 0.04066f
C6246 _459_.CLK _349_.A4 0.26454f
C6247 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN 0.00135f
C6248 a_33932_24073# a_34276_23705# 0.00275f
C6249 _237_.A1 _243_.B2 0.00148f
C6250 a_64660_23208# a_65668_23208# 0.00196f
C6251 _325_.ZN a_44459_18559# 0.00966f
C6252 _294_.A2 a_35710_28776# 0.00166f
C6253 a_43356_2727# a_43716_2824# 0.08717f
C6254 a_28000_29480# a_28388_29167# 0.00393f
C6255 _452_.CLK a_34939_23705# 0.03767f
C6256 _284_.B _447_.Q 0.01737f
C6257 a_65420_16839# a_65332_16936# 0.28563f
C6258 _437_.A1 _234_.ZN 0.03514f
C6259 _480_.Q a_44028_27815# 0.00539f
C6260 a_63516_18407# a_63964_18407# 0.0131f
C6261 a_20084_23588# a_19724_23544# 0.08707f
C6262 a_4964_25156# a_4604_25112# 0.08674f
C6263 a_2364_25112# a_2812_25112# 0.0131f
C6264 _284_.ZN a_43132_27815# 0.01309f
C6265 _459_.CLK a_30388_28776# 0.0257f
C6266 a_26580_20452# a_27028_20452# 0.01328f
C6267 _268_.A2 a_49112_29885# 0.06071f
C6268 a_49316_31048# a_49496_30345# 0.00192f
C6269 _359_.B a_40644_29480# 0.00199f
C6270 _459_.Q a_34700_28776# 0.00153f
C6271 _350_.A1 a_35652_31048# 0.01443f
C6272 _424_.B2 a_52512_19715# 0.00207f
C6273 a_19164_30951# _465_.D 0.00519f
C6274 a_1468_16839# a_1380_16936# 0.28563f
C6275 a_59484_11000# a_59396_9476# 0.00151f
C6276 _397_.A1 _389_.ZN 0.05599f
C6277 a_23332_1636# VPWR 0.20874f
C6278 a_61412_12612# a_61052_12568# 0.08707f
C6279 _448_.Q a_43750_23544# 0.07664f
C6280 a_64548_12612# a_64996_12612# 0.01328f
C6281 a_47412_23588# VPWR 0.00754f
C6282 _474_.CLK a_55340_19975# 0.02996f
C6283 a_25124_28776# a_28364_28776# 0.00576f
C6284 _260_.A1 a_40580_20452# 0.0027f
C6285 _459_.CLK _467_.D 0.31471f
C6286 _241_.I0 VPWR 0.96838f
C6287 a_63964_15271# a_64324_15368# 0.08717f
C6288 a_52452_11044# a_53124_11044# 0.00347f
C6289 a_61524_12232# a_61500_11000# 0.0016f
C6290 a_10564_1636# a_10428_1159# 0.00168f
C6291 a_35540_18504# VPWR 0.20605f
C6292 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN 0.00937f
C6293 vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN a_61724_18407# 0.00647f
C6294 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.79599f
C6295 a_2276_26724# a_2364_26680# 0.28563f
C6296 a_20672_30301# uio_out[4] 0.02732f
C6297 a_61300_16936# a_61300_15748# 0.05841f
C6298 _346_.B a_20756_26724# 0.03622f
C6299 _474_.CLK a_45904_30180# 0.00124f
C6300 a_65332_10664# a_65780_10664# 0.01328f
C6301 a_34620_1159# a_35292_1159# 0.00544f
C6302 _287_.A1 uo_out[5] 1.5124f
C6303 a_18096_27165# a_19164_26247# 0.03096f
C6304 a_16240_26795# a_16588_26247# 0.0074f
C6305 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I 0.00157f
C6306 vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I 0.71012f
C6307 a_1380_20452# VPWR 0.20348f
C6308 a_18628_31048# uio_out[5] 0.00152f
C6309 a_48868_12612# VPWR 0.21134f
C6310 a_60828_2727# VPWR 0.31143f
C6311 a_35728_29480# a_36608_29167# 0.00306f
C6312 _465_.D a_20003_29611# 0.00173f
C6313 a_66540_18407# a_66900_18504# 0.0869f
C6314 a_4852_20072# VPWR 0.22733f
C6315 a_38788_15368# a_39236_15368# 0.01328f
C6316 a_2364_29383# a_2276_29480# 0.28563f
C6317 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I 0.07983f
C6318 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I a_61300_16936# 0.07118f
C6319 _355_.C a_19372_30345# 0.01092f
C6320 a_64300_23544# a_64748_23544# 0.01255f
C6321 a_2364_15704# a_2364_15271# 0.05841f
C6322 _460_.Q a_35204_26344# 0.04682f
C6323 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.0068f
C6324 _459_.CLK a_30388_25156# 0.0015f
C6325 a_61612_10567# VPWR 0.31547f
C6326 a_40668_15271# a_40580_15368# 0.28563f
C6327 a_23556_23208# VPWR 0.20622f
C6328 a_63068_17272# a_63092_16936# 0.00172f
C6329 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN VPWR 1.01842f
C6330 a_35616_24776# a_36004_24463# 0.00393f
C6331 a_46198_27060# _402_.ZN 0.0013f
C6332 a_42236_15271# a_42684_15271# 0.0131f
C6333 a_24860_27209# VPWR 0.39942f
C6334 _452_.CLK a_34715_22137# 0.00111f
C6335 _270_.A2 _267_.A2 0.01448f
C6336 a_4604_21976# a_5052_21976# 0.01222f
C6337 a_54780_2727# a_54692_2824# 0.28563f
C6338 a_66204_17272# a_66652_17272# 0.01255f
C6339 a_26580_23588# a_27028_23588# 0.01328f
C6340 a_20420_23208# a_20508_21543# 0.00151f
C6341 a_23892_23588# a_23532_23544# 0.08717f
C6342 a_3172_1256# VPWR 0.20993f
C6343 _246_.B2 a_60656_29612# 0.00518f
C6344 a_35652_1256# a_36100_1256# 0.01328f
C6345 _402_.ZN clkbuf_1_0__f_clk.I 0.14393f
C6346 a_3620_31048# VPWR 0.22347f
C6347 a_18740_25156# a_18380_25112# 0.08707f
C6348 _436_.ZN _261_.ZN 0.15621f
C6349 a_50636_13703# a_50996_13800# 0.08707f
C6350 a_64300_13703# a_64972_13703# 0.00544f
C6351 a_32180_20452# a_32268_20408# 0.28563f
C6352 a_51240_23340# a_51428_23340# 0.00843f
C6353 a_14684_2727# a_15132_2727# 0.0131f
C6354 a_28054_30196# a_28000_29480# 0.00725f
C6355 vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I 0.1629f
C6356 a_58228_27912# VPWR 0.00904f
C6357 a_60516_27912# _245_.Z 0.00135f
C6358 a_37420_16839# a_37780_16936# 0.08707f
C6359 a_31396_26724# _358_.A3 0.00117f
C6360 a_19744_30301# uio_out[5] 0.04134f
C6361 a_54668_10567# a_54692_9476# 0.0016f
C6362 a_49828_22020# VPWR 0.00718f
C6363 a_29468_1592# VPWR 0.29679f
C6364 a_40668_1592# a_40804_1256# 0.00168f
C6365 _478_.D a_53908_24776# 0.00162f
C6366 a_61388_16839# VPWR 0.31552f
C6367 a_1828_1636# a_1468_1592# 0.08707f
C6368 a_29716_31048# _287_.A2 0.00268f
C6369 a_3708_25112# a_3708_24679# 0.05841f
C6370 a_60516_27912# a_60604_26247# 0.0027f
C6371 _417_.A2 _416_.A3 1.0808f
C6372 a_1828_17316# a_2276_17316# 0.01328f
C6373 a_67772_21543# VPWR 0.34683f
C6374 _284_.ZN _260_.A2 0.01006f
C6375 a_50772_16936# a_51220_16936# 0.01328f
C6376 a_45148_1592# a_45596_1592# 0.01288f
C6377 a_55812_11044# a_55900_11000# 0.28563f
C6378 a_59396_11044# a_59844_11044# 0.01328f
C6379 a_4964_11044# a_4940_10567# 0.00172f
C6380 _381_.Z _281_.ZN 0.04884f
C6381 a_16240_26795# a_16628_27209# 0.00393f
C6382 a_20308_26724# a_19948_26680# 0.08674f
C6383 a_17168_27165# a_16796_27209# 0.10745f
C6384 _433_.ZN _439_.ZN 0.06307f
C6385 _402_.A1 a_48384_26724# 0.02267f
C6386 a_4852_27912# a_4964_26724# 0.02666f
C6387 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_64300_23544# 0.00124f
C6388 _474_.Q a_51220_22504# 0.00164f
C6389 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN 0.68671f
C6390 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I a_57580_18840# 0.00712f
C6391 _249_.A2 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.00415f
C6392 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN 0.06071f
C6393 a_53348_18884# VPWR 0.14741f
C6394 a_20396_20408# VPWR 0.31143f
C6395 a_4156_27815# a_4940_27815# 0.00443f
C6396 _336_.A2 a_25796_24776# 0.00133f
C6397 a_60909_30600# ui_in[2] 0.04301f
C6398 _346_.B _378_.I 0.489f
C6399 _375_.Z a_21652_29480# 0.0013f
C6400 _397_.A2 a_47924_28292# 0.00333f
C6401 _355_.C a_25008_25597# 0.00315f
C6402 a_55004_12568# VPWR 0.31389f
C6403 _281_.ZN a_51540_24776# 0.00104f
C6404 a_932_15748# a_1020_15704# 0.28563f
C6405 a_15492_2824# a_16164_2824# 0.00347f
C6406 a_13340_29383# a_13700_29480# 0.08717f
C6407 VPWR uio_oe[6] 0.34414f
C6408 _355_.C a_20003_29611# 0.08688f
C6409 a_19035_28409# a_19500_27815# 0.02338f
C6410 a_55476_10664# VPWR 0.20614f
C6411 a_57580_18407# a_57492_18504# 0.28563f
C6412 a_1916_8999# a_1828_9096# 0.28563f
C6413 a_55228_27815# a_55140_27912# 0.28563f
C6414 a_2812_7431# a_2724_7528# 0.28563f
C6415 a_41488_24072# a_42796_23981# 0.0146f
C6416 _242_.Z _243_.B2 0.17666f
C6417 a_3708_5863# a_3620_5960# 0.28563f
C6418 a_51644_15271# a_52004_15368# 0.08717f
C6419 a_3172_21640# a_3172_20452# 0.05841f
C6420 a_39536_26795# _442_.ZN 0.24818f
C6421 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.02341f
C6422 a_60212_25156# a_61836_25515# 0.00523f
C6423 a_4940_4295# a_4852_4392# 0.28563f
C6424 a_30388_28776# uo_out[7] 0.07276f
C6425 a_3620_15368# VPWR 0.22347f
C6426 _355_.C a_26916_27912# 0.00203f
C6427 a_20980_22020# a_20620_21976# 0.08707f
C6428 a_65756_2727# a_66116_2824# 0.0869f
C6429 a_32156_15271# VPWR 0.29679f
C6430 a_1828_14180# a_2276_14180# 0.01328f
C6431 a_64772_17316# VPWR 0.20727f
C6432 a_28900_29535# VPWR 0.00246f
C6433 a_24080_25227# a_25936_25597# 0.02307f
C6434 a_25008_25597# a_24636_25641# 0.10745f
C6435 a_25572_1256# VPWR 0.20627f
C6436 a_1916_7431# VPWR 0.297f
C6437 a_3708_4295# VPWR 0.33374f
C6438 a_58028_17272# vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN 0.00332f
C6439 _437_.A1 a_39256_28292# 0.12988f
C6440 a_61612_13703# a_61524_13800# 0.28563f
C6441 a_16252_29383# VPWR 0.33444f
C6442 a_51084_28248# a_51048_26680# 0.00115f
C6443 a_7628_30951# VPWR 0.33205f
C6444 a_48396_16839# a_48308_16936# 0.28563f
C6445 a_18760_29032# uio_out[5] 0.01303f
C6446 _352_.ZN a_27228_26247# 0.01025f
C6447 a_40916_16936# VPWR 0.2076f
C6448 a_43268_1636# VPWR 0.20511f
C6449 a_51532_12135# a_51980_12135# 0.01288f
C6450 a_7068_1159# a_7428_1256# 0.08717f
C6451 a_65532_12568# a_65420_12135# 0.02634f
C6452 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN a_55340_25112# 0.00149f
C6453 a_22636_23544# a_22748_23111# 0.02634f
C6454 a_8188_1592# a_8772_1636# 0.01675f
C6455 a_7204_29860# a_6844_29816# 0.08707f
C6456 a_56572_29383# VPWR 0.32598f
C6457 _336_.Z a_28012_24679# 0.00506f
C6458 _317_.A2 a_34396_21543# 0.00136f
C6459 a_24900_27912# VPWR 0.60579f
C6460 a_5636_2824# VPWR 0.20815f
C6461 a_49404_11000# a_49292_10567# 0.02634f
C6462 a_52452_1636# a_52092_1592# 0.08707f
C6463 a_58476_17272# VPWR 0.3434f
C6464 _300_.ZN _438_.ZN 0.04869f
C6465 _416_.A1 a_46820_20569# 0.00132f
C6466 _242_.Z a_59172_26724# 0.00121f
C6467 a_28596_26725# VPWR 0.64228f
C6468 a_4940_24679# a_5388_24679# 0.01222f
C6469 _386_.ZN _404_.A1 0.13952f
C6470 _373_.A2 a_28000_29480# 0.00695f
C6471 a_57020_1159# a_57468_1159# 0.0131f
C6472 a_52204_18407# a_52116_18504# 0.28563f
C6473 a_51668_18504# VPWR 0.20595f
C6474 a_65756_18840# a_66204_18840# 0.01255f
C6475 a_15692_25112# VPWR 0.29679f
C6476 a_31372_20408# VPWR 0.31594f
C6477 a_20396_27815# a_20308_27912# 0.28563f
C6478 a_25100_30951# VPWR 0.32115f
C6479 _358_.A3 VPWR 1.83942f
C6480 a_34308_15748# a_34756_15748# 0.01328f
C6481 a_30724_15748# a_30812_15704# 0.28563f
C6482 a_1916_12135# VPWR 0.297f
C6483 _336_.Z a_29184_25597# 0.02001f
C6484 _319_.ZN _319_.A2 0.0988f
C6485 _450_.D a_43824_18147# 0.00516f
C6486 a_19500_27815# uio_out[7] 0.00294f
C6487 a_20672_30301# a_21740_29383# 0.03096f
C6488 _301_.A1 a_38228_20452# 0.00895f
C6489 a_27900_21543# a_27924_20452# 0.0016f
C6490 _324_.C a_44961_27912# 0.00368f
C6491 a_4068_15748# VPWR 0.2157f
C6492 a_51108_15368# VPWR 0.20353f
C6493 _402_.A1 _435_.A3 0.05902f
C6494 _419_.A4 a_48292_26369# 0.00137f
C6495 a_23892_22020# a_23980_21976# 0.28563f
C6496 _268_.A1 a_52756_29076# 0.33361f
C6497 a_27476_22020# a_27924_22020# 0.01328f
C6498 a_61836_25515# VPWR 0.61964f
C6499 a_54556_15271# VPWR 0.32938f
C6500 a_45708_16839# a_46156_16839# 0.01288f
C6501 a_36076_16839# VPWR 0.31389f
C6502 _474_.CLK a_54020_21640# 0.00555f
C6503 a_45060_31048# a_45088_29123# 0.00105f
C6504 a_40580_26344# _264_.B 0.00363f
C6505 a_24652_30951# a_25012_31048# 0.08674f
C6506 a_47972_1256# VPWR 0.20348f
C6507 a_58052_1256# a_58500_1256# 0.01328f
C6508 a_58388_13800# a_58836_13800# 0.01328f
C6509 a_4852_13800# a_4964_12612# 0.02666f
C6510 a_37084_2727# a_37532_2727# 0.0131f
C6511 _261_.ZN _439_.ZN 0.07004f
C6512 _358_.A2 _459_.D 0.13137f
C6513 _424_.A1 a_54244_20452# 0.00264f
C6514 a_25420_30345# VPWR 0.40008f
C6515 a_34308_17316# VPWR 0.21526f
C6516 _447_.Q a_38316_20408# 0.00983f
C6517 a_18492_1159# a_18404_1256# 0.28563f
C6518 a_49404_1592# VPWR 0.30187f
C6519 a_48508_12135# a_48420_12232# 0.28563f
C6520 a_15492_1636# a_15132_1592# 0.08707f
C6521 a_62396_12568# a_62420_12232# 0.00172f
C6522 _304_.B _324_.B 1.51427f
C6523 a_10116_29860# a_10204_29816# 0.28563f
C6524 a_13700_29860# a_14148_29860# 0.01328f
C6525 a_36188_17272# a_36636_17272# 0.01288f
C6526 _334_.A1 _290_.ZN 0.24568f
C6527 a_49628_17272# a_49652_16936# 0.00172f
C6528 a_65980_11000# a_66428_11000# 0.01288f
C6529 a_43736_25896# _448_.Q 0.00105f
C6530 a_58948_1636# a_59396_1636# 0.01328f
C6531 a_28036_2824# VPWR 0.20348f
C6532 _459_.CLK a_19948_27815# 0.00103f
C6533 _324_.C _480_.Q 0.09388f
C6534 a_24540_23111# a_24988_23111# 0.01288f
C6535 _350_.A1 _370_.ZN 0.07971f
C6536 a_3260_23111# a_3620_23208# 0.08717f
C6537 a_16140_24679# a_16500_24776# 0.08717f
C6538 a_55140_15748# a_54780_15704# 0.08663f
C6539 a_48868_14180# VPWR 0.21224f
C6540 a_8548_2824# a_8636_1159# 0.0027f
C6541 a_3708_18407# a_3620_18504# 0.28563f
C6542 a_36188_26680# a_36188_26247# 0.05841f
C6543 a_1380_31048# a_1380_29860# 0.05841f
C6544 a_33376_23659# a_34256_24073# 0.00306f
C6545 _351_.ZN a_24228_26344# 0.00447f
C6546 a_12804_29480# VPWR 0.20348f
C6547 a_63404_12135# VPWR 0.31547f
C6548 _336_.A2 _352_.ZN 0.33256f
C6549 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I 0.00652f
C6550 a_37892_2824# a_38340_2824# 0.01328f
C6551 a_25660_2727# a_25796_1636# 0.00154f
C6552 _416_.A1 a_44340_26183# 0.04682f
C6553 a_49764_31048# VPWR 0.21575f
C6554 _334_.A1 a_37396_29860# 0.00158f
C6555 _290_.ZN a_35156_29860# 0.00135f
C6556 _358_.A3 a_36100_26344# 0.00414f
C6557 a_25884_24679# VPWR 0.35314f
C6558 a_64324_7528# VPWR 0.22383f
C6559 a_26468_21640# a_26580_20452# 0.02666f
C6560 a_66116_4392# VPWR 0.23643f
C6561 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.00454f
C6562 a_5052_3160# a_5188_2824# 0.00168f
C6563 a_38564_15748# VPWR 0.22726f
C6564 a_55676_28248# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.00158f
C6565 _268_.A2 a_58116_30344# 0.00423f
C6566 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN a_54892_16839# 0.00404f
C6567 _398_.C a_51332_24072# 0.0078f
C6568 a_50748_14136# a_51196_14136# 0.01288f
C6569 a_54444_18407# VPWR 0.31547f
C6570 a_64324_15368# a_64188_14136# 0.00154f
C6571 _474_.D a_50300_20408# 0.02834f
C6572 _343_.A2 a_23920_27555# 0.0178f
C6573 _294_.A2 a_35728_29480# 0.0719f
C6574 a_28672_31048# uio_out[0] 0.00181f
C6575 _424_.B1 a_48384_26724# 0.00674f
C6576 a_28256_25597# VPWR 0.18826f
C6577 _324_.C _246_.B2 0.10926f
C6578 a_34292_28776# uo_out[7] 0.00118f
C6579 a_44252_30951# uio_in[5] 0.00117f
C6580 _290_.ZN a_35652_31048# 0.0014f
C6581 _409_.ZN _390_.ZN 0.02571f
C6582 _459_.CLK a_18400_28733# 0.00276f
C6583 a_66228_10664# a_66204_9432# 0.0016f
C6584 a_46404_17316# VPWR 0.23079f
C6585 a_63068_1592# VPWR 0.35728f
C6586 a_29468_1159# a_29828_1256# 0.08717f
C6587 a_30924_23544# a_30948_23208# 0.00172f
C6588 a_18404_1636# a_18492_1592# 0.28563f
C6589 a_21988_1636# a_22436_1636# 0.01328f
C6590 a_56796_12568# a_56708_11044# 0.0027f
C6591 a_59372_12135# a_59732_12232# 0.08707f
C6592 a_45284_12232# a_45732_12232# 0.01328f
C6593 _324_.B VPWR 4.1551f
C6594 a_56148_23588# a_56124_23111# 0.00172f
C6595 _287_.A1 _460_.Q 0.06649f
C6596 _474_.CLK a_53460_18504# 0.00546f
C6597 a_19164_21543# VPWR 0.33846f
C6598 a_19164_26247# a_19188_25156# 0.0016f
C6599 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_62956_23111# 0.03454f
C6600 _474_.Q a_49404_18407# 0.00251f
C6601 a_63292_11000# a_63404_10567# 0.02634f
C6602 a_53212_11000# a_53236_10664# 0.00172f
C6603 a_50436_2824# VPWR 0.27305f
C6604 _324_.C _281_.ZN 0.86966f
C6605 a_23644_23111# a_23556_23208# 0.28563f
C6606 _404_.A1 a_47476_28292# 0.00127f
C6607 a_18628_24776# a_19076_24776# 0.01328f
C6608 a_55228_28248# a_55676_28248# 0.01222f
C6609 a_49628_9432# VPWR 0.31767f
C6610 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I VPWR 0.73599f
C6611 _451_.Q _284_.B 0.0959f
C6612 a_59844_2824# a_59844_1636# 0.05841f
C6613 a_56036_2824# a_55900_1592# 0.00154f
C6614 _452_.Q _452_.D 0.00345f
C6615 a_26916_31048# VPWR 0.22322f
C6616 a_55900_14136# VPWR 0.31389f
C6617 _474_.CLK _397_.A4 0.05192f
C6618 a_33860_18504# a_34644_18504# 0.00276f
C6619 a_55956_25940# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.05394f
C6620 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_56516_26344# 0.62304f
C6621 _452_.CLK a_34844_24679# 0.04684f
C6622 a_40444_15704# a_40892_15704# 0.01288f
C6623 a_44388_15748# a_44476_15704# 0.28563f
C6624 a_57492_12232# VPWR 0.21191f
C6625 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I a_65196_23544# 0.00304f
C6626 ui_in[7] ui_in[6] 0.01143f
C6627 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I a_56684_18407# 0.00681f
C6628 a_40132_20452# a_39772_20408# 0.08674f
C6629 _248_.B1 a_65668_27912# 0.00221f
C6630 a_31803_24831# VPWR 0.37274f
C6631 a_49496_30345# _409_.ZN 0.00787f
C6632 a_62980_20072# VPWR 0.20348f
C6633 a_9532_2727# a_9892_2824# 0.08717f
C6634 a_52228_15748# VPWR 0.20622f
C6635 a_61724_19975# a_62172_19975# 0.0131f
C6636 hold2.Z a_43126_24119# 0.00896f
C6637 _386_.A4 _404_.A1 0.13621f
C6638 a_46716_30951# _393_.ZN 0.00111f
C6639 a_50436_9476# a_50524_9432# 0.28563f
C6640 _461_.D a_32352_29535# 0.00242f
C6641 a_24652_30951# uio_out[2] 0.00531f
C6642 a_59284_14180# a_58924_14136# 0.0869f
C6643 _379_.Z _378_.ZN 0.01654f
C6644 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_65668_27912# 0.0206f
C6645 _447_.Q a_36548_21640# 0.09439f
C6646 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN VPWR 0.69986f
C6647 _336_.Z a_28372_23588# 0.0013f
C6648 _437_.A1 a_37084_26680# 0.0012f
C6649 _384_.ZN clkbuf_1_0__f_clk.I 0.14968f
C6650 _388_.B _397_.A2 0.10316f
C6651 a_47524_12612# a_47972_12612# 0.01328f
C6652 a_59484_2727# a_59932_2727# 0.0131f
C6653 a_37892_26344# VPWR 0.2115f
C6654 a_30948_23208# a_30924_21976# 0.0016f
C6655 _252_.ZN a_60940_28248# 0.01168f
C6656 a_40892_1159# a_40804_1256# 0.28563f
C6657 _460_.D a_33520_25597# 0.00851f
C6658 a_13340_1159# VPWR 0.29679f
C6659 a_3172_20072# a_3620_20072# 0.01328f
C6660 a_2724_12232# a_2724_11044# 0.05841f
C6661 a_932_4772# a_1020_4728# 0.28563f
C6662 a_64772_4392# a_64772_3204# 0.05841f
C6663 a_16052_21640# VPWR 0.20348f
C6664 _251_.A1 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN 0.40347f
C6665 _241_.I0 a_57156_27912# 0.03783f
C6666 hold2.Z a_43192_25640# 0.00108f
C6667 a_52228_17316# a_52316_17272# 0.28563f
C6668 a_48284_17272# a_48732_17272# 0.01288f
C6669 a_46268_10567# a_46628_10664# 0.08717f
C6670 a_60268_10567# a_60716_10567# 0.01288f
C6671 _340_.A2 _349_.A4 0.45414f
C6672 a_1020_1159# a_1468_1159# 0.0131f
C6673 a_45596_1592# a_45596_1159# 0.05841f
C6674 a_6532_2824# a_6396_1592# 0.00154f
C6675 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN VPWR 0.84569f
C6676 a_22212_23208# a_22660_23208# 0.01328f
C6677 a_54692_18884# a_54332_18840# 0.08674f
C6678 a_57940_18884# a_58388_18884# 0.01328f
C6679 _452_.CLK a_36636_25112# 0.00272f
C6680 a_30240_24776# a_30796_24463# 0.8399f
C6681 a_60604_9432# VPWR 0.31605f
C6682 _316_.ZN _317_.A2 0.10339f
C6683 a_63316_23588# clk 0.00148f
C6684 a_28796_21543# a_29244_21543# 0.01288f
C6685 a_4604_6296# VPWR 0.33016f
C6686 a_16588_21543# a_16500_21640# 0.28563f
C6687 a_4604_23544# VPWR 0.33016f
C6688 a_65220_3204# VPWR 0.20921f
C6689 a_3708_13703# VPWR 0.33374f
C6690 _404_.A1 _407_.A1 0.00305f
C6691 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN 0.0075f
C6692 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN 0.03675f
C6693 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_55340_26680# 0.09282f
C6694 _355_.C a_30388_23588# 0.00249f
C6695 _256_.A2 clk 0.02956f
C6696 _452_.CLK a_36432_19325# 0.02445f
C6697 _427_.ZN a_53572_21640# 0.01058f
C6698 a_17284_31048# a_17148_29816# 0.00154f
C6699 a_47748_15748# a_47388_15704# 0.08707f
C6700 a_46628_11044# VPWR 0.20348f
C6701 a_60292_2824# a_60740_2824# 0.01328f
C6702 a_67436_19975# a_67348_20072# 0.28563f
C6703 a_10540_30951# a_10564_29860# 0.0016f
C6704 _459_.Q a_30388_28776# 0.01163f
C6705 a_67861_30644# ena 0.00145f
C6706 a_33500_18840# VPWR 0.30042f
C6707 a_16588_26247# VPWR 0.31848f
C6708 a_20956_2727# a_20868_2824# 0.28563f
C6709 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN 0.01887f
C6710 _261_.ZN _303_.ZN 0.00684f
C6711 a_48956_30951# _392_.A2 0.00208f
C6712 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN 0.80566f
C6713 a_4964_9476# a_4940_8999# 0.00172f
C6714 a_55676_9432# a_56124_9432# 0.0131f
C6715 a_1828_1256# a_2276_1256# 0.01328f
C6716 a_2276_31048# a_2724_31048# 0.01328f
C6717 a_66340_14180# a_66788_14180# 0.01328f
C6718 a_63204_14180# a_62844_14136# 0.08707f
C6719 _336_.Z a_29268_22020# 0.00263f
C6720 _474_.Q a_50300_20408# 0.02088f
C6721 _327_.Z a_40684_19368# 0.00105f
C6722 _459_.CLK a_25124_28776# 0.03204f
C6723 a_49652_13800# a_49740_12135# 0.00151f
C6724 a_63316_13800# a_63292_12568# 0.0016f
C6725 _474_.CLK a_52756_29076# 0.00536f
C6726 _313_.ZN a_36772_23208# 0.11088f
C6727 a_43232_29480# a_43296_28733# 0.00781f
C6728 _255_.ZN vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I 0.0311f
C6729 a_58063_30644# _272_.A2 0.00283f
C6730 a_35740_1159# VPWR 0.3289f
C6731 a_51868_1159# a_52228_1256# 0.08717f
C6732 a_28124_1592# a_28572_1592# 0.01288f
C6733 a_57020_23111# vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.00111f
C6734 a_67124_12232# a_67572_12232# 0.01328f
C6735 a_50996_12232# a_51108_11044# 0.02666f
C6736 _345_.A2 _346_.A2 0.63307f
C6737 a_65196_23544# VPWR 0.33397f
C6738 a_57580_10567# a_57492_10664# 0.28563f
C6739 a_34448_25597# a_34844_24679# 0.00201f
C6740 _424_.B1 _419_.Z 0.04041f
C6741 _250_.B a_62279_28293# 0.0286f
C6742 _381_.A2 a_48292_26369# 0.0229f
C6743 _424_.ZN a_53380_20127# 0.00159f
C6744 a_52024_20083# VPWR 1.09802f
C6745 a_14708_22020# VPWR 0.22176f
C6746 a_45396_28292# _404_.A1 0.00414f
C6747 _256_.A2 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I 0.04285f
C6748 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.02977f
C6749 _459_.Q a_30388_25156# 0.0159f
C6750 _245_.Z a_59652_25640# 0.00158f
C6751 _352_.A2 a_29244_23111# 0.00118f
C6752 _246_.B2 _252_.ZN 0.56161f
C6753 a_3172_18884# a_2812_18840# 0.08717f
C6754 _424_.B1 _399_.A2 0.00717f
C6755 a_27476_23588# VPWR 0.21464f
C6756 a_27452_21543# a_27812_21640# 0.08707f
C6757 _397_.A4 _398_.C 0.03824f
C6758 a_50732_23233# VPWR 0.01343f
C6759 a_15580_2727# VPWR 0.33981f
C6760 a_65420_13703# VPWR 0.32215f
C6761 _467_.D a_16140_28248# 0.01305f
C6762 _399_.A1 a_50420_23233# 0.02533f
C6763 a_932_29860# VPWR 0.22176f
C6764 a_54244_15748# a_54692_15748# 0.01328f
C6765 a_60292_11044# VPWR 0.21241f
C6766 _275_.A2 _409_.ZN 0.00826f
C6767 _251_.A1 a_56404_27208# 0.83439f
C6768 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN 0.00785f
C6769 a_5388_27815# VPWR 0.35574f
C6770 a_65668_15748# a_65756_15704# 0.28563f
C6771 a_37444_26344# a_37444_25156# 0.05841f
C6772 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I 0.63026f
C6773 a_31932_2727# a_32292_2824# 0.08717f
C6774 _457_.D a_25936_25597# 0.03607f
C6775 a_26468_31048# uio_out[2] 0.00296f
C6776 a_61748_23588# a_62196_23588# 0.01328f
C6777 a_47724_18840# a_48172_18840# 0.01222f
C6778 a_48888_19243# a_49896_18909# 0.02307f
C6779 a_4964_7908# a_5052_7864# 0.28563f
C6780 _437_.A1 a_39760_23588# 0.0122f
C6781 a_61412_9476# a_61500_9432# 0.28563f
C6782 _365_.ZN a_35008_27533# 0.02696f
C6783 a_21204_20452# a_20844_20408# 0.08717f
C6784 a_58028_18840# a_57940_17316# 0.0027f
C6785 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN 0.00115f
C6786 a_19052_20408# a_19500_20408# 0.0131f
C6787 a_4156_30951# a_4740_31048# 0.01675f
C6788 a_9220_1636# VPWR 0.2085f
C6789 a_26332_1592# a_26468_1256# 0.00168f
C6790 _459_.CLK a_19724_25112# 0.00182f
C6791 a_53660_12568# a_54108_12568# 0.01288f
C6792 a_57604_12612# a_57692_12568# 0.28563f
C6793 _281_.ZN _281_.A1 0.4796f
C6794 _388_.B a_42908_30951# 0.01934f
C6795 a_24900_24776# a_24876_23544# 0.0016f
C6796 _325_.A2 a_43916_16839# 0.03577f
C6797 _304_.B a_56124_28248# 0.00221f
C6798 a_63292_1159# a_63204_1256# 0.28563f
C6799 _274_.ZN _274_.A3 0.21666f
C6800 a_8860_29816# a_8996_29480# 0.00168f
C6801 a_34644_18504# a_34732_16839# 0.00151f
C6802 a_58140_1159# VPWR 0.33803f
C6803 a_66676_20452# VPWR 0.20851f
C6804 a_35652_25156# a_35740_25112# 0.28563f
C6805 a_57940_12232# a_58052_11044# 0.02666f
C6806 a_54132_12232# a_54108_11000# 0.0016f
C6807 _416_.ZN a_46128_20127# 0.00159f
C6808 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I 0.00108f
C6809 a_66652_18840# VPWR 0.31547f
C6810 _416_.A3 a_45920_20523# 0.07686f
C6811 a_35428_1636# a_35068_1592# 0.08707f
C6812 _398_.C a_51956_26183# 0.04515f
C6813 _452_.CLK _439_.ZN 0.00363f
C6814 _474_.Q _421_.B 0.26217f
C6815 a_49764_26724# a_51048_26680# 0.01082f
C6816 a_54132_10664# a_54580_10664# 0.01328f
C6817 a_23196_1159# a_23868_1159# 0.00544f
C6818 _395_.A1 _384_.A1 0.00513f
C6819 _272_.A2 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I 0.00169f
C6820 a_61412_17316# a_61388_16839# 0.00172f
C6821 a_28372_22020# VPWR 0.20622f
C6822 a_66787_30600# _256_.A2 0.26056f
C6823 _358_.A3 _360_.ZN 0.58159f
C6824 _355_.C a_21287_29076# 0.00105f
C6825 a_25796_21640# a_26468_21640# 0.00347f
C6826 a_37980_2727# VPWR 0.31143f
C6827 a_59284_13800# VPWR 0.20595f
C6828 a_53124_2824# a_53212_1159# 0.0027f
C6829 _465_.D a_19744_30301# 0.02149f
C6830 a_1468_26247# a_1380_26344# 0.28563f
C6831 a_2276_15368# a_2724_15368# 0.01328f
C6832 _267_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.40275f
C6833 a_14596_29860# VPWR 0.2085f
C6834 a_66876_11000# VPWR 0.31589f
C6835 a_4156_15271# a_4068_15368# 0.28563f
C6836 _393_.A3 _397_.A4 0.0106f
C6837 _470_.Q _470_.D 0.00693f
C6838 a_25436_23111# VPWR 0.31768f
C6839 a_30812_15271# a_31260_15271# 0.0131f
C6840 _424_.B1 _424_.A1 0.2167f
C6841 _325_.ZN a_43452_18191# 0.03282f
C6842 a_67548_17272# a_67460_15748# 0.00151f
C6843 a_43356_2727# a_43268_2824# 0.28563f
C6844 a_54892_26680# a_55340_26680# 0.01255f
C6845 _452_.CLK a_35232_24029# 0.0496f
C6846 a_28556_29167# a_28900_29535# 0.00275f
C6847 a_63428_17316# a_63876_17316# 0.01328f
C6848 a_64972_16839# a_65332_16936# 0.08674f
C6849 _437_.A1 a_40038_28720# 0.01484f
C6850 _480_.Q a_43580_27815# 0.00131f
C6851 a_66652_9432# a_67100_9432# 0.0131f
C6852 a_19636_23588# a_19724_23544# 0.28563f
C6853 a_15692_23544# a_16140_23544# 0.01288f
C6854 a_24228_1256# a_24676_1256# 0.01328f
C6855 a_1468_5863# a_1916_5863# 0.0131f
C6856 _284_.ZN a_42684_27815# 0.0048f
C6857 a_64860_6296# a_64860_5863# 0.05841f
C6858 a_4516_25156# a_4604_25112# 0.28563f
C6859 a_67324_14136# a_67212_13703# 0.02634f
C6860 a_2364_4295# a_2812_4295# 0.0131f
C6861 a_65756_4728# a_65756_4295# 0.05841f
C6862 a_53324_13703# a_53772_13703# 0.01288f
C6863 a_3260_2727# a_3708_2727# 0.0131f
C6864 a_35540_16936# a_35516_15271# 0.00134f
C6865 a_19164_30951# a_19076_31048# 0.28563f
C6866 a_14684_29383# a_15132_29383# 0.0131f
C6867 _218_.ZN _419_.Z 0.02634f
C6868 _424_.B2 a_52024_20083# 0.07114f
C6869 _452_.CLK _330_.ZN 0.15155f
C6870 _350_.A1 a_35204_31048# 0.01443f
C6871 a_1020_16839# a_1380_16936# 0.08717f
C6872 _403_.ZN VPWR 0.42658f
C6873 _355_.C a_27228_26680# 0.00318f
C6874 a_18816_29931# a_19696_30345# 0.00306f
C6875 a_22884_1636# VPWR 0.2085f
C6876 a_51196_12568# a_51084_12135# 0.02634f
C6877 a_6172_30951# a_6723_30644# 0.03643f
C6878 _448_.Q a_43126_24119# 0.0023f
C6879 _384_.A3 _474_.Q 2.223f
C6880 a_60964_12612# a_61052_12568# 0.28563f
C6881 _474_.CLK a_54892_19975# 0.02923f
C6882 _325_.B a_42392_19243# 0.05438f
C6883 a_47172_23588# VPWR 0.00677f
C6884 _399_.A2 _218_.ZN 0.01229f
C6885 a_25124_28776# a_27868_28776# 0.00582f
C6886 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN VPWR 0.80065f
C6887 _459_.CLK a_17060_29480# 0.04864f
C6888 _251_.A1 _238_.I 0.07857f
C6889 a_56124_28248# VPWR 0.3101f
C6890 a_63964_15271# a_63876_15368# 0.28563f
C6891 a_52452_11044# a_52540_11000# 0.28563f
C6892 a_64884_12232# a_64996_11044# 0.02666f
C6893 a_48508_11000# a_48956_11000# 0.01288f
C6894 a_39572_16936# a_40020_16936# 0.01328f
C6895 a_41924_1636# a_42372_1636# 0.01328f
C6896 a_35092_18504# VPWR 0.2323f
C6897 _476_.Q _424_.ZN 0.00722f
C6898 a_65756_15704# a_65892_15368# 0.00168f
C6899 a_58476_20408# vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.0105f
C6900 VPWR uo_out[1] 0.79394f
C6901 a_2276_26724# a_1916_26680# 0.08717f
C6902 a_4068_26724# a_4516_26724# 0.01328f
C6903 a_20379_29977# uio_out[4] 0.00244f
C6904 _474_.CLK a_45416_29885# 0.0059f
C6905 a_1020_1159# a_932_1256# 0.28563f
C6906 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN clk 0.04366f
C6907 a_18096_27165# a_18716_26247# 0.02396f
C6908 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN 0.00156f
C6909 a_932_20452# VPWR 0.22176f
C6910 a_60380_2727# VPWR 0.31143f
C6911 a_48420_12612# VPWR 0.20348f
C6912 _465_.D a_18760_29032# 0.00133f
C6913 _402_.A1 _411_.A2 1.35182f
C6914 a_66540_18407# a_66452_18504# 0.28563f
C6915 a_4068_2824# a_4740_2824# 0.00347f
C6916 a_49764_26724# _381_.A2 0.00122f
C6917 a_16052_26344# a_16500_26344# 0.01328f
C6918 a_1916_29383# a_2276_29480# 0.08717f
C6919 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.00222f
C6920 a_4068_20072# VPWR 0.22146f
C6921 _260_.ZN _324_.B 0.08516f
C6922 a_57132_17272# a_57580_17272# 0.01255f
C6923 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I 0.00748f
C6924 _355_.C a_19744_30301# 0.03493f
C6925 a_58063_30644# _228_.ZN 0.00345f
C6926 _460_.Q a_34308_26344# 0.14134f
C6927 _416_.A1 a_40092_27209# 0.00167f
C6928 a_61164_10567# VPWR 0.31547f
C6929 a_40220_15271# a_40580_15368# 0.08717f
C6930 a_29804_21976# a_29692_21543# 0.02634f
C6931 a_58836_18884# VPWR 0.20893f
C6932 a_23108_23208# VPWR 0.20622f
C6933 _284_.A2 a_43736_25896# 0.05983f
C6934 _274_.ZN _324_.C 0.00104f
C6935 a_25232_27165# VPWR 0.1886f
C6936 a_3708_28248# a_4156_28248# 0.0131f
C6937 a_54332_2727# a_54692_2824# 0.08717f
C6938 _260_.A2 a_39985_24372# 0.00512f
C6939 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I 0.0996f
C6940 a_20172_23544# a_20084_22020# 0.00151f
C6941 a_31620_16936# a_31620_15748# 0.05841f
C6942 a_50324_18504# a_50772_18504# 0.01328f
C6943 a_23444_23588# a_23532_23544# 0.28563f
C6944 a_2724_1256# VPWR 0.20782f
C6945 _246_.B2 a_59796_29480# 0.00287f
C6946 a_18292_25156# a_18380_25112# 0.28563f
C6947 a_3172_31048# VPWR 0.20993f
C6948 a_50636_13703# a_50548_13800# 0.28563f
C6949 a_5052_18840# a_4940_18407# 0.02634f
C6950 a_64188_14136# a_64212_13800# 0.00172f
C6951 a_30028_20408# a_30476_20408# 0.0131f
C6952 a_32180_20452# a_31820_20408# 0.08717f
C6953 a_23084_30951# a_24196_31048# 0.00193f
C6954 a_37420_16839# a_37332_16936# 0.28563f
C6955 a_39268_18840# a_39648_19435# 0.00372f
C6956 a_18816_29931# uio_out[5] 0.0504f
C6957 a_31396_26724# a_31484_26680# 0.28563f
C6958 a_29020_1592# VPWR 0.29679f
C6959 a_49604_22020# VPWR 0.01537f
C6960 _478_.D a_53460_24776# 0.00356f
C6961 a_1380_1636# a_1468_1592# 0.28563f
C6962 a_4964_1636# a_5412_1636# 0.01328f
C6963 a_58140_12568# a_58028_12135# 0.02634f
C6964 _460_.Q a_35652_25156# 0.04816f
C6965 a_18740_23588# a_18716_23111# 0.00172f
C6966 a_14796_23544# a_14796_23111# 0.05841f
C6967 a_61836_25515# a_62796_25640# 0.00284f
C6968 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN 0.0053f
C6969 a_58388_12232# a_58476_10567# 0.00151f
C6970 a_2364_11000# a_2364_10567# 0.05841f
C6971 a_55812_11044# a_55452_11000# 0.08707f
C6972 VPWR uio_oe[0] 0.08962f
C6973 _371_.ZN _352_.A2 0.01394f
C6974 _350_.A1 _296_.ZN 0.5907f
C6975 a_16240_26795# a_16796_27209# 0.8399f
C6976 a_19860_26724# a_19948_26680# 0.28563f
C6977 _343_.A2 _340_.ZN 0.57168f
C6978 a_49896_18909# a_51308_18407# 0.00984f
C6979 _268_.A2 _274_.A2 0.48079f
C6980 a_45596_1159# a_46044_1159# 0.0131f
C6981 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_63852_23544# 0.01466f
C6982 _474_.Q a_47524_22021# 0.10776f
C6983 a_49492_18840# VPWR 0.36635f
C6984 a_63428_18884# a_63876_18884# 0.01328f
C6985 _395_.A3 _427_.B2 1.48483f
C6986 a_19948_20408# VPWR 0.31239f
C6987 _397_.A2 a_47700_28292# 0.00179f
C6988 a_60285_30600# ui_in[2] 0.03039f
C6989 a_54556_12568# VPWR 0.31389f
C6990 a_2724_15748# a_3172_15748# 0.01328f
C6991 _402_.A1 _399_.ZN 0.06572f
C6992 _355_.C a_24080_25227# 0.01209f
C6993 a_11324_2727# a_11460_1636# 0.00154f
C6994 a_13340_29383# a_13252_29480# 0.28563f
C6995 a_21540_28292# _455_.D 0.00124f
C6996 a_49764_15368# a_50212_15368# 0.01328f
C6997 _355_.C a_18760_29032# 0.00788f
C6998 _251_.A1 _272_.B1 0.91391f
C6999 _395_.A2 _384_.A3 0.18478f
C7000 _447_.Q _301_.Z 0.05018f
C7001 a_57132_18407# a_57492_18504# 0.08663f
C7002 a_2364_7431# a_2724_7528# 0.08717f
C7003 a_51644_15271# a_51556_15368# 0.28563f
C7004 a_1468_8999# a_1828_9096# 0.08717f
C7005 _252_.B a_60068_27912# 0.05918f
C7006 a_55028_10664# VPWR 0.20614f
C7007 a_3260_5863# a_3620_5960# 0.08717f
C7008 _294_.A2 a_40264_30320# 0.21963f
C7009 a_60212_25156# a_60524_25640# 0.00685f
C7010 a_4156_4295# a_4852_4392# 0.01227f
C7011 _250_.B _250_.A2 0.00443f
C7012 a_56036_23208# _427_.ZN 0.01116f
C7013 a_52988_15271# a_53660_15271# 0.00544f
C7014 a_3172_15368# VPWR 0.20993f
C7015 _437_.A1 _443_.D 1.04896f
C7016 a_20532_22020# a_20620_21976# 0.28563f
C7017 a_16588_21976# a_17036_21976# 0.01288f
C7018 a_31708_15271# VPWR 0.29679f
C7019 _355_.C a_26468_27912# 0.04118f
C7020 a_65756_2727# a_65668_2824# 0.28563f
C7021 a_38576_22504# _302_.Z 0.36671f
C7022 a_34732_16839# a_35180_16839# 0.01288f
C7023 a_49852_30951# a_49764_31048# 0.28563f
C7024 a_23980_23544# a_23892_22020# 0.00151f
C7025 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN 0.00984f
C7026 a_38676_16936# a_38564_15748# 0.02666f
C7027 a_64324_17316# VPWR 0.20554f
C7028 _452_.CLK a_42932_16936# 0.00139f
C7029 a_30948_23208# a_31036_21543# 0.00151f
C7030 _404_.A1 a_47600_27912# 0.01483f
C7031 _251_.A1 a_60212_25156# 0.28547f
C7032 a_30388_23588# a_30836_23588# 0.01328f
C7033 a_1468_7431# VPWR 0.29679f
C7034 a_25124_1256# VPWR 0.20348f
C7035 a_3260_4295# VPWR 0.30487f
C7036 a_24080_25227# a_24636_25641# 0.8399f
C7037 a_46628_1256# a_47076_1256# 0.01328f
C7038 a_57580_17272# vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN 0.00262f
C7039 a_25660_2727# a_26108_2727# 0.0131f
C7040 a_61164_13703# a_61524_13800# 0.08707f
C7041 a_15580_29383# VPWR 0.32517f
C7042 a_47076_13800# a_47524_13800# 0.01328f
C7043 _437_.A1 a_38772_28292# 0.00717f
C7044 a_7180_30951# VPWR 0.31145f
C7045 _452_.CLK _303_.ZN 0.00229f
C7046 a_19164_23111# a_19188_22020# 0.0016f
C7047 a_47948_16839# a_48308_16936# 0.08707f
C7048 a_7068_1159# a_6980_1256# 0.28563f
C7049 a_22059_26399# a_22344_26399# 0.00277f
C7050 a_51444_10664# a_51420_9432# 0.0016f
C7051 a_42820_1636# VPWR 0.23424f
C7052 a_40468_16936# VPWR 0.20637f
C7053 a_55004_12568# a_55028_12232# 0.00172f
C7054 a_6756_29860# a_6844_29816# 0.28563f
C7055 a_2812_29816# a_3260_29816# 0.01288f
C7056 a_19724_25112# a_19612_24679# 0.02634f
C7057 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _268_.A1 0.02509f
C7058 a_32964_17316# a_33412_17316# 0.01328f
C7059 a_62620_15271# a_62756_14180# 0.00154f
C7060 _459_.CLK a_34084_28776# 0.0088f
C7061 _251_.A1 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN 0.02768f
C7062 a_5188_2824# VPWR 0.20815f
C7063 a_24452_1636# a_24316_1159# 0.00168f
C7064 a_48060_1592# a_48508_1592# 0.01288f
C7065 a_52004_1636# a_52092_1592# 0.28563f
C7066 _384_.A3 a_50196_22805# 0.0047f
C7067 a_62308_11044# a_62756_11044# 0.01328f
C7068 a_58028_17272# VPWR 0.35213f
C7069 _452_.CLK a_33164_20408# 0.01227f
C7070 a_32516_20072# a_32516_18884# 0.05841f
C7071 a_26152_26841# VPWR 0.00224f
C7072 _337_.ZN a_29348_25940# 0.00718f
C7073 a_4156_23111# a_4940_23111# 0.00443f
C7074 _242_.Z a_58052_26724# 0.04119f
C7075 a_39256_18559# VPWR 0.00204f
C7076 a_51756_18407# a_52116_18504# 0.08717f
C7077 _373_.A2 a_26970_29480# 0.011f
C7078 a_53460_18504# a_53548_16839# 0.00151f
C7079 _395_.A1 clk 0.12402f
C7080 a_41700_2824# a_41564_1592# 0.00154f
C7081 a_45508_2824# a_45508_1636# 0.05841f
C7082 a_51220_18504# VPWR 0.20595f
C7083 a_15244_25112# VPWR 0.29679f
C7084 a_30924_20408# VPWR 0.31594f
C7085 a_19948_27815# a_20308_27912# 0.08663f
C7086 _475_.Q _473_.Q 0.97272f
C7087 a_4852_27912# a_5300_27912# 0.01328f
C7088 a_24652_30951# VPWR 0.31184f
C7089 a_31484_26680# VPWR 0.3205f
C7090 _435_.A3 _304_.A1 0.00305f
C7091 a_1468_12135# VPWR 0.29679f
C7092 a_34160_20523# _319_.A2 0.04554f
C7093 a_26468_2824# a_26916_2824# 0.01328f
C7094 a_39548_15704# a_39684_15368# 0.00168f
C7095 _450_.D a_42896_18504# 0.25728f
C7096 a_17932_27815# uio_out[7] 0.00512f
C7097 a_19076_21640# a_18964_20452# 0.02666f
C7098 _397_.A2 a_48708_29816# 0.00584f
C7099 a_3620_15748# VPWR 0.22347f
C7100 a_50660_15368# VPWR 0.2267f
C7101 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN a_63068_19975# 0.00154f
C7102 a_23892_22020# a_23532_21976# 0.08707f
C7103 a_54108_15271# VPWR 0.32871f
C7104 a_47524_14180# a_47972_14180# 0.01328f
C7105 a_35292_17272# a_35204_15748# 0.00151f
C7106 _452_.CLK a_36100_17316# 0.002f
C7107 a_35628_16839# VPWR 0.31389f
C7108 a_47524_1256# VPWR 0.20348f
C7109 _404_.A1 _424_.A2 0.00743f
C7110 a_24652_30951# a_24564_31048# 0.28563f
C7111 a_61948_14136# a_61860_12612# 0.00151f
C7112 _358_.A2 a_31732_25156# 0.00474f
C7113 _251_.A1 VPWR 4.37176f
C7114 a_25792_30301# VPWR 0.19143f
C7115 _424_.A1 a_53796_20452# 0.00597f
C7116 a_33860_17316# VPWR 0.20799f
C7117 _371_.A1 a_33476_27912# 0.00505f
C7118 a_48956_1592# VPWR 0.30013f
C7119 a_17844_23208# a_17844_22020# 0.05841f
C7120 a_18044_1159# a_18404_1256# 0.08717f
C7121 a_48060_12135# a_48420_12232# 0.08717f
C7122 _424_.B1 _411_.A2 0.04447f
C7123 a_62060_12135# a_62508_12135# 0.01288f
C7124 a_31820_23544# a_31932_23111# 0.02634f
C7125 a_11100_1592# a_11548_1592# 0.01288f
C7126 a_15044_1636# a_15132_1592# 0.28563f
C7127 a_11236_29480# a_11684_29480# 0.01328f
C7128 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I a_64884_26724# 0.03821f
C7129 a_10116_29860# a_9756_29816# 0.08707f
C7130 _350_.A2 _369_.ZN 0.06507f
C7131 a_48420_31048# a_48868_31048# 0.01328f
C7132 a_55812_15368# a_55812_14180# 0.05841f
C7133 _390_.ZN _267_.ZN 0.00317f
C7134 a_59844_11044# a_59820_10567# 0.00172f
C7135 a_27588_2824# VPWR 0.2304f
C7136 _438_.A2 _434_.ZN 0.00372f
C7137 a_55900_11000# a_56012_10567# 0.02634f
C7138 vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I 0.00176f
C7139 _251_.A1 a_59332_29816# 0.01325f
C7140 _324_.C a_43232_29480# 0.00126f
C7141 _459_.CLK a_19500_27815# 0.00525f
C7142 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN a_57604_14180# 0.0404f
C7143 a_16140_24679# a_16052_24776# 0.28563f
C7144 _350_.A1 a_29232_29931# 0.05806f
C7145 a_3260_23111# a_3172_23208# 0.28563f
C7146 a_24540_24679# a_24988_24679# 0.01288f
C7147 a_54692_15748# a_54780_15704# 0.28563f
C7148 a_32604_19975# a_33052_19975# 0.0131f
C7149 a_4068_7528# a_4852_7528# 0.00276f
C7150 a_3172_9096# a_3620_9096# 0.01328f
C7151 a_48420_14180# VPWR 0.20952f
C7152 a_33948_18407# a_34732_18407# 0.00443f
C7153 a_3260_18407# a_3620_18504# 0.08717f
C7154 a_64772_4392# a_65220_4392# 0.01328f
C7155 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN 0.623f
C7156 a_33376_23659# a_33764_24073# 0.00393f
C7157 a_55700_25156# vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN 0.00236f
C7158 a_12356_29480# VPWR 0.22423f
C7159 a_62956_12135# VPWR 0.31547f
C7160 _386_.ZN _411_.A2 0.00348f
C7161 a_37084_15704# a_37532_15704# 0.01288f
C7162 a_49316_31048# VPWR 0.20832f
C7163 _340_.ZN a_24952_29032# 0.01768f
C7164 _290_.ZN a_34708_29860# 0.0029f
C7165 _358_.A3 a_35652_26344# 0.02091f
C7166 a_48284_15704# a_48284_15271# 0.05841f
C7167 a_52228_15748# a_52092_15271# 0.00168f
C7168 a_25436_24679# VPWR 0.299f
C7169 a_65668_4392# VPWR 0.21209f
C7170 a_5300_7528# VPWR 0.21406f
C7171 _437_.A1 a_39796_27912# 0.12547f
C7172 a_37980_15704# VPWR 0.3582f
C7173 a_30795_29977# uo_out[6] 0.01182f
C7174 a_53100_18407# a_53548_18407# 0.0131f
C7175 _409_.ZN a_49740_29383# 0.00275f
C7176 a_30388_22020# a_30836_22020# 0.01328f
C7177 a_38506_26724# VPWR 0.01466f
C7178 a_67684_15368# a_67684_14180# 0.05841f
C7179 a_53996_18407# VPWR 0.3305f
C7180 _384_.A3 _427_.A2 0.50108f
C7181 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN a_55140_28292# 0.01924f
C7182 _384_.A3 a_51196_21543# 0.00175f
C7183 _455_.Q a_25300_26344# 0.00127f
C7184 a_5052_1592# a_5188_1256# 0.00168f
C7185 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN VPWR 0.79218f
C7186 a_1380_12612# a_1828_12612# 0.01328f
C7187 a_34084_28776# uo_out[7] 0.08134f
C7188 a_48060_2727# a_48508_2727# 0.0131f
C7189 _388_.B _393_.A1 0.12388f
C7190 a_48956_18407# a_49092_17316# 0.00154f
C7191 _325_.A2 _325_.ZN 0.93177f
C7192 _290_.ZN a_35204_31048# 0.01535f
C7193 a_50884_17316# a_50860_16839# 0.00172f
C7194 _231_.ZN vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN 0.11579f
C7195 a_46940_17272# a_47052_16839# 0.02634f
C7196 a_45708_17272# VPWR 0.31817f
C7197 a_24900_23208# a_24788_22020# 0.02666f
C7198 a_29468_1159# a_29380_1256# 0.28563f
C7199 a_59372_12135# a_59284_12232# 0.28563f
C7200 a_62620_1592# VPWR 0.3289f
C7201 _424_.B1 _399_.ZN 1.42143f
C7202 a_18404_1636# a_18044_1592# 0.08707f
C7203 _474_.CLK a_53012_18504# 0.00546f
C7204 a_47860_23208# VPWR 0.14301f
C7205 a_18716_21543# VPWR 0.32683f
C7206 a_16612_29860# a_17060_29860# 0.01328f
C7207 _397_.A1 clk 0.00278f
C7208 a_44340_26183# a_44688_26399# 0.00277f
C7209 _474_.Q a_48956_18407# 0.00393f
C7210 _237_.A1 a_59572_29076# 0.00418f
C7211 a_44812_17272# a_45260_17272# 0.01255f
C7212 a_49764_2824# VPWR 0.21599f
C7213 a_66788_11044# a_66764_10567# 0.00172f
C7214 a_49292_10567# a_49740_10567# 0.01288f
C7215 a_61724_1592# a_62172_1592# 0.01288f
C7216 _402_.ZN _473_.Q 0.0038f
C7217 _324_.C a_46156_25112# 0.0181f
C7218 a_1828_23208# a_2276_23208# 0.01328f
C7219 _248_.B1 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN 0.05831f
C7220 a_23196_23111# a_23556_23208# 0.08707f
C7221 a_55452_21543# VPWR 0.30531f
C7222 _404_.A1 a_46804_28292# 0.00106f
C7223 _362_.B a_33188_25940# 0.00103f
C7224 _397_.A2 _402_.A1 0.29081f
C7225 a_60401_30300# _255_.I 0.18586f
C7226 a_49180_9432# VPWR 0.32016f
C7227 a_55452_14136# VPWR 0.31389f
C7228 a_17484_21543# a_17932_21543# 0.0131f
C7229 _325_.A1 a_41440_23208# 0.01251f
C7230 a_26468_31048# VPWR 0.20586f
C7231 a_29716_31048# a_29856_29123# 0.00145f
C7232 _452_.CLK a_34396_24679# 0.01103f
C7233 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I a_57604_14180# 0.00109f
C7234 a_55956_25940# a_56516_26344# 0.3026f
C7235 a_57044_12232# VPWR 0.23066f
C7236 a_44388_15748# a_44028_15704# 0.08707f
C7237 a_3260_29816# a_3260_29383# 0.05841f
C7238 a_7204_29860# a_7068_29383# 0.00168f
C7239 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I a_64748_23544# 0.0016f
C7240 a_48868_2824# a_49316_2824# 0.01328f
C7241 a_23196_29816# a_23084_29383# 0.02634f
C7242 _384_.ZN _412_.A1 0.0209f
C7243 _303_.ZN a_43668_19668# 0.01165f
C7244 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.01028f
C7245 a_35723_20569# a_36008_20569# 0.00277f
C7246 a_39684_20452# a_39772_20408# 0.28563f
C7247 a_49600_30180# _409_.ZN 0.22193f
C7248 a_30796_24463# VPWR 0.39641f
C7249 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN 0.00147f
C7250 a_62532_20072# VPWR 0.20348f
C7251 _448_.Q _323_.A3 0.80014f
C7252 a_9532_2727# a_9444_2824# 0.28563f
C7253 a_51780_15748# VPWR 0.20622f
C7254 a_54556_21543# a_55004_21543# 0.01255f
C7255 _362_.ZN VPWR 0.33617f
C7256 hold2.Z a_42796_23981# 0.27406f
C7257 a_50436_9476# a_50076_9432# 0.08717f
C7258 a_51780_9476# a_52228_9476# 0.01328f
C7259 a_24196_31048# uio_out[2] 0.00329f
C7260 a_36288_31048# _462_.D 0.02546f
C7261 a_54556_14136# a_55004_14136# 0.0131f
C7262 _379_.Z a_17472_28363# 0.00665f
C7263 a_58836_14180# a_58924_14136# 0.28563f
C7264 a_61188_15368# a_61164_13703# 0.00131f
C7265 _412_.ZN a_51332_24372# 0.44033f
C7266 a_20672_30301# a_22100_29480# 0.00172f
C7267 _237_.A1 _257_.B 0.00437f
C7268 a_59732_13800# a_59844_12612# 0.02666f
C7269 a_55924_13800# a_55900_12568# 0.0016f
C7270 _325_.B a_43892_20072# 0.01325f
C7271 _287_.A2 a_31396_26724# 0.0016f
C7272 _252_.ZN a_60492_28248# 0.04943f
C7273 a_37444_26344# VPWR 0.20348f
C7274 a_31844_23208# a_31732_22020# 0.02666f
C7275 a_18716_24679# a_18740_23588# 0.0016f
C7276 _345_.A2 _454_.D 0.12082f
C7277 a_3172_24776# a_3172_23588# 0.05841f
C7278 _460_.D a_32592_25227# 0.2885f
C7279 a_12892_1159# VPWR 0.29679f
C7280 a_55924_12232# a_56372_12232# 0.01328f
C7281 a_932_7908# a_1380_7908# 0.01328f
C7282 a_40444_1159# a_40804_1256# 0.08717f
C7283 a_24900_1636# a_25348_1636# 0.01328f
C7284 a_15604_21640# VPWR 0.20348f
C7285 hold2.Z a_42784_25640# 0.00225f
C7286 a_52228_17316# a_51868_17272# 0.08707f
C7287 a_58020_27508# VPWR 0.88418f
C7288 _427_.B1 _427_.B2 0.35812f
C7289 a_46268_10567# a_46180_10664# 0.28563f
C7290 _327_.A2 a_45260_17272# 0.00176f
C7291 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _474_.CLK 0.02002f
C7292 a_54244_18884# a_54332_18840# 0.28563f
C7293 _459_.CLK _336_.A1 0.15425f
C7294 a_65756_23111# VPWR 0.34587f
C7295 _452_.CLK a_36188_25112# 0.00442f
C7296 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN 0.0139f
C7297 a_30240_24776# a_31168_24419# 1.16391f
C7298 a_4156_23544# VPWR 0.30552f
C7299 _474_.CLK a_52852_24372# 0.00205f
C7300 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN _427_.ZN 0.01628f
C7301 a_63652_9476# VPWR 0.21214f
C7302 a_64772_3204# VPWR 0.20727f
C7303 a_16140_21543# a_16500_21640# 0.08717f
C7304 a_61636_20072# a_62084_20072# 0.01328f
C7305 a_62196_23588# clk 0.00646f
C7306 a_4156_6296# VPWR 0.30552f
C7307 a_3260_13703# VPWR 0.30487f
C7308 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_54892_26680# 0.00426f
C7309 _416_.A1 _436_.B 0.02526f
C7310 _452_.CLK a_35504_18955# 0.11297f
C7311 _427_.ZN a_53108_21640# 0.01608f
C7312 a_50884_15748# a_51332_15748# 0.01328f
C7313 a_47300_15748# a_47388_15704# 0.28563f
C7314 a_46180_11044# VPWR 0.20348f
C7315 a_66988_19975# a_67348_20072# 0.0869f
C7316 _231_.ZN vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN 0.09978f
C7317 _350_.A1 a_30596_28292# 0.00798f
C7318 a_33052_18840# VPWR 0.29736f
C7319 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I VPWR 0.79508f
C7320 a_16140_26247# VPWR 0.31993f
C7321 a_20508_2727# a_20868_2824# 0.08717f
C7322 _275_.A2 _267_.ZN 0.04102f
C7323 _399_.ZN _218_.ZN 0.00594f
C7324 _304_.B _421_.A1 0.03808f
C7325 _330_.A2 a_39324_17272# 0.01121f
C7326 a_2364_9432# a_2364_8999# 0.05841f
C7327 _359_.B _455_.Q 0.00683f
C7328 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN clk 0.08707f
C7329 a_28460_21976# a_28372_20452# 0.00151f
C7330 a_15156_20452# a_15604_20452# 0.01328f
C7331 a_52092_14136# a_51980_13703# 0.02634f
C7332 _474_.Q a_49856_20936# 0.00269f
C7333 a_62756_14180# a_62844_14136# 0.28563f
C7334 _417_.Z _474_.D 0.0066f
C7335 a_50300_12568# a_50748_12568# 0.01288f
C7336 a_66676_13800# a_66788_12612# 0.02666f
C7337 _313_.ZN a_36288_23208# 0.00988f
C7338 _424_.A1 a_51877_21236# 0.00101f
C7339 _335_.ZN a_37324_28776# 0.00371f
C7340 vgaringosc.workerclkbuff_notouch_.I uio_in[1] 0.03938f
C7341 a_20868_24776# a_20980_23588# 0.02666f
C7342 a_35292_1159# VPWR 0.34116f
C7343 a_51868_1159# a_51780_1256# 0.28563f
C7344 a_56572_23111# vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.00111f
C7345 _451_.Q _301_.Z 0.10529f
C7346 a_58388_20452# vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN 0.00602f
C7347 a_31620_1636# a_32292_1636# 0.00347f
C7348 a_45508_31048# a_45416_29885# 0.00998f
C7349 _319_.A3 VPWR 1.66847f
C7350 a_36548_26344# a_36996_26344# 0.01328f
C7351 a_64748_23544# VPWR 0.30098f
C7352 _424_.A2 a_47259_20127# 0.00145f
C7353 a_34448_25597# a_34396_24679# 0.00818f
C7354 a_3172_10664# a_3620_10664# 0.01328f
C7355 a_57132_10567# a_57492_10664# 0.08707f
C7356 a_11772_1159# a_12444_1159# 0.00544f
C7357 _324_.C vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.06002f
C7358 _455_.D a_20956_24679# 0.00173f
C7359 _355_.C _457_.D 1.08963f
C7360 a_32740_23208# a_33188_23208# 0.01328f
C7361 a_5052_21976# VPWR 0.33516f
C7362 a_64996_31048# vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.00439f
C7363 _256_.A2 a_60793_29860# 0.00106f
C7364 _402_.A1 _330_.A1 0.5006f
C7365 a_36172_24463# a_36516_24831# 0.00275f
C7366 a_27028_23588# VPWR 0.23512f
C7367 a_16612_29480# a_16588_28248# 0.0016f
C7368 a_27452_21543# a_27364_21640# 0.28563f
C7369 a_14708_21640# a_15156_21640# 0.01328f
C7370 _467_.D a_15692_28248# 0.0048f
C7371 a_64972_13703# VPWR 0.3241f
C7372 a_2724_18884# a_2812_18840# 0.28563f
C7373 a_15132_2727# VPWR 0.31143f
C7374 a_41700_2824# a_41788_1159# 0.0027f
C7375 _246_.B2 a_60276_29032# 0.05637f
C7376 _399_.A1 a_48321_23208# 0.03435f
C7377 a_50420_23233# VPWR 0.03902f
C7378 _355_.C _454_.Q 0.14661f
C7379 _459_.CLK a_33776_29123# 0.03161f
C7380 _284_.B _441_.A2 0.00118f
C7381 _448_.Q a_37964_18191# 0.00132f
C7382 _287_.A2 VPWR 1.0991f
C7383 a_50436_30689# _409_.ZN 0.00216f
C7384 _274_.ZN a_51457_29861# 0.07271f
C7385 a_59844_11044# VPWR 0.20622f
C7386 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN a_56720_26344# 0.00192f
C7387 a_16796_27209# VPWR 0.3968f
C7388 a_17820_30951# a_17956_29860# 0.00154f
C7389 _371_.A3 _336_.A1 0.05376f
C7390 _260_.ZN a_44290_21236# 0.00132f
C7391 _462_.D a_36160_29535# 0.00242f
C7392 a_62172_15704# a_62620_15704# 0.0131f
C7393 a_65668_15748# a_65308_15704# 0.0869f
C7394 a_4940_27815# VPWR 0.31954f
C7395 _407_.A1 _411_.A2 0.02645f
C7396 a_64300_23111# a_64748_23111# 0.012f
C7397 a_31932_2727# a_31844_2824# 0.28563f
C7398 _282_.ZN _279_.Z 0.0197f
C7399 _457_.D a_24636_25641# 0.2313f
C7400 a_26020_31048# uio_out[2] 0.01582f
C7401 _421_.A1 VPWR 1.17941f
C7402 a_61412_9476# a_61052_9432# 0.08717f
C7403 a_62756_9476# a_63204_9476# 0.01328f
C7404 a_2364_7864# a_2812_7864# 0.0131f
C7405 a_4964_7908# a_4604_7864# 0.08674f
C7406 _437_.A1 a_39536_23588# 0.01692f
C7407 a_3260_6296# a_3708_6296# 0.0131f
C7408 a_3260_23544# a_3708_23544# 0.0131f
C7409 a_12804_1256# a_13252_1256# 0.01328f
C7410 a_18628_31048# a_19076_31048# 0.01328f
C7411 a_27228_26680# a_27676_26680# 0.01222f
C7412 a_4156_4728# a_4604_4728# 0.01222f
C7413 a_49652_29480# _395_.A1 0.00273f
C7414 a_59820_14136# a_59820_13703# 0.05841f
C7415 a_2364_13703# a_2812_13703# 0.0131f
C7416 a_20756_20452# a_20844_20408# 0.28563f
C7417 _441_.A2 a_43245_24373# 0.0016f
C7418 a_4156_30951# a_4068_31048# 0.28563f
C7419 a_3260_29383# a_3708_29383# 0.0131f
C7420 a_51791_30644# _268_.A2 0.00149f
C7421 _397_.A2 _424_.B1 0.02546f
C7422 a_57604_12612# a_57244_12568# 0.08707f
C7423 a_4156_12568# a_4156_12135# 0.05841f
C7424 a_8772_1636# VPWR 0.22925f
C7425 a_60180_13800# a_60268_12135# 0.00151f
C7426 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN VPWR 0.7334f
C7427 _412_.B2 a_50084_24328# 0.00116f
C7428 _474_.CLK a_56036_23208# 0.04935f
C7429 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN a_62420_22020# 0.00722f
C7430 a_66228_20452# VPWR 0.21556f
C7431 a_57468_1159# VPWR 0.36405f
C7432 _304_.B a_55676_28248# 0.00464f
C7433 a_62844_1159# a_63204_1256# 0.08717f
C7434 _350_.A1 _223_.I 0.08343f
C7435 a_34980_1636# a_35068_1592# 0.28563f
C7436 a_38564_1636# a_39012_1636# 0.01328f
C7437 _431_.A3 _452_.Q 0.00386f
C7438 a_3172_16936# a_3620_16936# 0.01328f
C7439 a_67660_12135# a_67684_11044# 0.0016f
C7440 a_66204_18840# VPWR 0.33522f
C7441 a_45284_11044# a_45732_11044# 0.01328f
C7442 _268_.A1 _416_.A1 0.08786f
C7443 a_68108_10567# a_68020_10664# 0.28563f
C7444 _304_.B _409_.ZN 0.02139f
C7445 a_59484_1592# a_59484_1159# 0.05841f
C7446 a_33412_18504# a_33412_17316# 0.05841f
C7447 _437_.A1 a_35616_24776# 0.00233f
C7448 _424_.A2 _419_.Z 1.22711f
C7449 a_20420_2824# a_20284_1592# 0.00154f
C7450 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_55700_25156# 0.00136f
C7451 _358_.A3 a_32380_26247# 0.01752f
C7452 a_27924_22020# VPWR 0.20622f
C7453 _397_.A2 _386_.ZN 0.7362f
C7454 _398_.C a_52852_24372# 0.29825f
C7455 a_34308_18884# a_34396_18840# 0.28563f
C7456 _419_.A4 _417_.A2 0.41746f
C7457 _465_.D a_18816_29931# 0.28627f
C7458 _359_.B a_42908_30951# 0.00129f
C7459 a_32156_18840# a_32604_18840# 0.0131f
C7460 a_37532_2727# VPWR 0.31143f
C7461 a_59260_23111# a_59708_23111# 0.01222f
C7462 a_58836_13800# VPWR 0.20657f
C7463 a_1020_26247# a_1380_26344# 0.08717f
C7464 a_15244_26247# a_15692_26247# 0.0131f
C7465 _352_.A2 _336_.A2 2.31621f
C7466 a_14148_29860# VPWR 0.20845f
C7467 a_58364_25112# vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN 0.00114f
C7468 a_66428_11000# VPWR 0.32178f
C7469 a_63988_16936# a_63876_15748# 0.02666f
C7470 _290_.ZN _335_.ZN 0.07308f
C7471 a_3708_15271# a_4068_15368# 0.08717f
C7472 a_24988_23111# VPWR 0.31547f
C7473 a_64300_23544# a_64300_23111# 0.05841f
C7474 a_33708_22505# a_34052_22137# 0.00275f
C7475 a_43400_18909# a_44752_18147# 0.00388f
C7476 _325_.ZN a_43824_18147# 0.03995f
C7477 a_42908_2727# a_43268_2824# 0.08717f
C7478 _452_.CLK a_33932_24073# 0.02788f
C7479 a_64972_16839# a_64884_16936# 0.28563f
C7480 a_63068_18407# a_63516_18407# 0.0131f
C7481 _437_.A1 a_38584_28292# 0.40753f
C7482 a_19636_23588# a_19276_23544# 0.08707f
C7483 _274_.A2 a_56572_29383# 0.00184f
C7484 a_4516_25156# a_4156_25112# 0.08674f
C7485 _267_.A2 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I 0.05248f
C7486 a_1916_25112# a_2364_25112# 0.0131f
C7487 a_62060_20408# a_62084_20072# 0.00172f
C7488 _474_.Q _417_.Z 0.44535f
C7489 a_67796_20072# a_67908_18884# 0.02666f
C7490 a_56348_14136# a_56372_13800# 0.00172f
C7491 a_49316_31048# a_49112_29885# 0.00809f
C7492 _459_.Q a_34084_28776# 1.27795f
C7493 a_26132_20452# a_26580_20452# 0.01328f
C7494 _359_.B a_39748_29480# 0.00182f
C7495 a_18716_30951# a_19076_31048# 0.08663f
C7496 _250_.A2 a_62644_26724# 0.00108f
C7497 a_1020_16839# a_932_16936# 0.28563f
C7498 _452_.CLK a_37408_18504# 0.06278f
C7499 a_59036_11000# a_58948_9476# 0.00151f
C7500 a_64100_12612# a_64548_12612# 0.01328f
C7501 a_22436_1636# VPWR 0.2085f
C7502 a_60380_12568# a_61052_12568# 0.00544f
C7503 a_19744_30301# a_19372_30345# 0.10745f
C7504 a_18816_29931# a_19204_30345# 0.00393f
C7505 _474_.CLK a_54444_19975# 0.02892f
C7506 _251_.A1 a_57156_27912# 0.04429f
C7507 _284_.ZN _284_.B 0.56346f
C7508 a_25124_28776# a_27460_28776# 0.00589f
C7509 a_54780_15704# a_55228_15704# 0.012f
C7510 _459_.CLK a_16612_29480# 0.00745f
C7511 a_55676_28248# VPWR 0.29679f
C7512 a_63516_15271# a_63876_15368# 0.08717f
C7513 a_10116_1636# a_9980_1159# 0.00168f
C7514 _424_.B1 a_48308_23588# 0.00391f
C7515 a_52452_11044# a_52092_11000# 0.08663f
C7516 a_61076_12232# a_61052_11000# 0.0016f
C7517 a_34644_18504# VPWR 0.24097f
C7518 a_58028_20408# vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.00224f
C7519 a_1828_26724# a_1916_26680# 0.28563f
C7520 a_42908_30951# _495_.I 0.00239f
C7521 a_64884_10664# a_65332_10664# 0.01328f
C7522 _409_.ZN VPWR 0.76155f
C7523 a_33776_29123# uo_out[7] 0.01101f
C7524 a_34172_1159# a_34620_1159# 0.0131f
C7525 _384_.ZN _473_.Q 0.10795f
C7526 a_18096_27165# a_17932_26247# 0.00119f
C7527 a_67684_21640# VPWR 0.20429f
C7528 _451_.Q _436_.ZN 0.02037f
C7529 a_37084_21543# a_37532_21543# 0.012f
C7530 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_63852_23111# 0.00424f
C7531 a_47972_12612# VPWR 0.20348f
C7532 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I a_63316_20452# 0.0015f
C7533 a_59932_2727# VPWR 0.31143f
C7534 a_66092_18407# a_66452_18504# 0.0869f
C7535 _412_.A1 a_51576_25896# 0.05401f
C7536 a_1916_29383# a_1828_29480# 0.28563f
C7537 a_38340_15368# a_38788_15368# 0.01328f
C7538 a_3620_20072# VPWR 0.22347f
C7539 _355_.C a_18816_29931# 0.06124f
C7540 a_63852_23544# a_64300_23544# 0.01255f
C7541 a_1916_15704# a_1916_15271# 0.05841f
C7542 a_60716_10567# VPWR 0.33016f
C7543 a_40220_15271# a_40132_15368# 0.28563f
C7544 _274_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN 0.06982f
C7545 a_58388_18884# VPWR 0.23728f
C7546 a_22660_23208# VPWR 0.20622f
C7547 a_62620_17272# a_62644_16936# 0.00172f
C7548 _252_.ZN a_60276_26724# 0.00441f
C7549 a_41564_15271# a_42236_15271# 0.00544f
C7550 _447_.Q _303_.ZN 0.47942f
C7551 _452_.CLK a_33708_22505# 0.00806f
C7552 a_4156_21976# a_4604_21976# 0.01222f
C7553 _424_.A2 _424_.A1 0.74625f
C7554 a_54332_2727# a_54244_2824# 0.28563f
C7555 a_65756_17272# a_66204_17272# 0.01255f
C7556 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN a_58500_21640# 0.0063f
C7557 _260_.A2 a_39781_24372# 0.00499f
C7558 a_19972_23208# a_20060_21543# 0.00151f
C7559 a_35204_1256# a_35652_1256# 0.01328f
C7560 a_18292_25156# a_17932_25112# 0.08707f
C7561 a_23444_23588# a_23084_23544# 0.08717f
C7562 a_26132_23588# a_26580_23588# 0.01328f
C7563 a_2724_31048# VPWR 0.20782f
C7564 a_2276_1256# VPWR 0.20634f
C7565 a_14236_2727# a_14684_2727# 0.0131f
C7566 a_63852_13703# a_64300_13703# 0.012f
C7567 a_50188_13703# a_50548_13800# 0.08707f
C7568 a_31732_20452# a_31820_20408# 0.28563f
C7569 _330_.A1 _424_.B1 0.04182f
C7570 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN 0.02297f
C7571 a_37067_19001# a_37352_19001# 0.00277f
C7572 _336_.Z _358_.A3 0.01633f
C7573 a_36972_16839# a_37332_16936# 0.08707f
C7574 _317_.A2 a_38228_20452# 0.00123f
C7575 a_48921_22020# VPWR 0.00558f
C7576 a_54220_10567# a_54244_9476# 0.0016f
C7577 a_40220_1592# a_40356_1256# 0.00168f
C7578 _478_.D a_53076_24776# 0.01415f
C7579 a_28572_1592# VPWR 0.29679f
C7580 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I 0.02461f
C7581 a_18716_30951# a_19164_30951# 0.012f
C7582 _460_.Q a_34155_25273# 0.00503f
C7583 a_1380_1636# a_1020_1592# 0.08707f
C7584 a_3260_25112# a_3260_24679# 0.05841f
C7585 _473_.Q a_49068_20408# 0.29514f
C7586 a_61836_25515# a_62404_25640# 0.00685f
C7587 a_1380_17316# a_1828_17316# 0.01328f
C7588 a_55364_11044# a_55452_11000# 0.28563f
C7589 a_58948_11044# a_59396_11044# 0.01328f
C7590 a_50324_16936# a_50772_16936# 0.01328f
C7591 a_44700_1592# a_45148_1592# 0.01288f
C7592 _474_.CLK _392_.A2 0.03214f
C7593 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN a_62084_18504# 0.0012f
C7594 _371_.ZN a_28364_28776# 0.00222f
C7595 _255_.I _238_.I 0.14707f
C7596 a_23084_29383# _340_.ZN 0.00299f
C7597 a_16240_26795# a_17168_27165# 1.16391f
C7598 a_18096_27165# a_19948_26680# 0.00553f
C7599 a_49896_18909# a_50860_18407# 0.00107f
C7600 _251_.A1 a_62796_25640# 0.00448f
C7601 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_63404_23544# 0.01876f
C7602 _402_.A1 a_43908_26841# 0.00101f
C7603 _324_.C _402_.ZN 0.75457f
C7604 a_48172_18840# VPWR 0.32769f
C7605 a_3708_27815# a_4156_27815# 0.0131f
C7606 a_19500_20408# VPWR 0.34288f
C7607 _370_.ZN _369_.ZN 0.26211f
C7608 _397_.A2 a_47476_28292# 0.02244f
C7609 a_54040_22366# a_54556_21543# 0.00664f
C7610 _281_.ZN a_50464_24908# 0.01099f
C7611 a_54108_12568# VPWR 0.31389f
C7612 a_15044_2824# a_15492_2824# 0.01328f
C7613 a_12892_29383# a_13252_29480# 0.08717f
C7614 a_56348_30951# _272_.B1 0.0057f
C7615 _409_.ZN a_50068_27508# 0.44477f
C7616 _419_.Z a_52136_20936# 0.00147f
C7617 a_1468_8999# a_1380_9096# 0.28563f
C7618 a_54580_10664# VPWR 0.20614f
C7619 a_33948_15704# a_33948_15271# 0.05841f
C7620 a_37892_15748# a_37756_15271# 0.00168f
C7621 a_57132_18407# a_57044_18504# 0.28563f
C7622 a_51196_15271# a_51556_15368# 0.08717f
C7623 a_53660_27815# a_53572_27912# 0.28563f
C7624 _424_.A2 _416_.A2 0.03096f
C7625 _324_.C vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.0319f
C7626 _252_.B a_59172_27912# 0.12604f
C7627 a_2364_7431# a_2276_7528# 0.28563f
C7628 a_3260_5863# a_3172_5960# 0.28563f
C7629 a_4156_4295# a_4068_4392# 0.28563f
C7630 a_2724_21640# a_2724_20452# 0.05841f
C7631 a_60212_25156# a_60084_25640# 0.00284f
C7632 _250_.B a_60940_28248# 0.00111f
C7633 a_45232_25987# a_45128_26031# 0.10745f
C7634 _362_.ZN _360_.ZN 0.00882f
C7635 hold2.I _305_.A2 0.00197f
C7636 _430_.ZN _304_.A1 0.41709f
C7637 a_2724_15368# VPWR 0.20782f
C7638 _437_.A1 a_36960_27912# 0.07002f
C7639 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN clk 0.12367f
C7640 a_65084_2727# a_65668_2824# 0.01675f
C7641 a_20532_22020# a_20172_21976# 0.08707f
C7642 a_38576_22504# a_39172_22504# 0.00736f
C7643 a_31260_15271# VPWR 0.29679f
C7644 a_55340_26680# VPWR 0.31744f
C7645 a_49404_30951# a_49764_31048# 0.08717f
C7646 a_1380_14180# a_1828_14180# 0.01328f
C7647 _473_.Q a_48776_20204# 0.05298f
C7648 a_63876_17316# VPWR 0.20348f
C7649 _404_.A1 a_47376_27912# 0.01896f
C7650 a_1020_7431# VPWR 0.30073f
C7651 a_24676_1256# VPWR 0.20348f
C7652 _397_.A2 _386_.A4 0.51669f
C7653 _287_.A2 _370_.B 0.02674f
C7654 a_24080_25227# a_25008_25597# 1.16391f
C7655 a_2812_4295# VPWR 0.30213f
C7656 a_15132_29383# VPWR 0.29679f
C7657 a_61164_13703# a_61076_13800# 0.28563f
C7658 a_56596_18504# vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I 0.00245f
C7659 a_6723_30644# VPWR 0.18305f
C7660 a_44276_17316# a_43664_17317# 0.09638f
C7661 a_47948_16839# a_47860_16936# 0.28563f
C7662 a_40020_16936# VPWR 0.20637f
C7663 a_42372_1636# VPWR 0.2184f
C7664 a_6620_1159# a_6980_1256# 0.08717f
C7665 a_65084_12568# a_64972_12135# 0.02634f
C7666 a_7740_1592# a_8188_1592# 0.012f
C7667 a_51084_12135# a_51532_12135# 0.01288f
C7668 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN _250_.A2 0.01897f
C7669 _452_.CLK _452_.D 0.11024f
C7670 a_6756_29860# a_6396_29816# 0.08707f
C7671 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN 0.02196f
C7672 a_35008_27533# VPWR 0.51906f
C7673 _251_.A1 a_62844_27815# 0.01396f
C7674 a_52004_1636# a_51644_1592# 0.08707f
C7675 a_4740_2824# VPWR 0.22891f
C7676 a_57580_17272# VPWR 0.3228f
C7677 _452_.CLK a_32716_20408# 0.00212f
C7678 a_49034_21640# VPWR 0.01498f
C7679 _475_.Q _281_.A1 1.21027f
C7680 a_38308_18559# VPWR 0.00246f
C7681 _337_.ZN a_29164_25940# 0.00775f
C7682 a_25204_26841# VPWR 0.00246f
C7683 _242_.Z a_56964_26724# 0.05375f
C7684 a_4156_24679# a_4940_24679# 0.00443f
C7685 _384_.ZN _381_.Z 0.03955f
C7686 _325_.B a_43380_16936# 0.00221f
C7687 a_51756_18407# a_51668_18504# 0.28563f
C7688 a_56572_1159# a_57020_1159# 0.0131f
C7689 a_65308_18840# a_65756_18840# 0.01255f
C7690 a_50772_18504# VPWR 0.21545f
C7691 a_14796_25112# VPWR 0.30073f
C7692 _474_.CLK _416_.A1 0.08308f
C7693 a_19948_27815# a_19860_27912# 0.28563f
C7694 _287_.A1 uo_out[2] 1.69228f
C7695 a_24196_31048# VPWR 0.36801f
C7696 a_30476_20408# VPWR 0.33105f
C7697 a_1020_12135# VPWR 0.30073f
C7698 a_33860_15748# a_34308_15748# 0.01328f
C7699 _451_.Q _439_.ZN 0.06039f
C7700 a_26468_27912# a_26916_27912# 0.01328f
C7701 _397_.A2 _407_.A1 0.48059f
C7702 a_17484_27815# uio_out[7] 0.00241f
C7703 _304_.B _305_.A2 1.82536f
C7704 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN a_57940_18884# 0.00102f
C7705 _346_.B uio_out[6] 0.09319f
C7706 _229_.I _267_.A2 0.00718f
C7707 a_27452_21543# a_27476_20452# 0.0016f
C7708 _452_.CLK a_37420_16839# 0.00239f
C7709 _251_.A1 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN 0.161f
C7710 a_3172_15748# VPWR 0.20993f
C7711 a_50212_15368# VPWR 0.2189f
C7712 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN a_62620_19975# 0.001f
C7713 a_23444_22020# a_23532_21976# 0.28563f
C7714 a_27028_22020# a_27476_22020# 0.01328f
C7715 _474_.CLK vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN 0.02092f
C7716 a_53660_15271# VPWR 0.30141f
C7717 a_45260_16839# a_45708_16839# 0.01288f
C7718 a_35180_16839# VPWR 0.32427f
C7719 a_57380_1256# a_58052_1256# 0.00347f
C7720 a_24196_31048# a_24564_31048# 0.02601f
C7721 a_47076_1256# VPWR 0.20348f
C7722 a_32476_29167# _223_.ZN 0.00205f
C7723 a_36636_2727# a_37084_2727# 0.0131f
C7724 a_57940_13800# a_58388_13800# 0.01328f
C7725 _358_.A2 a_30476_25112# 0.00501f
C7726 _362_.B a_35740_26247# 0.03367f
C7727 a_56348_30951# VPWR 0.32213f
C7728 a_33412_17316# VPWR 0.20644f
C7729 a_48508_1592# VPWR 0.29679f
C7730 vgaringosc.workerclkbuff_notouch_.I _275_.ZN 0.02495f
C7731 a_18044_1159# a_17956_1256# 0.28563f
C7732 a_61948_12568# a_61972_12232# 0.00172f
C7733 _395_.A3 a_52452_21236# 0.00133f
C7734 a_15044_1636# a_14684_1592# 0.08707f
C7735 a_48060_12135# a_47972_12232# 0.28563f
C7736 _474_.CLK a_49896_18909# 0.00401f
C7737 a_60964_27912# a_60828_26680# 0.00154f
C7738 a_67796_20072# a_67884_18407# 0.00151f
C7739 a_13252_29860# a_13700_29860# 0.01328f
C7740 a_9668_29860# a_9756_29816# 0.28563f
C7741 a_56404_27208# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.07819f
C7742 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_59260_23544# 0.00221f
C7743 a_35740_17272# a_36188_17272# 0.01288f
C7744 a_65532_11000# a_65980_11000# 0.01288f
C7745 a_49180_17272# a_49204_16936# 0.00172f
C7746 _294_.A2 _285_.Z 0.33328f
C7747 a_26916_2824# VPWR 0.23308f
C7748 _251_.A1 a_58116_30344# 0.02123f
C7749 a_58500_1636# a_58948_1636# 0.01328f
C7750 _438_.ZN _302_.Z 0.40946f
C7751 _293_.A2 uo_out[2] 0.02909f
C7752 a_2812_23111# a_3172_23208# 0.08717f
C7753 _459_.CLK a_17932_27815# 0.01166f
C7754 a_24092_23111# a_24540_23111# 0.01288f
C7755 a_15692_24679# a_16052_24776# 0.08717f
C7756 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN clk 0.08095f
C7757 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I 0.00209f
C7758 a_54692_15748# a_54332_15704# 0.08674f
C7759 a_47972_14180# VPWR 0.20952f
C7760 a_7876_2824# a_7964_1159# 0.0027f
C7761 a_3260_18407# a_3172_18504# 0.28563f
C7762 _287_.A2 _360_.ZN 0.00104f
C7763 _238_.ZN _247_.B 0.0013f
C7764 a_54892_18407# vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN 0.0195f
C7765 a_932_31048# a_932_29860# 0.05841f
C7766 a_11684_29480# VPWR 0.24433f
C7767 a_62508_12135# VPWR 0.31547f
C7768 a_25212_2727# a_25348_1636# 0.00154f
C7769 a_37444_2824# a_37892_2824# 0.01328f
C7770 _340_.ZN a_24304_29480# 0.0171f
C7771 a_54804_18504# vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN 0.04047f
C7772 a_48868_31048# VPWR 0.2062f
C7773 _358_.A3 a_35204_26344# 0.0128f
C7774 _290_.ZN a_34260_29860# 0.00342f
C7775 _330_.A1 a_39236_26344# 0.00184f
C7776 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN 0.09137f
C7777 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN 0.02571f
C7778 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN 0.00304f
C7779 a_24988_24679# VPWR 0.29679f
C7780 _305_.A2 VPWR 1.25377f
C7781 a_4852_7528# VPWR 0.22733f
C7782 a_65220_4392# VPWR 0.20921f
C7783 a_4604_3160# a_4740_2824# 0.00168f
C7784 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN VPWR 0.74741f
C7785 a_37532_15704# VPWR 0.3289f
C7786 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN 0.67418f
C7787 a_31088_30301# uo_out[6] 0.03415f
C7788 a_4604_9432# a_5052_9432# 0.01222f
C7789 _402_.A1 a_46580_23588# 0.00149f
C7790 a_63876_15368# a_63740_14136# 0.00154f
C7791 a_50300_14136# a_50748_14136# 0.01288f
C7792 _330_.A1 _330_.A2 0.25506f
C7793 _384_.A3 a_51332_24072# 0.10619f
C7794 _459_.CLK a_27676_26247# 0.01893f
C7795 a_53548_18407# VPWR 0.31547f
C7796 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN clk 0.02523f
C7797 _441_.A3 _304_.A1 0.03661f
C7798 a_33720_28776# uo_out[7] 0.00118f
C7799 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN VPWR 0.75126f
C7800 _388_.B a_47525_29480# 0.11737f
C7801 _325_.A2 a_43784_19369# 0.06886f
C7802 _334_.A1 _462_.D 0.00466f
C7803 _231_.ZN a_58364_25112# 0.0023f
C7804 a_45260_17272# VPWR 0.29679f
C7805 a_62172_1592# VPWR 0.3289f
C7806 a_29020_1159# a_29380_1256# 0.08717f
C7807 a_65780_10664# a_65756_9432# 0.0016f
C7808 a_67572_10664# a_67460_9476# 0.02666f
C7809 a_56348_12568# a_56260_11044# 0.00151f
C7810 a_58924_12135# a_59284_12232# 0.08707f
C7811 a_17956_1636# a_18044_1592# 0.28563f
C7812 a_21540_1636# a_21988_1636# 0.01328f
C7813 _279_.Z _324_.B 0.15654f
C7814 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN 0.79649f
C7815 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN a_56596_17316# 0.07124f
C7816 _383_.A2 _384_.ZN 0.60775f
C7817 a_30476_23544# a_30500_23208# 0.00172f
C7818 a_41440_23208# VPWR 0.01466f
C7819 _355_.ZN a_29163_24394# 0.00603f
C7820 _474_.CLK a_52564_18504# 0.00546f
C7821 _255_.I VPWR 0.99328f
C7822 a_17932_21543# VPWR 0.32173f
C7823 _395_.A1 a_49044_28292# 0.02001f
C7824 a_18716_26247# a_18740_25156# 0.0016f
C7825 _416_.A1 _261_.ZN 0.04785f
C7826 a_62844_11000# a_62956_10567# 0.02634f
C7827 _459_.Q a_33776_29123# 0.03353f
C7828 a_49316_2824# VPWR 0.20761f
C7829 _324_.C a_46068_25156# 0.0356f
C7830 _247_.ZN a_59260_26680# 0.00232f
C7831 a_23196_23111# a_23108_23208# 0.28563f
C7832 a_27172_24328# a_26548_24372# 0.00587f
C7833 a_28012_24679# a_27924_24776# 0.28563f
C7834 a_17844_24776# a_18628_24776# 0.00276f
C7835 _359_.B _393_.A1 0.00108f
C7836 _404_.A1 a_46580_28292# 0.00314f
C7837 a_55004_21543# VPWR 0.31233f
C7838 a_59332_29816# _255_.I 0.61549f
C7839 a_26020_31048# VPWR 0.20607f
C7840 a_52228_9476# VPWR 0.21296f
C7841 a_55004_14136# VPWR 0.31389f
C7842 a_59396_2824# a_59396_1636# 0.05841f
C7843 a_33412_18504# a_33860_18504# 0.01328f
C7844 _392_.A2 _393_.A3 0.04853f
C7845 _452_.CLK a_33612_24679# 0.00649f
C7846 a_56372_12232# VPWR 0.21291f
C7847 a_43940_15748# a_44028_15704# 0.28563f
C7848 a_39996_15704# a_40444_15704# 0.01288f
C7849 _407_.A1 _330_.A1 0.04736f
C7850 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN VPWR 0.74204f
C7851 a_52228_19368# a_52884_18884# 0.01565f
C7852 _419_.Z a_49988_21236# 0.00159f
C7853 a_49600_30180# a_49496_30345# 0.10745f
C7854 a_49112_29885# _409_.ZN 0.2489f
C7855 a_31168_24419# VPWR 0.18833f
C7856 a_62084_20072# VPWR 0.20348f
C7857 _416_.ZN a_46716_18407# 0.00627f
C7858 a_53548_16839# a_53572_15748# 0.0016f
C7859 a_9084_2727# a_9444_2824# 0.08717f
C7860 a_33188_21640# a_33164_20408# 0.0016f
C7861 a_61276_19975# a_61724_19975# 0.0131f
C7862 a_51332_15748# VPWR 0.20622f
C7863 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN a_59260_23544# 0.00153f
C7864 a_26712_29977# VPWR 0.00231f
C7865 a_46044_30951# a_45800_30345# 0.00105f
C7866 hold2.Z a_41488_24072# 0.00846f
C7867 _412_.A1 clkload0.Z 0.02319f
C7868 a_49988_9476# a_50076_9432# 0.28563f
C7869 a_20672_30301# a_21652_29480# 0.00172f
C7870 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN 0.00266f
C7871 a_59036_2727# a_59484_2727# 0.0131f
C7872 a_47076_12612# a_47524_12612# 0.01328f
C7873 _395_.A1 _284_.A2 0.03284f
C7874 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN VPWR 0.77878f
C7875 a_36996_26344# VPWR 0.20348f
C7876 a_30500_23208# a_30476_21976# 0.0016f
C7877 a_12444_1159# VPWR 0.30141f
C7878 a_40444_1159# a_40356_1256# 0.28563f
C7879 _345_.A2 a_22064_27912# 0.05215f
C7880 a_2724_20072# a_3172_20072# 0.01328f
C7881 a_2276_12232# a_2276_11044# 0.05841f
C7882 _424_.A2 _399_.ZN 0.03532f
C7883 a_64324_4392# a_64324_3204# 0.05841f
C7884 _324_.B _304_.ZN 0.62666f
C7885 a_59620_27208# _251_.ZN 0.00345f
C7886 a_15156_21640# VPWR 0.20348f
C7887 a_48384_26724# clkbuf_1_0__f_clk.I 0.00323f
C7888 a_20496_26344# a_21068_25112# 0.00105f
C7889 a_47836_17272# a_48284_17272# 0.01288f
C7890 a_51780_17316# a_51868_17272# 0.28563f
C7891 _340_.A2 a_25744_30345# 0.00121f
C7892 _451_.Q _303_.ZN 0.74233f
C7893 a_45820_10567# a_46180_10664# 0.08717f
C7894 a_59820_10567# a_60268_10567# 0.01288f
C7895 a_45148_1592# a_45148_1159# 0.05841f
C7896 a_22636_28248# a_22620_27599# 0.0019f
C7897 a_6084_2824# a_5948_1592# 0.00154f
C7898 a_35740_30951# _365_.ZN 0.07104f
C7899 a_64748_23111# VPWR 0.32068f
C7900 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I a_52639_30644# 0.00111f
C7901 a_57492_18884# a_57940_18884# 0.01328f
C7902 a_53436_18840# a_54332_18840# 0.00373f
C7903 a_33724_23111# _312_.ZN 0.00109f
C7904 _388_.B vgaringosc.workerclkbuff_notouch_.I 0.5005f
C7905 a_21764_23208# a_22212_23208# 0.01328f
C7906 _452_.CLK a_35740_25112# 0.01421f
C7907 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN a_63105_28293# 0.07802f
C7908 a_3708_6296# VPWR 0.33374f
C7909 a_3708_23544# VPWR 0.33374f
C7910 _324_.C _384_.ZN 0.05819f
C7911 a_63204_9476# VPWR 0.20595f
C7912 a_54420_21976# _427_.ZN 0.0147f
C7913 a_61748_23588# clk 0.00645f
C7914 a_2812_13703# VPWR 0.30213f
C7915 a_4068_29480# a_4068_28292# 0.05841f
C7916 a_59955_30600# a_60405_30644# 0.00184f
C7917 a_28348_21543# a_28796_21543# 0.01288f
C7918 a_16140_21543# a_16052_21640# 0.28563f
C7919 a_64324_3204# VPWR 0.22383f
C7920 a_55252_26724# a_55340_26680# 0.28563f
C7921 _325_.A1 _327_.A2 1.52508f
C7922 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_54444_26680# 0.00214f
C7923 _294_.A2 _371_.A1 0.2882f
C7924 _419_.A4 a_45920_20523# 0.00403f
C7925 a_45732_11044# VPWR 0.20348f
C7926 _274_.A1 a_53212_27815# 0.00156f
C7927 a_47300_15748# a_46940_15704# 0.08707f
C7928 a_59844_2824# a_60292_2824# 0.01328f
C7929 a_66988_19975# a_66900_20072# 0.28563f
C7930 a_10092_30951# a_10116_29860# 0.0016f
C7931 _416_.A1 _393_.A3 0.00316f
C7932 _397_.A4 _421_.B 0.0084f
C7933 _474_.CLK vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN 0.00297f
C7934 _350_.A1 a_29575_28293# 0.00161f
C7935 a_15692_26247# VPWR 0.32732f
C7936 a_32604_18840# VPWR 0.29679f
C7937 _438_.A2 a_39772_20408# 0.00506f
C7938 a_59708_23111# VPWR 0.34138f
C7939 a_20508_2727# a_20420_2824# 0.28563f
C7940 _448_.Q _437_.ZN 0.00517f
C7941 _304_.B a_45128_26031# 0.02099f
C7942 _330_.A2 a_40040_17675# 0.00123f
C7943 a_1380_1256# a_1828_1256# 0.01328f
C7944 a_55228_9432# a_55676_9432# 0.0131f
C7945 a_1828_31048# a_2276_31048# 0.01328f
C7946 _417_.Z a_50196_21640# 0.002f
C7947 a_62756_14180# a_62396_14136# 0.08707f
C7948 a_65892_14180# a_66340_14180# 0.01328f
C7949 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I 0.13053f
C7950 a_62868_13800# a_62844_12568# 0.0016f
C7951 a_49204_13800# a_49292_12135# 0.00151f
C7952 _313_.ZN a_36084_23208# 0.00292f
C7953 _379_.A2 a_22188_29383# 0.00297f
C7954 _335_.ZN a_36828_28776# 0.00371f
C7955 a_50548_12232# a_50660_11044# 0.02666f
C7956 a_51420_1159# a_51780_1256# 0.08717f
C7957 a_66676_12232# a_67124_12232# 0.01328f
C7958 _330_.A1 _304_.A1 0.69937f
C7959 a_34620_1159# VPWR 0.33964f
C7960 a_27676_1592# a_28124_1592# 0.01288f
C7961 a_31620_1636# a_31708_1592# 0.28563f
C7962 a_37532_21543# VPWR 0.32983f
C7963 _302_.Z a_43192_22504# 0.00259f
C7964 _267_.A1 a_56036_28292# 0.00449f
C7965 _424_.A2 a_46252_19759# 0.00219f
C7966 a_64300_23544# VPWR 0.29893f
C7967 a_57132_10567# a_57044_10664# 0.28563f
C7968 _231_.ZN clk 0.0416f
C7969 a_51620_19911# VPWR 0.36983f
C7970 uio_in[3] uio_in[2] 0.01021f
C7971 a_4604_21976# VPWR 0.33016f
C7972 a_57580_23544# vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN 0.00119f
C7973 _402_.A1 a_44388_27912# 0.00311f
C7974 a_37179_24831# a_37472_24419# 0.49319f
C7975 a_26580_23588# VPWR 0.21327f
C7976 a_27004_21543# a_27364_21640# 0.08707f
C7977 a_64300_13703# VPWR 0.34608f
C7978 a_2724_18884# a_2364_18840# 0.08717f
C7979 a_14684_2727# VPWR 0.31143f
C7980 _386_.ZN _393_.A1 0.33251f
C7981 _467_.D a_15244_28248# 0.00241f
C7982 a_4516_18884# a_4964_18884# 0.01328f
C7983 a_48321_23208# VPWR 1.23563f
C7984 a_38340_21327# a_38676_20452# 0.02511f
C7985 _459_.CLK a_33483_29535# 0.02343f
C7986 _304_.B _267_.ZN 0.00425f
C7987 _355_.C a_23084_28248# 0.0144f
C7988 a_29716_31048# VPWR 0.20777f
C7989 a_53660_15704# a_54244_15748# 0.01675f
C7990 a_59396_11044# VPWR 0.20622f
C7991 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN rst_n 0.0023f
C7992 a_56516_26344# a_56720_26344# 0.03324f
C7993 _478_.D _424_.A1 0.00481f
C7994 a_17168_27165# VPWR 0.18702f
C7995 a_65220_15748# a_65308_15704# 0.28563f
C7996 _304_.B _390_.ZN 0.19793f
C7997 _330_.A1 _448_.D 0.67136f
C7998 VPWR uio_oe[4] 0.30805f
C7999 a_36996_26344# a_36996_25156# 0.05841f
C8000 a_4156_27815# VPWR 0.3269f
C8001 a_31484_2727# a_31844_2824# 0.08717f
C8002 _282_.ZN a_47297_25596# 0.01609f
C8003 a_25012_31048# uio_out[2] 0.00726f
C8004 _457_.D a_25008_25597# 0.03113f
C8005 a_45128_26031# VPWR 0.1863f
C8006 a_60964_9476# a_61052_9432# 0.28563f
C8007 _397_.A1 _284_.A2 0.07317f
C8008 _325_.A2 a_40580_20072# 0.00861f
C8009 a_4516_7908# a_4604_7864# 0.28563f
C8010 a_18604_20408# a_19052_20408# 0.0131f
C8011 a_20756_20452# a_20396_20408# 0.08717f
C8012 _427_.B1 a_52452_21236# 0.46374f
C8013 a_8996_31048# a_9084_29383# 0.0027f
C8014 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I a_61724_15271# 0.0019f
C8015 a_3708_30951# a_4068_31048# 0.08717f
C8016 _350_.A1 _363_.Z 0.05346f
C8017 _229_.I _256_.A2 0.06365f
C8018 _397_.A2 a_47600_27912# 0.01308f
C8019 a_61500_17272# a_61388_16839# 0.02634f
C8020 a_8188_1592# VPWR 0.3582f
C8021 a_25884_1592# a_26020_1256# 0.00168f
C8022 a_57156_12612# a_57244_12568# 0.28563f
C8023 _459_.CLK a_18828_25112# 0.00189f
C8024 a_53212_12568# a_53660_12568# 0.01288f
C8025 _281_.ZN _476_.Q 0.59899f
C8026 _371_.ZN _459_.CLK 0.07401f
C8027 a_24452_24776# a_24428_23544# 0.0016f
C8028 _350_.A1 a_31396_31048# 0.01343f
C8029 a_63404_20408# VPWR 0.33437f
C8030 a_57020_1159# VPWR 0.33328f
C8031 _304_.B a_55228_28248# 0.01719f
C8032 a_62844_1159# a_62756_1256# 0.28563f
C8033 a_53684_12232# a_53660_11000# 0.0016f
C8034 a_57492_12232# a_57604_11044# 0.02666f
C8035 a_34980_1636# a_34620_1592# 0.08707f
C8036 a_34448_25597# a_35740_25112# 0.00486f
C8037 a_65756_18840# VPWR 0.34838f
C8038 _287_.A1 _358_.A3 0.0017f
C8039 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN a_61612_20408# 0.0053f
C8040 _246_.B2 _245_.Z 0.06775f
C8041 a_41140_27912# a_42148_27912# 0.00196f
C8042 _460_.Q _452_.CLK 0.71757f
C8043 a_67660_10567# a_68020_10664# 0.08717f
C8044 a_22748_1159# a_23196_1159# 0.0131f
C8045 a_53684_10664# a_54132_10664# 0.01328f
C8046 _371_.A2 _355_.B 0.00133f
C8047 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_55252_25156# 0.03524f
C8048 _304_.A1 _226_.ZN 0.34726f
C8049 _427_.B2 a_51108_21640# 0.00207f
C8050 _358_.A3 a_31932_26247# 0.01835f
C8051 a_27476_22020# VPWR 0.21518f
C8052 a_46356_24072# a_46984_23588# 0.00899f
C8053 _478_.D a_54804_23588# 0.00627f
C8054 _398_.C a_51332_24372# 0.07335f
C8055 a_19076_31048# a_18816_29931# 0.00187f
C8056 a_52676_2824# a_52764_1159# 0.0027f
C8057 a_58388_13800# VPWR 0.23551f
C8058 a_25348_21640# a_25796_21640# 0.01328f
C8059 a_37084_2727# VPWR 0.31143f
C8060 a_34308_18884# a_33948_18840# 0.08663f
C8061 _251_.A1 a_65072_29860# 0.00129f
C8062 a_1020_26247# a_932_26344# 0.28563f
C8063 _267_.ZN VPWR 0.67103f
C8064 _352_.A2 a_28036_26724# 0.00827f
C8065 a_1828_15368# a_2276_15368# 0.01328f
C8066 _438_.A2 _432_.ZN 0.00133f
C8067 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I VPWR 1.29622f
C8068 a_13700_29860# VPWR 0.20823f
C8069 a_3708_15271# a_3620_15368# 0.28563f
C8070 _350_.A2 a_31964_28292# 0.02456f
C8071 a_65980_11000# VPWR 0.36386f
C8072 a_24540_23111# VPWR 0.31547f
C8073 _231_.ZN a_59260_23544# 0.03631f
C8074 clkbuf_1_0__f_clk.I _399_.A2 0.00112f
C8075 _390_.ZN VPWR 0.66485f
C8076 _304_.A1 _300_.ZN 0.0867f
C8077 a_67100_17272# a_67012_15748# 0.00151f
C8078 a_64212_23208# a_64660_23208# 0.01328f
C8079 _325_.ZN a_42896_18504# 0.0482f
C8080 a_54444_26680# a_54892_26680# 0.01255f
C8081 a_42908_2727# a_42820_2824# 0.28563f
C8082 a_62980_17316# a_63428_17316# 0.01328f
C8083 _452_.CLK a_34304_24029# 0.02285f
C8084 a_29563_29535# a_29856_29123# 0.49319f
C8085 a_64524_16839# a_64884_16936# 0.08674f
C8086 _246_.B2 _252_.B 0.25028f
C8087 a_15244_23544# a_15692_23544# 0.01288f
C8088 a_66204_9432# a_66652_9432# 0.0131f
C8089 a_19188_23588# a_19276_23544# 0.28563f
C8090 a_23780_1256# a_24228_1256# 0.01328f
C8091 a_4068_25156# a_4156_25112# 0.28563f
C8092 a_64412_6296# a_64412_5863# 0.05841f
C8093 a_1020_5863# a_1468_5863# 0.0131f
C8094 _267_.A2 a_56484_29480# 0.0186f
C8095 a_67548_7864# a_67996_7864# 0.012f
C8096 a_2812_2727# a_3260_2727# 0.0131f
C8097 a_1916_4295# a_2364_4295# 0.0131f
C8098 a_65308_4728# a_65308_4295# 0.05841f
C8099 a_52876_13703# a_53324_13703# 0.01288f
C8100 _281_.ZN a_50084_24328# 0.1962f
C8101 _337_.A3 _371_.A1 0.07262f
C8102 a_35092_16936# a_35068_15271# 0.00134f
C8103 a_66876_14136# a_66764_13703# 0.02634f
C8104 _359_.B a_39300_29480# 0.00374f
C8105 _355_.C a_23060_26724# 0.01583f
C8106 _350_.A1 a_29371_30644# 0.00957f
C8107 _424_.B2 a_51620_19911# 0.03355f
C8108 a_18716_30951# a_18628_31048# 0.28563f
C8109 a_14236_29383# a_14684_29383# 0.0131f
C8110 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN 0.02591f
C8111 _452_.CLK a_36436_18504# 0.00737f
C8112 a_21988_1636# VPWR 0.2085f
C8113 a_18816_29931# a_19372_30345# 0.8399f
C8114 a_5724_30951# a_6172_30951# 0.01255f
C8115 _260_.ZN _305_.A2 0.0718f
C8116 a_50748_12568# a_50636_12135# 0.02634f
C8117 _474_.CLK a_52408_19759# 0.00603f
C8118 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I 0.00318f
C8119 a_55228_28248# VPWR 0.29679f
C8120 _459_.CLK a_16164_29480# 0.00204f
C8121 _355_.ZN a_28260_23208# 0.00235f
C8122 a_63516_15271# a_63428_15368# 0.28563f
C8123 _384_.ZN _281_.A1 0.00497f
C8124 a_48060_11000# a_48508_11000# 0.01288f
C8125 a_52004_11044# a_52092_11000# 0.28563f
C8126 a_39124_16936# a_39572_16936# 0.01328f
C8127 a_33860_18504# VPWR 0.21375f
C8128 a_41476_1636# a_41924_1636# 0.01328f
C8129 a_56236_24679# vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN 0.01518f
C8130 a_65308_15704# a_65444_15368# 0.00168f
C8131 a_3620_26724# a_4068_26724# 0.01328f
C8132 a_1828_26724# a_1468_26680# 0.08717f
C8133 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN 0.03773f
C8134 a_49496_30345# VPWR 0.19192f
C8135 a_33483_29535# uo_out[7] 0.00542f
C8136 _371_.ZN _371_.A3 0.07212f
C8137 _243_.B2 a_59172_27912# 0.00323f
C8138 _256_.A2 rst_n 0.0089f
C8139 _324_.C vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I 0.04097f
C8140 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I 0.00251f
C8141 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_63404_23111# 0.00533f
C8142 a_50436_30689# _275_.A2 0.00702f
C8143 a_47524_12612# VPWR 0.20348f
C8144 a_59484_2727# VPWR 0.31143f
C8145 a_35816_21192# _319_.A3 0.24626f
C8146 _416_.A1 _452_.CLK 0.12408f
C8147 a_15604_26344# a_16052_26344# 0.01328f
C8148 a_66092_18407# a_66004_18504# 0.28563f
C8149 a_3620_2824# a_4068_2824# 0.01328f
C8150 a_58948_26344# _231_.ZN 0.00598f
C8151 a_3172_20072# VPWR 0.20993f
C8152 a_56684_17272# a_57132_17272# 0.01255f
C8153 a_1468_29383# a_1828_29480# 0.08717f
C8154 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_54780_26247# 0.00174f
C8155 a_60268_10567# VPWR 0.31389f
C8156 a_35723_20569# _448_.D 0.00455f
C8157 _365_.ZN VPWR 1.10493f
C8158 a_29356_21976# a_29244_21543# 0.02634f
C8159 a_39772_15271# a_40132_15368# 0.08717f
C8160 a_22212_23208# VPWR 0.20862f
C8161 a_57940_18884# VPWR 0.21986f
C8162 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN 0.00226f
C8163 _256_.A2 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN 0.13777f
C8164 _452_.CLK a_34080_22461# 0.00354f
C8165 a_3260_28248# a_3708_28248# 0.0131f
C8166 _251_.A1 _274_.A2 0.04573f
C8167 a_53660_2727# a_54244_2824# 0.01675f
C8168 a_31172_16936# a_31172_15748# 0.05841f
C8169 _304_.B a_54892_26680# 0.00277f
C8170 a_19724_23544# a_19636_22020# 0.00151f
C8171 _274_.A3 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN 0.04474f
C8172 a_22996_23588# a_23084_23544# 0.28563f
C8173 _350_.A1 uo_out[3] 0.15563f
C8174 a_2276_31048# VPWR 0.20634f
C8175 a_1828_1256# VPWR 0.20348f
C8176 _371_.ZN uo_out[7] 0.00543f
C8177 a_17844_25156# a_17932_25112# 0.28563f
C8178 a_21428_25156# a_21876_25156# 0.01328f
C8179 _386_.A4 _393_.A1 0.04965f
C8180 _383_.ZN _390_.ZN 0.02098f
C8181 _476_.Q a_50660_20452# 0.00108f
C8182 _349_.A4 a_25884_27815# 0.00169f
C8183 a_31732_20452# a_31372_20408# 0.08717f
C8184 a_50188_13703# a_50100_13800# 0.28563f
C8185 a_46068_16936# a_46044_15271# 0.00144f
C8186 a_63740_14136# a_63764_13800# 0.00172f
C8187 _427_.A2 _424_.ZN 0.00162f
C8188 _384_.A1 clk 0.0107f
C8189 a_22636_30951# a_23084_30951# 0.012f
C8190 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN 0.0138f
C8191 a_36972_16839# a_36884_16936# 0.28563f
C8192 a_54040_22366# VPWR 0.50875f
C8193 _311_.A2 _313_.ZN 0.76929f
C8194 a_28124_1592# VPWR 0.29679f
C8195 _422_.ZN a_52452_21236# 0.17044f
C8196 a_67324_12568# a_67772_12568# 0.01288f
C8197 a_57692_12568# a_57580_12135# 0.02634f
C8198 a_18816_29931# a_20003_29611# 0.01007f
C8199 _337_.ZN a_29680_26724# 0.00293f
C8200 a_4516_1636# a_4964_1636# 0.01328f
C8201 _460_.Q a_34448_25597# 0.23215f
C8202 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN 0.00414f
C8203 a_1916_11000# a_1916_10567# 0.05841f
C8204 a_55364_11044# a_55004_11000# 0.08707f
C8205 a_57940_12232# a_58028_10567# 0.00151f
C8206 _324_.C vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.00423f
C8207 vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I 0.51221f
C8208 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN a_61636_18504# 0.07278f
C8209 a_45148_1159# a_45596_1159# 0.0131f
C8210 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_62284_23544# 0.0546f
C8211 a_4068_27912# a_4068_26724# 0.05841f
C8212 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN 0.0011f
C8213 vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I 0.66565f
C8214 a_54804_20072# a_54780_18840# 0.0016f
C8215 a_62980_18884# a_63428_18884# 0.01328f
C8216 a_47724_18840# VPWR 0.31595f
C8217 a_19052_20408# VPWR 0.32276f
C8218 a_54040_22366# a_54108_21543# 0.01908f
C8219 _355_.C a_23084_25112# 0.00613f
C8220 a_53660_12568# VPWR 0.31389f
C8221 a_2276_15748# a_2724_15748# 0.01328f
C8222 a_10876_2727# a_11012_1636# 0.00154f
C8223 a_12892_29383# a_12804_29480# 0.28563f
C8224 a_49092_15368# a_49764_15368# 0.00347f
C8225 _251_.A1 a_56260_31048# 0.00189f
C8226 a_54132_10664# VPWR 0.20614f
C8227 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN 0.01222f
C8228 a_56684_18407# a_57044_18504# 0.08674f
C8229 a_1020_8999# a_1380_9096# 0.08717f
C8230 a_53212_27815# a_53572_27912# 0.0869f
C8231 a_1916_7431# a_2276_7528# 0.08717f
C8232 a_51196_15271# a_51108_15368# 0.28563f
C8233 a_2812_5863# a_3172_5960# 0.08717f
C8234 a_3708_4295# a_4068_4392# 0.08717f
C8235 a_52540_15271# a_52988_15271# 0.0131f
C8236 a_44744_26355# a_45128_26031# 1.16391f
C8237 a_2276_15368# VPWR 0.20634f
C8238 a_58364_25112# clk 0.00333f
C8239 a_53548_24679# a_52852_24372# 0.00604f
C8240 a_16140_21976# a_16588_21976# 0.01288f
C8241 a_38576_22504# a_38968_22504# 0.00629f
C8242 a_20084_22020# a_20172_21976# 0.28563f
C8243 _355_.C a_25796_27912# 0.00773f
C8244 a_65084_2727# a_64996_2824# 0.28563f
C8245 a_30812_15271# VPWR 0.30073f
C8246 a_33948_16839# a_34732_16839# 0.00443f
C8247 a_5052_17272# a_4964_15748# 0.00151f
C8248 a_49404_30951# a_49316_31048# 0.28563f
C8249 a_23532_23544# a_23444_22020# 0.00151f
C8250 a_54892_26680# VPWR 0.31547f
C8251 a_29856_29123# VPWR 0.50544f
C8252 _473_.Q a_47552_19715# 0.19413f
C8253 a_63428_17316# VPWR 0.20348f
C8254 _404_.A1 a_47172_27912# 0.00248f
C8255 a_30500_23208# a_30588_21543# 0.00151f
C8256 a_29804_23544# a_30388_23588# 0.01675f
C8257 a_45956_1256# a_46628_1256# 0.00347f
C8258 a_2364_4295# VPWR 0.30029f
C8259 a_24228_1256# VPWR 0.20348f
C8260 a_67996_7864# VPWR 0.35142f
C8261 a_25212_2727# a_25660_2727# 0.0131f
C8262 a_14684_29383# VPWR 0.29679f
C8263 a_57692_14136# a_57604_12612# 0.00151f
C8264 a_60716_13703# a_61076_13800# 0.08707f
C8265 a_46628_13800# a_47076_13800# 0.01328f
C8266 a_6172_30951# VPWR 0.32306f
C8267 _311_.A2 _316_.ZN 0.00351f
C8268 a_47500_16839# a_47860_16936# 0.08707f
C8269 _480_.Q a_43664_29535# 0.00159f
C8270 _330_.A1 _424_.A2 0.04243f
C8271 a_18716_23111# a_18740_22020# 0.0016f
C8272 a_932_9476# a_1020_9432# 0.28563f
C8273 a_50996_10664# a_50972_9432# 0.0016f
C8274 a_21052_26031# a_21396_26399# 0.00275f
C8275 a_39572_16936# VPWR 0.20637f
C8276 a_41924_1636# VPWR 0.21436f
C8277 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN VPWR 0.7944f
C8278 a_6620_1159# a_6532_1256# 0.28563f
C8279 a_54556_12568# a_54580_12232# 0.00172f
C8280 _268_.A2 _268_.A1 2.08974f
C8281 _452_.CLK a_41776_18504# 0.00156f
C8282 a_19276_25112# a_19164_24679# 0.02634f
C8283 a_2364_29816# a_2812_29816# 0.01288f
C8284 a_6308_29860# a_6396_29816# 0.28563f
C8285 a_5052_15704# a_4964_14180# 0.00151f
C8286 a_32516_17316# a_32964_17316# 0.01328f
C8287 _275_.A2 VPWR 0.92432f
C8288 a_62172_15271# a_62308_14180# 0.00154f
C8289 a_61860_11044# a_62308_11044# 0.01328f
C8290 a_4068_2824# VPWR 0.22189f
C8291 a_52452_11044# a_52428_10567# 0.00172f
C8292 a_48508_11000# a_48508_10567# 0.05841f
C8293 _251_.A1 a_62396_27815# 0.03252f
C8294 a_51556_1636# a_51644_1592# 0.28563f
C8295 a_23868_1592# a_23868_1159# 0.05841f
C8296 a_57132_17272# VPWR 0.33195f
C8297 _337_.ZN a_28756_25940# 0.00181f
C8298 a_32068_20072# a_32068_18884# 0.05841f
C8299 _371_.A1 a_29828_26344# 0.00239f
C8300 _424_.ZN a_52228_19368# 0.42528f
C8301 _324_.B _328_.A2 0.13226f
C8302 a_3708_23111# a_4156_23111# 0.0131f
C8303 a_51308_18407# a_51668_18504# 0.08717f
C8304 _336_.A1 a_29176_25273# 0.00151f
C8305 a_45060_2824# a_45060_1636# 0.05841f
C8306 a_41252_2824# a_41116_1592# 0.00154f
C8307 a_53012_18504# a_53100_16839# 0.00151f
C8308 a_50324_18504# VPWR 0.25458f
C8309 a_21876_25156# VPWR 0.20983f
C8310 _452_.D a_41432_17801# 0.00911f
C8311 a_4068_27912# a_4852_27912# 0.00276f
C8312 a_30028_20408# VPWR 0.31605f
C8313 a_19500_27815# a_19860_27912# 0.08674f
C8314 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN _324_.C 0.00261f
C8315 a_23084_30951# VPWR 0.33606f
C8316 vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN VPWR 0.89309f
C8317 _303_.ZN _325_.B 0.01939f
C8318 _393_.A1 a_45396_28292# 0.00462f
C8319 a_67772_12568# VPWR 0.33516f
C8320 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN _249_.A2 0.73848f
C8321 a_39100_15704# a_39236_15368# 0.00168f
C8322 a_26020_2824# a_26468_2824# 0.01328f
C8323 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN a_58924_14136# 0.00378f
C8324 vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN 0.00215f
C8325 a_56596_17316# vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I 0.00803f
C8326 a_18628_21640# a_18516_20452# 0.02666f
C8327 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN a_57492_18884# 0.07232f
C8328 vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN 0.00102f
C8329 _251_.A1 a_58340_29860# 0.00173f
C8330 a_38764_20408# a_38876_19975# 0.02634f
C8331 a_2724_15748# VPWR 0.20782f
C8332 a_49764_15368# VPWR 0.23042f
C8333 _474_.CLK a_54420_21976# 0.00556f
C8334 a_23444_22020# a_23084_21976# 0.08707f
C8335 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_56388_25940# 0.00172f
C8336 a_47689_25156# VPWR 0.00561f
C8337 a_52988_15271# VPWR 0.3577f
C8338 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.01285f
C8339 a_47076_14180# a_47524_14180# 0.01328f
C8340 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN a_55228_27815# 0.00323f
C8341 a_34844_17272# a_34756_15748# 0.00151f
C8342 _452_.CLK a_35204_17316# 0.00146f
C8343 a_34732_16839# VPWR 0.34674f
C8344 a_24196_31048# a_22996_31048# 0.00154f
C8345 a_46628_1256# VPWR 0.22423f
C8346 _230_.I _243_.A1 0.06023f
C8347 a_23084_30951# a_24564_31048# 0.00188f
C8348 a_32848_29123# _223_.ZN 0.00497f
C8349 a_4068_13800# a_4068_12612# 0.05841f
C8350 a_61500_14136# a_61412_12612# 0.00151f
C8351 _358_.A2 a_30388_25156# 0.00733f
C8352 a_50748_20408# a_49896_18909# 0.00106f
C8353 a_50300_20408# a_50384_19204# 0.00131f
C8354 _362_.B a_35292_26247# 0.00156f
C8355 _363_.Z _290_.ZN 0.06404f
C8356 a_17396_23208# a_17396_22020# 0.05841f
C8357 a_32964_17316# VPWR 0.20348f
C8358 _417_.A2 _427_.B2 0.20222f
C8359 a_17596_1159# a_17956_1256# 0.08717f
C8360 _371_.A1 a_32580_27912# 0.00194f
C8361 a_61612_12135# a_62060_12135# 0.01288f
C8362 a_47612_12135# a_47972_12232# 0.08717f
C8363 vgaringosc.workerclkbuff_notouch_.I a_48708_29816# 0.02589f
C8364 a_48060_1592# VPWR 0.30141f
C8365 a_31372_23544# a_31484_23111# 0.02634f
C8366 a_10788_29480# a_11236_29480# 0.01328f
C8367 a_10652_1592# a_11100_1592# 0.01288f
C8368 a_14596_1636# a_14684_1592# 0.28563f
C8369 VPWR ena 0.33188f
C8370 _331_.ZN a_41188_18840# 0.02523f
C8371 _428_.Z _475_.Q 0.00132f
C8372 a_55252_26724# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.00875f
C8373 a_9668_29860# a_9308_29816# 0.08707f
C8374 a_55364_15368# a_55364_14180# 0.05841f
C8375 _304_.B _325_.A1 0.05925f
C8376 a_55452_11000# a_55564_10567# 0.02634f
C8377 a_47972_31048# a_48420_31048# 0.01328f
C8378 a_59396_11044# a_59372_10567# 0.00172f
C8379 a_26468_2824# VPWR 0.21447f
C8380 _451_.Q a_37408_18504# 0.00269f
C8381 a_30812_1592# a_30812_1159# 0.05841f
C8382 _459_.CLK a_17484_27815# 0.02224f
C8383 a_37968_31048# uo_out[2] 0.00128f
C8384 a_2812_23111# a_2724_23208# 0.28563f
C8385 a_15692_24679# a_15604_24776# 0.28563f
C8386 a_24092_24679# a_24540_24679# 0.01288f
C8387 a_2724_9096# a_3172_9096# 0.01328f
C8388 a_67548_1159# a_67996_1159# 0.01222f
C8389 a_54244_15748# a_54332_15704# 0.28563f
C8390 a_32156_19975# a_32604_19975# 0.0131f
C8391 a_4940_5863# a_4964_4772# 0.0016f
C8392 a_4852_5960# a_5300_5960# 0.01328f
C8393 a_47524_14180# VPWR 0.20952f
C8394 a_3620_7528# a_4068_7528# 0.01328f
C8395 a_64324_4392# a_64772_4392# 0.01328f
C8396 a_2812_18407# a_3172_18504# 0.08717f
C8397 a_33500_18407# a_33948_18407# 0.0131f
C8398 _247_.ZN _243_.ZN 0.25392f
C8399 _438_.A2 _260_.A2 0.05592f
C8400 a_55252_25156# a_55700_25156# 0.01328f
C8401 a_36636_15704# a_37084_15704# 0.01288f
C8402 a_62060_12135# VPWR 0.31547f
C8403 a_11236_29480# VPWR 0.21187f
C8404 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_64772_26344# 0.00546f
C8405 a_48420_31048# VPWR 0.20938f
C8406 _340_.ZN a_24100_29480# 0.00427f
C8407 _324_.C vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN 0.11832f
C8408 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN a_64884_26724# 0.00225f
C8409 _358_.A3 a_34308_26344# 0.10518f
C8410 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN VPWR 0.96077f
C8411 a_24540_24679# VPWR 0.32114f
C8412 a_51780_15748# a_51644_15271# 0.00168f
C8413 a_47836_15704# a_47836_15271# 0.05841f
C8414 a_61972_23208# vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN 0.0356f
C8415 a_4068_7528# VPWR 0.22146f
C8416 _275_.ZN a_51050_29480# 0.02622f
C8417 a_34396_21543# _319_.ZN 0.00193f
C8418 a_64772_4392# VPWR 0.20727f
C8419 a_45036_28248# a_45484_28248# 0.01222f
C8420 a_55700_25156# VPWR 0.21119f
C8421 a_37084_15704# VPWR 0.3289f
C8422 _379_.A2 uio_out[4] 0.00117f
C8423 a_41099_26841# a_41344_27209# 0.00232f
C8424 a_29788_30345# uo_out[6] 0.00152f
C8425 a_52652_18407# a_53100_18407# 0.0131f
C8426 a_29804_21976# a_30388_22020# 0.01675f
C8427 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN a_59620_23208# 0.00137f
C8428 _436_.ZN a_40565_24394# 0.00616f
C8429 a_53100_18407# VPWR 0.329f
C8430 a_67236_15368# a_67236_14180# 0.05841f
C8431 _459_.CLK a_27228_26247# 0.05214f
C8432 _359_.ZN a_34516_25940# 0.00922f
C8433 _455_.Q a_23780_26344# 0.0025f
C8434 _399_.A1 VPWR 0.55595f
C8435 a_4604_1592# a_4740_1256# 0.00168f
C8436 a_47612_2727# a_48060_2727# 0.0131f
C8437 a_52340_13800# a_52452_12612# 0.02666f
C8438 a_932_12612# a_1380_12612# 0.01328f
C8439 a_48508_18407# a_48644_17316# 0.00154f
C8440 _324_.C a_59948_30352# 0.00271f
C8441 a_33312_28776# uo_out[7] 0.0013f
C8442 _231_.ZN a_57916_25112# 0.00122f
C8443 a_46492_17272# a_46604_16839# 0.02634f
C8444 a_50436_17316# a_50412_16839# 0.00172f
C8445 _325_.A2 a_43888_19204# 0.01863f
C8446 a_24452_23208# a_24340_22020# 0.02666f
C8447 a_44812_17272# VPWR 0.29679f
C8448 a_61724_1592# VPWR 0.32824f
C8449 a_29020_1159# a_28932_1256# 0.28563f
C8450 a_17956_1636# a_17596_1592# 0.08707f
C8451 _346_.A2 a_23420_26247# 0.02316f
C8452 a_58924_12135# a_58836_12232# 0.28563f
C8453 a_41216_23208# VPWR 0.0143f
C8454 _474_.CLK a_52116_18504# 0.00546f
C8455 a_17484_21543# VPWR 0.29719f
C8456 a_60401_30300# VPWR 0.47715f
C8457 a_16028_29816# a_16612_29860# 0.01675f
C8458 _448_.Q a_39669_21236# 0.00449f
C8459 _304_.B _327_.A2 0.03438f
C8460 a_44364_17272# a_44812_17272# 0.01255f
C8461 _237_.A1 a_58709_29076# 0.00927f
C8462 _325_.A1 VPWR 2.7364f
C8463 a_66340_11044# a_66316_10567# 0.00172f
C8464 a_48508_10567# a_49292_10567# 0.00443f
C8465 a_48868_2824# VPWR 0.2062f
C8466 a_61276_1592# a_61724_1592# 0.01288f
C8467 _430_.ZN _301_.A1 0.63193f
C8468 a_22748_23111# a_23108_23208# 0.08707f
C8469 _251_.A1 a_62756_27912# 0.02975f
C8470 a_1380_23208# a_1828_23208# 0.01328f
C8471 a_27172_24328# a_27924_24776# 0.09971f
C8472 a_51780_9476# VPWR 0.20677f
C8473 a_54556_21543# VPWR 0.32433f
C8474 a_25012_31048# VPWR 0.20513f
C8475 a_17036_21543# a_17484_21543# 0.0131f
C8476 a_54556_14136# VPWR 0.31389f
C8477 _325_.A1 a_41012_23208# 0.00275f
C8478 _474_.Q a_47948_23111# 0.05577f
C8479 _452_.CLK a_33164_24679# 0.00625f
C8480 _362_.B _437_.A1 0.00364f
C8481 a_6756_29860# a_6620_29383# 0.00168f
C8482 a_2812_29816# a_2812_29383# 0.05841f
C8483 a_43940_15748# a_43580_15704# 0.08707f
C8484 a_55924_12232# VPWR 0.20622f
C8485 _397_.A1 _419_.A4 0.04051f
C8486 a_48420_2824# a_48868_2824# 0.01328f
C8487 a_20396_27815# a_21044_27508# 0.00223f
C8488 a_57156_27912# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.04067f
C8489 a_52228_19368# a_52436_18884# 0.02745f
C8490 a_49112_29885# a_49496_30345# 1.16391f
C8491 _441_.A2 _439_.ZN 0.01736f
C8492 a_30240_24776# VPWR 1.09923f
C8493 a_61636_20072# VPWR 0.20812f
C8494 _371_.ZN _340_.A2 0.04479f
C8495 _459_.Q a_35140_26680# 0.00811f
C8496 _416_.ZN a_46268_18407# 0.00254f
C8497 a_9084_2727# a_8996_2824# 0.28563f
C8498 _395_.A2 _412_.B2 0.2462f
C8499 a_50884_15748# VPWR 0.21255f
C8500 a_54108_21543# a_54556_21543# 0.01255f
C8501 _412_.A1 a_48384_26724# 0.04747f
C8502 _424_.B1 _395_.A3 0.04533f
C8503 a_25764_29977# VPWR 0.00258f
C8504 a_51332_9476# a_51780_9476# 0.01328f
C8505 a_49988_9476# a_49628_9432# 0.08717f
C8506 a_24564_31048# a_25012_31048# 0.01328f
C8507 a_57604_14180# a_57692_14136# 0.28563f
C8508 _452_.CLK _431_.A3 0.00715f
C8509 a_5052_14136# a_4940_13703# 0.02634f
C8510 a_54108_14136# a_54556_14136# 0.0131f
C8511 _287_.A1 uo_out[1] 0.00751f
C8512 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I 0.25671f
C8513 a_11548_1592# a_11684_1256# 0.00168f
C8514 a_59284_13800# a_59396_12612# 0.02666f
C8515 a_55476_13800# a_55452_12568# 0.0016f
C8516 a_58388_20452# VPWR 0.23732f
C8517 _395_.A1 a_51048_26680# 0.01209f
C8518 a_36548_26344# VPWR 0.20348f
C8519 _346_.A2 _346_.ZN 0.60797f
C8520 a_31396_23208# a_31284_22020# 0.02666f
C8521 a_2724_24776# a_2724_23588# 0.05841f
C8522 _355_.C _343_.A2 0.42649f
C8523 a_39996_1159# a_40356_1256# 0.08717f
C8524 a_11772_1159# VPWR 0.37894f
C8525 a_4852_9096# a_4964_7908# 0.02666f
C8526 a_55476_12232# a_55924_12232# 0.01328f
C8527 a_24452_1636# a_24900_1636# 0.01328f
C8528 vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I 0.00117f
C8529 a_14708_21640# VPWR 0.22176f
C8530 _327_.A2 VPWR 1.8463f
C8531 a_59260_26680# _251_.ZN 0.00963f
C8532 a_51780_17316# a_51420_17272# 0.08707f
C8533 a_45820_10567# a_45732_10664# 0.28563f
C8534 _238_.I a_60852_28292# 0.02459f
C8535 a_35292_30951# _365_.ZN 0.00169f
C8536 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I a_52415_31220# 0.00232f
C8537 a_64300_23111# VPWR 0.29893f
C8538 _459_.CLK _336_.A2 0.10817f
C8539 _268_.A2 _474_.CLK 1.16666f
C8540 a_33724_23111# a_33636_23208# 0.28563f
C8541 clkbuf_1_0__f_clk.I _399_.ZN 0.10808f
C8542 a_62756_9476# VPWR 0.20595f
C8543 a_3260_23544# VPWR 0.30487f
C8544 a_54420_21976# a_55208_22505# 0.02112f
C8545 a_15692_21543# a_16052_21640# 0.08717f
C8546 a_61188_20072# a_61636_20072# 0.01328f
C8547 a_59260_23544# clk 0.00531f
C8548 a_3260_6296# VPWR 0.30487f
C8549 _350_.A1 _294_.ZN 0.02168f
C8550 a_5052_3160# VPWR 0.34934f
C8551 _325_.A1 a_40452_22504# 0.00491f
C8552 a_2364_13703# VPWR 0.30029f
C8553 a_55252_26724# a_54892_26680# 0.0869f
C8554 _264_.B _304_.A1 0.00324f
C8555 _294_.A2 a_30388_28776# 0.01171f
C8556 _474_.D a_51252_19001# 0.00159f
C8557 _452_.CLK a_34396_18840# 0.01266f
C8558 _424_.A2 a_47483_20569# 0.00426f
C8559 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN a_58500_21640# 0.00328f
C8560 a_37444_25156# VPWR 0.20924f
C8561 a_50436_15748# a_50884_15748# 0.01328f
C8562 a_46852_15748# a_46940_15704# 0.28563f
C8563 a_45284_11044# VPWR 0.22176f
C8564 _435_.ZN a_39760_23588# 0.0063f
C8565 a_66540_19975# a_66900_20072# 0.0869f
C8566 _474_.CLK a_54892_18407# 0.00211f
C8567 _237_.A1 a_60909_30600# 0.02482f
C8568 a_32156_18840# VPWR 0.29679f
C8569 a_15244_26247# VPWR 0.29679f
C8570 _359_.B vgaringosc.workerclkbuff_notouch_.I 0.11724f
C8571 a_43804_30951# a_43828_29860# 0.0016f
C8572 a_59260_23111# VPWR 0.29802f
C8573 a_20060_2727# a_20420_2824# 0.08717f
C8574 _293_.A2 uo_out[1] 1.91637f
C8575 a_1916_9432# a_1916_8999# 0.05841f
C8576 _330_.A2 a_39236_17316# 0.07238f
C8577 _304_.B a_45232_25987# 0.03068f
C8578 a_28012_21976# a_27924_20452# 0.00151f
C8579 _459_.Q _460_.D 0.20773f
C8580 a_51644_14136# a_51532_13703# 0.02634f
C8581 a_62308_14180# a_62396_14136# 0.28563f
C8582 a_14708_20452# a_15156_20452# 0.01328f
C8583 _447_.Q a_37196_23544# 0.02725f
C8584 _459_.CLK _346_.A2 0.86815f
C8585 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN VPWR 0.71289f
C8586 _250_.ZN _250_.C 0.21206f
C8587 a_66228_13800# a_66340_12612# 0.02666f
C8588 _397_.A1 a_48820_28292# 0.00157f
C8589 a_49852_12568# a_50300_12568# 0.01288f
C8590 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I a_58164_18504# 0.00339f
C8591 _313_.ZN a_36860_23111# 0.00598f
C8592 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN VPWR 0.99694f
C8593 a_20420_24776# a_20532_23588# 0.02666f
C8594 a_21204_31048# _346_.B 0.00121f
C8595 _416_.A1 a_45820_18840# 0.00246f
C8596 _335_.ZN a_36420_28776# 0.00371f
C8597 _379_.A2 a_21740_29383# 0.00518f
C8598 a_57940_20452# a_58388_20452# 0.01328f
C8599 a_34172_1159# VPWR 0.30352f
C8600 a_51420_1159# a_51332_1256# 0.28563f
C8601 a_31620_1636# a_31260_1592# 0.08663f
C8602 a_60268_12135# a_60292_11044# 0.0016f
C8603 _296_.ZN _462_.D 0.01586f
C8604 a_46984_23588# a_47948_23111# 0.02974f
C8605 a_18028_28777# a_18372_28409# 0.00275f
C8606 a_45508_31048# a_45012_29816# 0.00123f
C8607 a_37084_21543# VPWR 0.31591f
C8608 _302_.Z a_42784_22504# 0.00353f
C8609 a_36100_26344# a_36548_26344# 0.01328f
C8610 a_63852_23544# VPWR 0.29679f
C8611 _452_.Q _324_.B 0.05189f
C8612 a_56460_10567# a_57044_10664# 0.01675f
C8613 a_2724_10664# a_3172_10664# 0.01328f
C8614 _381_.Z a_50120_26476# 0.03756f
C8615 _395_.A1 _381_.A2 0.04538f
C8616 _267_.A1 a_55588_28292# 0.0146f
C8617 a_11324_1159# a_11772_1159# 0.0131f
C8618 a_4940_18407# a_4964_17316# 0.0016f
C8619 a_49448_20072# VPWR 0.61855f
C8620 VPWR uio_out[2] 0.08141f
C8621 a_4156_21976# VPWR 0.30552f
C8622 a_32292_23208# a_32740_23208# 0.01328f
C8623 _402_.A1 a_43940_27912# 0.02975f
C8624 a_2276_18884# a_2364_18840# 0.28563f
C8625 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN 0.00155f
C8626 a_26132_23588# VPWR 0.21395f
C8627 a_27004_21543# a_26916_21640# 0.28563f
C8628 _386_.ZN a_47525_29480# 0.04111f
C8629 a_41252_2824# a_41340_1159# 0.0027f
C8630 a_52920_22760# VPWR 0.51559f
C8631 a_14236_2727# VPWR 0.31143f
C8632 a_63852_13703# VPWR 0.31556f
C8633 a_16164_29480# a_16140_28248# 0.0016f
C8634 _218_.ZN _395_.A3 0.04059f
C8635 _399_.A1 a_51240_23340# 0.00608f
C8636 _355_.C a_22636_28248# 0.03264f
C8637 _459_.CLK a_32476_29167# 0.01498f
C8638 a_39772_26247# _436_.ZN 0.00139f
C8639 a_67861_31220# VPWR 0.00437f
C8640 _495_.I vgaringosc.workerclkbuff_notouch_.I 0.01485f
C8641 a_58948_11044# VPWR 0.20622f
C8642 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN 0.00552f
C8643 a_56516_26344# a_56368_26344# 0.00128f
C8644 _371_.A3 _336_.A2 0.00494f
C8645 a_16240_26795# VPWR 1.09532f
C8646 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN 0.01949f
C8647 a_17372_30951# a_17508_29860# 0.00154f
C8648 a_65220_15748# a_64860_15704# 0.08717f
C8649 _330_.A1 a_35716_20072# 0.00119f
C8650 _438_.A2 _311_.A2 0.21444f
C8651 a_3708_27815# VPWR 0.33374f
C8652 _265_.ZN a_43008_26795# 0.00346f
C8653 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I 0.00365f
C8654 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.18341f
C8655 a_63852_23111# a_64300_23111# 0.0131f
C8656 a_31484_2727# a_31396_2824# 0.28563f
C8657 _457_.D a_24080_25227# 0.28107f
C8658 _421_.A1 _279_.Z 0.00373f
C8659 a_24564_31048# uio_out[2] 0.00354f
C8660 a_45232_25987# VPWR 0.39609f
C8661 a_48888_19243# a_49492_18840# 0.49241f
C8662 a_2812_23544# a_3260_23544# 0.0131f
C8663 a_12356_1256# a_12804_1256# 0.01328f
C8664 a_1916_7864# a_2364_7864# 0.0131f
C8665 a_4516_7908# a_4156_7864# 0.08674f
C8666 _397_.A1 a_51048_26680# 0.00374f
C8667 a_60964_9476# a_60604_9432# 0.08717f
C8668 a_62308_9476# a_62756_9476# 0.01328f
C8669 _325_.A2 a_40132_20072# 0.00699f
C8670 _229_.I _238_.ZN 0.0153f
C8671 a_3708_4728# a_4156_4728# 0.0131f
C8672 a_18180_31048# a_18628_31048# 0.01328f
C8673 a_2812_6296# a_3260_6296# 0.0131f
C8674 a_1916_13703# a_2364_13703# 0.0131f
C8675 a_4604_3160# a_5052_3160# 0.01222f
C8676 _448_.Q _316_.A3 0.01134f
C8677 _316_.ZN _319_.ZN 0.00479f
C8678 a_59372_14136# a_59372_13703# 0.05841f
C8679 a_20308_20452# a_20396_20408# 0.28563f
C8680 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I a_61276_15271# 0.00606f
C8681 a_2812_29383# a_3260_29383# 0.0131f
C8682 a_3708_30951# a_3620_31048# 0.28563f
C8683 a_59955_30600# ui_in[3] 0.01621f
C8684 _397_.A2 a_47376_27912# 0.00344f
C8685 a_7740_1592# VPWR 0.3289f
C8686 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN 0.0058f
C8687 a_59732_13800# a_59820_12135# 0.00151f
C8688 a_3708_12568# a_3708_12135# 0.05841f
C8689 _459_.CLK a_18380_25112# 0.00189f
C8690 vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN 0.02902f
C8691 a_57156_12612# a_56796_12568# 0.08707f
C8692 _267_.A1 a_55588_27912# 0.00265f
C8693 a_27924_24776# a_27924_23588# 0.05841f
C8694 a_62396_1159# a_62756_1256# 0.08717f
C8695 a_56572_1159# VPWR 0.33158f
C8696 a_62060_20408# VPWR 0.32563f
C8697 a_36996_25156# a_37444_25156# 0.01328f
C8698 _350_.A1 a_30778_31048# 0.00188f
C8699 _416_.A1 _447_.Q 0.00198f
C8700 _402_.A1 a_48292_26369# 0.00175f
C8701 a_67212_12135# a_67236_11044# 0.0016f
C8702 a_65308_18840# VPWR 0.30377f
C8703 a_38116_1636# a_38564_1636# 0.01328f
C8704 a_34532_1636# a_34620_1592# 0.28563f
C8705 a_2724_16936# a_3172_16936# 0.01328f
C8706 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN a_61164_20408# 0.0016f
C8707 _441_.ZN a_39760_23588# 0.0096f
C8708 _246_.B2 a_59172_26724# 0.01596f
C8709 _474_.Q a_48529_22460# 0.00255f
C8710 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN 0.75003f
C8711 a_32964_18504# a_32964_17316# 0.05841f
C8712 a_62980_1636# a_62844_1159# 0.00168f
C8713 a_59036_1592# a_59036_1159# 0.05841f
C8714 a_67660_10567# a_67572_10664# 0.28563f
C8715 a_23780_2824# a_23780_1636# 0.05841f
C8716 a_19972_2824# a_19836_1592# 0.00154f
C8717 a_27028_22020# VPWR 0.23583f
C8718 _358_.A3 a_30724_26020# 0.18445f
C8719 _355_.C a_24952_29032# 0.02706f
C8720 _478_.D a_54356_23588# 0.00727f
C8721 a_31708_18840# a_32156_18840# 0.0131f
C8722 a_33860_18884# a_33948_18840# 0.28563f
C8723 a_13700_29860# uio_oe[2] 0.0058f
C8724 _441_.A2 _303_.ZN 0.02404f
C8725 a_36636_2727# VPWR 0.31143f
C8726 a_57940_13800# VPWR 0.21723f
C8727 a_14796_26247# a_15244_26247# 0.0131f
C8728 a_49740_29383# VPWR 0.32863f
C8729 _352_.A2 a_27588_26724# 0.00121f
C8730 a_57916_25112# a_58364_25112# 0.01222f
C8731 a_13252_29860# VPWR 0.20614f
C8732 a_56404_27208# VPWR 0.55961f
C8733 a_63540_16936# a_63428_15748# 0.02666f
C8734 a_65532_11000# VPWR 0.32454f
C8735 a_3260_15271# a_3620_15368# 0.08717f
C8736 _350_.A2 a_31516_28292# 0.02109f
C8737 a_24092_23111# VPWR 0.31547f
C8738 a_63852_23544# a_63852_23111# 0.05841f
C8739 a_48141_29480# VPWR 0.00658f
C8740 _349_.A4 _337_.A3 0.03648f
C8741 a_42236_2727# a_42820_2824# 0.01675f
C8742 a_64524_16839# a_64436_16936# 0.28563f
C8743 a_62620_18407# a_63068_18407# 0.0131f
C8744 a_61612_20408# a_61636_20072# 0.00172f
C8745 a_19188_23588# a_18828_23544# 0.08707f
C8746 a_1468_25112# a_1916_25112# 0.0131f
C8747 a_4068_25156# a_3708_25112# 0.08717f
C8748 a_55900_14136# a_55924_13800# 0.00172f
C8749 a_67348_20072# a_67460_18884# 0.02666f
C8750 a_25548_20408# a_26132_20452# 0.01675f
C8751 a_18268_30951# a_18628_31048# 0.0869f
C8752 _452_.CLK a_35988_18504# 0.00599f
C8753 a_67996_17272# a_67884_16839# 0.02634f
C8754 _350_.A1 a_34404_31048# 0.00234f
C8755 a_58588_11000# a_58500_9476# 0.00151f
C8756 a_61836_23544# vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I 0.00656f
C8757 a_18816_29931# a_19744_30301# 1.16391f
C8758 a_21540_1636# VPWR 0.2085f
C8759 a_63652_12612# a_64100_12612# 0.01328f
C8760 _274_.A3 a_53616_29480# 0.01837f
C8761 _474_.CLK a_52512_19715# 0.00775f
C8762 _397_.A1 _381_.A2 1.17067f
C8763 _459_.CLK a_32292_26344# 0.03226f
C8764 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I 0.75757f
C8765 a_54332_15704# a_54780_15704# 0.01222f
C8766 _390_.ZN _407_.ZN 0.04044f
C8767 a_60852_28292# VPWR 0.21094f
C8768 a_52004_11044# a_51644_11000# 0.08707f
C8769 a_63068_15271# a_63428_15368# 0.08717f
C8770 a_64212_12232# a_64100_11044# 0.02666f
C8771 a_9668_1636# a_9532_1159# 0.00168f
C8772 a_33412_18504# VPWR 0.20644f
C8773 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN a_61076_20452# 0.00636f
C8774 _397_.A2 clkbuf_1_0__f_clk.I 0.82141f
C8775 a_1380_26724# a_1468_26680# 0.28563f
C8776 a_49600_30180# VPWR 0.4074f
C8777 a_33724_1159# a_34172_1159# 0.0131f
C8778 a_64212_10664# a_64884_10664# 0.00347f
C8779 a_32476_29167# uo_out[7] 0.00412f
C8780 _371_.ZN a_27004_27815# 0.00818f
C8781 _274_.A1 _258_.I 0.00883f
C8782 a_26916_2824# a_26780_1592# 0.00154f
C8783 a_30724_2824# a_30724_1636# 0.05841f
C8784 _381_.Z a_50308_26476# 0.00171f
C8785 _303_.ZN a_39772_19975# 0.00158f
C8786 _324_.C a_56036_28292# 0.00984f
C8787 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I VPWR 1.00569f
C8788 _462_.D _335_.ZN 0.00121f
C8789 a_39796_27912# _442_.ZN 0.01084f
C8790 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_62956_23111# 0.00737f
C8791 a_59036_2727# VPWR 0.31143f
C8792 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I 0.84058f
C8793 a_36636_21543# a_37084_21543# 0.01222f
C8794 a_47076_12612# VPWR 0.20348f
C8795 _381_.Z _404_.A1 0.8538f
C8796 a_65308_18407# a_66004_18504# 0.01227f
C8797 a_1468_29383# a_1380_29480# 0.28563f
C8798 a_2724_20072# VPWR 0.20782f
C8799 a_63404_23544# a_63852_23544# 0.01255f
C8800 a_37668_15368# a_38340_15368# 0.00347f
C8801 a_1468_15704# a_1468_15271# 0.05841f
C8802 _474_.CLK _282_.ZN 0.00939f
C8803 _424_.B1 _427_.B1 0.00519f
C8804 a_36016_20893# _448_.D 0.00508f
C8805 a_59820_10567# VPWR 0.31389f
C8806 a_39772_15271# a_39684_15368# 0.28563f
C8807 a_57492_18884# VPWR 0.15752f
C8808 a_21764_23208# VPWR 0.20595f
C8809 a_35740_30951# VPWR 0.31353f
C8810 a_62172_17272# a_62196_16936# 0.00172f
C8811 _256_.A2 a_64412_29816# 0.0064f
C8812 a_41116_15271# a_41564_15271# 0.0131f
C8813 _330_.A1 _301_.A1 0.07367f
C8814 _427_.ZN vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I 0.01924f
C8815 _409_.ZN a_50704_27912# 0.00104f
C8816 a_56348_30951# _274_.A2 0.00302f
C8817 a_3708_21976# a_4156_21976# 0.0131f
C8818 a_53660_2727# a_53572_2824# 0.28563f
C8819 a_65308_17272# a_65756_17272# 0.01255f
C8820 _304_.B a_54444_26680# 0.00453f
C8821 a_49316_18504# a_50324_18504# 0.00196f
C8822 _419_.Z a_51912_20452# 0.10241f
C8823 a_19524_23208# a_19612_21543# 0.00151f
C8824 a_1380_1256# VPWR 0.20348f
C8825 a_25684_23588# a_26132_23588# 0.01328f
C8826 a_34532_1256# a_35204_1256# 0.00347f
C8827 a_22996_23588# a_22636_23544# 0.08717f
C8828 a_17844_25156# a_17484_25112# 0.08707f
C8829 a_1828_31048# VPWR 0.20348f
C8830 _383_.ZN a_48141_29480# 0.00406f
C8831 a_49740_13703# a_50100_13800# 0.08707f
C8832 a_63404_13703# a_63852_13703# 0.01288f
C8833 a_13788_2727# a_14236_2727# 0.0131f
C8834 a_4156_18840# a_4156_18407# 0.05841f
C8835 a_51240_23340# a_52920_22760# 0.00672f
C8836 _304_.B hold2.I 0.09776f
C8837 a_31284_20452# a_31372_20408# 0.28563f
C8838 a_36524_16839# a_36884_16936# 0.08707f
C8839 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN a_57468_16839# 0.00676f
C8840 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I a_58924_18840# 0.00497f
C8841 a_27676_1592# VPWR 0.29903f
C8842 _238_.I VPWR 0.88188f
C8843 a_53772_10567# a_53796_9476# 0.0016f
C8844 a_18268_30951# a_18716_30951# 0.01255f
C8845 _284_.B _281_.ZN 0.13296f
C8846 a_2812_25112# a_2812_24679# 0.05841f
C8847 _350_.A2 _334_.A1 0.00906f
C8848 _371_.A2 a_28112_27912# 0.0212f
C8849 a_932_17316# a_1380_17316# 0.01328f
C8850 a_54916_11044# a_55004_11000# 0.28563f
C8851 a_58500_11044# a_58948_11044# 0.01328f
C8852 _324_.C a_56036_27912# 0.00238f
C8853 a_44252_1592# a_44700_1592# 0.01288f
C8854 a_49652_16936# a_50324_16936# 0.00347f
C8855 a_17803_26841# a_18048_27209# 0.00232f
C8856 _402_.A1 a_49764_26724# 0.45219f
C8857 _324_.C a_50120_26476# 0.05065f
C8858 a_3260_27815# a_3708_27815# 0.0131f
C8859 _246_.B2 a_59397_26344# 0.0024f
C8860 a_18604_20408# VPWR 0.32267f
C8861 a_5052_29816# a_4964_28292# 0.0027f
C8862 a_53212_12568# VPWR 0.3185f
C8863 _290_.ZN _294_.ZN 0.09067f
C8864 _287_.A1 _362_.ZN 1.04695f
C8865 a_14596_2824# a_15044_2824# 0.01328f
C8866 a_12444_29383# a_12804_29480# 0.08717f
C8867 a_56348_30951# a_56260_31048# 0.28563f
C8868 a_56684_18407# a_56596_18504# 0.28563f
C8869 a_37444_15748# a_37308_15271# 0.00168f
C8870 a_33500_15704# a_33500_15271# 0.05841f
C8871 _342_.ZN _349_.A4 0.05271f
C8872 a_1916_7431# a_1828_7528# 0.28563f
C8873 a_54892_26680# a_54804_25156# 0.00151f
C8874 a_50748_15271# a_51108_15368# 0.08717f
C8875 a_53684_10664# VPWR 0.20614f
C8876 a_53212_27815# a_53124_27912# 0.28563f
C8877 a_2812_5863# a_2724_5960# 0.28563f
C8878 _476_.Q a_51240_19624# 0.1893f
C8879 a_19164_26247# uio_out[7] 0.0012f
C8880 _294_.A2 a_38472_30169# 0.04477f
C8881 a_2276_21640# a_2276_20452# 0.05841f
C8882 a_3708_4295# a_3620_4392# 0.28563f
C8883 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I 0.06546f
C8884 a_44744_26355# a_45232_25987# 0.8399f
C8885 a_56036_23208# a_54824_22045# 0.00187f
C8886 a_1828_15368# VPWR 0.20348f
C8887 a_57916_25112# clk 0.00706f
C8888 _416_.A1 a_40668_26247# 0.00387f
C8889 _475_.D a_46800_20937# 0.00108f
C8890 a_20084_22020# a_19724_21976# 0.08707f
C8891 vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN 0.0175f
C8892 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN 0.02642f
C8893 a_64636_2727# a_64996_2824# 0.08717f
C8894 a_38576_22504# a_38784_22504# 0.00403f
C8895 a_5388_15271# VPWR 0.35526f
C8896 a_932_14180# a_1380_14180# 0.01328f
C8897 a_48956_30951# a_49316_31048# 0.08717f
C8898 a_54444_26680# VPWR 0.32229f
C8899 _473_.Q a_47259_20127# 0.00231f
C8900 a_42982_21730# a_44038_21236# 0.00231f
C8901 a_29563_29535# VPWR 0.35863f
C8902 a_62980_17316# VPWR 0.20348f
C8903 a_1916_4295# VPWR 0.297f
C8904 a_67548_7864# VPWR 0.29679f
C8905 a_23780_1256# VPWR 0.22423f
C8906 _325_.A2 _330_.A2 0.02008f
C8907 a_60716_13703# a_60628_13800# 0.28563f
C8908 hold2.I VPWR 1.31608f
C8909 a_14236_29383# VPWR 0.29679f
C8910 a_5724_30951# VPWR 0.31143f
C8911 _311_.A2 a_33152_22091# 0.00248f
C8912 _470_.D a_44571_26841# 0.02698f
C8913 _330_.A1 a_46198_27060# 0.46741f
C8914 _480_.Q a_45088_29123# 0.00126f
C8915 a_47500_16839# a_47412_16936# 0.28563f
C8916 a_6172_1159# a_6532_1256# 0.08717f
C8917 a_41476_1636# VPWR 0.21238f
C8918 _452_.CLK a_45564_21236# 0.00172f
C8919 a_39124_16936# VPWR 0.20637f
C8920 a_50636_12135# a_51084_12135# 0.01288f
C8921 a_56236_24679# VPWR 0.33506f
C8922 a_7292_1592# a_7740_1592# 0.01288f
C8923 a_6308_29860# a_5948_29816# 0.08707f
C8924 vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN 0.00173f
C8925 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN 0.00112f
C8926 a_5052_20408# a_4964_18884# 0.00151f
C8927 a_50436_30689# VPWR 0.58776f
C8928 a_3620_2824# VPWR 0.22347f
C8929 a_51556_1636# a_51196_1592# 0.08707f
C8930 a_23196_29816# uio_out[4] 0.00152f
C8931 _243_.ZN a_58588_26247# 0.00241f
C8932 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I VPWR 0.90514f
C8933 a_56684_17272# VPWR 0.32009f
C8934 _407_.A1 a_51084_28248# 0.00991f
C8935 _475_.Q _476_.Q 0.41102f
C8936 _300_.ZN _301_.A1 0.37326f
C8937 _337_.ZN a_28552_25940# 0.00122f
C8938 _384_.ZN _470_.Q 0.00445f
C8939 _424_.A1 a_51912_20452# 0.02603f
C8940 _359_.B a_35292_26247# 0.00841f
C8941 a_3708_24679# a_4156_24679# 0.0131f
C8942 _343_.A2 uio_out[3] 0.0013f
C8943 a_44459_18559# a_44704_18191# 0.00232f
C8944 a_51308_18407# a_51220_18504# 0.28563f
C8945 _459_.CLK a_19612_26247# 0.03238f
C8946 a_56124_1159# a_56572_1159# 0.0131f
C8947 a_61612_20408# a_62060_20408# 0.012f
C8948 _346_.ZN _455_.D 0.05089f
C8949 a_64860_18840# a_65308_18840# 0.0131f
C8950 _460_.Q _288_.ZN 0.64047f
C8951 a_21428_25156# VPWR 0.20595f
C8952 _452_.D a_41536_17636# 0.22107f
C8953 a_19500_27815# a_19412_27912# 0.28563f
C8954 a_33076_20452# VPWR 0.21355f
C8955 a_31396_26724# VPWR 0.12433f
C8956 _272_.B1 VPWR 0.37011f
C8957 a_22636_30951# VPWR 0.31143f
C8958 _393_.A1 a_44948_28292# 0.00159f
C8959 a_67324_12568# VPWR 0.31547f
C8960 a_33412_15748# a_33860_15748# 0.01328f
C8961 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN a_57692_14136# 0.03478f
C8962 _381_.Z a_48384_26724# 0.00183f
C8963 _397_.A2 a_49637_28776# 0.00928f
C8964 _398_.C _282_.ZN 0.607f
C8965 _424_.A1 a_54332_20408# 0.00193f
C8966 a_27004_21543# a_27028_20452# 0.0016f
C8967 _424_.B1 _422_.ZN 0.00286f
C8968 a_2276_15748# VPWR 0.20634f
C8969 a_49092_15368# VPWR 0.21839f
C8970 a_22996_22020# a_23084_21976# 0.28563f
C8971 a_60212_25156# VPWR 0.6091f
C8972 a_26580_22020# a_27028_22020# 0.01328f
C8973 a_52540_15271# VPWR 0.32932f
C8974 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I a_50996_28292# 0.01018f
C8975 a_44812_16839# a_45260_16839# 0.01288f
C8976 _402_.A1 _437_.A1 0.98131f
C8977 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN a_53660_27815# 0.01499f
C8978 a_33948_16839# VPWR 0.32378f
C8979 _408_.ZN _411_.A2 0.43793f
C8980 a_45956_1256# VPWR 0.20968f
C8981 a_23084_30951# a_22996_31048# 0.28563f
C8982 a_56932_1256# a_57380_1256# 0.01328f
C8983 _473_.Q _419_.Z 0.09148f
C8984 _304_.B VPWR 6.47945f
C8985 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN a_66316_20408# 0.0032f
C8986 a_31920_29480# _223_.ZN 0.0152f
C8987 a_57492_13800# a_57940_13800# 0.01328f
C8988 a_36188_2727# a_36636_2727# 0.0131f
C8989 a_40644_17272# a_40556_16839# 0.02951f
C8990 a_32516_17316# VPWR 0.20348f
C8991 a_59732_10664# a_59844_9476# 0.02666f
C8992 a_55140_1636# VPWR 0.20968f
C8993 _371_.A1 a_32132_27912# 0.00264f
C8994 a_17596_1159# a_17508_1256# 0.28563f
C8995 _399_.A2 _473_.Q 0.00736f
C8996 a_47612_12135# a_47524_12232# 0.28563f
C8997 a_61500_12568# a_61524_12232# 0.00172f
C8998 _331_.ZN a_40684_19368# 0.00878f
C8999 a_14596_1636# a_14236_1592# 0.08707f
C9000 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN VPWR 0.67182f
C9001 a_54804_26724# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.00117f
C9002 a_67348_20072# a_67436_18407# 0.00151f
C9003 a_12804_29860# a_13252_29860# 0.01328f
C9004 a_9220_29860# a_9308_29816# 0.28563f
C9005 _474_.CLK a_53348_18884# 0.02283f
C9006 a_33776_29123# uo_out[4] 0.00181f
C9007 a_35292_17272# a_35740_17272# 0.01288f
C9008 a_48732_17272# a_48756_16936# 0.00172f
C9009 _287_.A2 _287_.A1 1.80873f
C9010 _424_.A2 a_44786_24120# 0.02176f
C9011 a_58052_1636# a_58500_1636# 0.01328f
C9012 a_65084_11000# a_65532_11000# 0.01288f
C9013 _459_.CLK _455_.D 0.24283f
C9014 a_26020_2824# VPWR 0.21239f
C9015 a_37386_31048# uo_out[2] 0.00182f
C9016 _459_.CLK a_17036_27815# 0.05931f
C9017 a_15244_24679# a_15604_24776# 0.08717f
C9018 a_23644_23111# a_24092_23111# 0.01288f
C9019 a_2364_23111# a_2724_23208# 0.08717f
C9020 a_53660_15704# a_54332_15704# 0.00544f
C9021 a_7428_2824# a_7516_1159# 0.0027f
C9022 a_47076_14180# VPWR 0.20952f
C9023 a_2812_18407# a_2724_18504# 0.28563f
C9024 a_61612_12135# VPWR 0.31547f
C9025 a_10788_29480# VPWR 0.20914f
C9026 a_24764_2727# a_24900_1636# 0.00154f
C9027 a_36996_2824# a_37444_2824# 0.01328f
C9028 _324_.C _404_.A1 0.07596f
C9029 a_47972_31048# VPWR 0.20452f
C9030 a_65668_23208# vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I 0.00107f
C9031 _419_.Z _475_.D 0.24907f
C9032 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN 0.06518f
C9033 a_24092_24679# VPWR 0.32732f
C9034 a_61524_23208# vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN 0.00593f
C9035 _416_.A1 _421_.B 0.18126f
C9036 a_64324_4392# VPWR 0.22383f
C9037 a_3620_7528# VPWR 0.22347f
C9038 _452_.CLK a_43008_26795# 0.00384f
C9039 _330_.A1 a_37296_22020# 0.00131f
C9040 _416_.A1 _451_.Q 0.28823f
C9041 a_55252_25156# VPWR 0.20525f
C9042 a_36636_15704# VPWR 0.3289f
C9043 a_30160_30301# uo_out[6] 0.00236f
C9044 _369_.ZN a_29575_28293# 0.06688f
C9045 a_4156_9432# a_4604_9432# 0.01222f
C9046 _230_.I _250_.C 1.1412f
C9047 a_37384_19624# a_37360_19325# 0.00918f
C9048 _330_.A1 a_39268_18840# 0.00683f
C9049 a_63428_15368# a_63292_14136# 0.00154f
C9050 a_49852_14136# a_50300_14136# 0.01288f
C9051 a_52652_18407# VPWR 0.31585f
C9052 _359_.ZN a_33188_25940# 0.39463f
C9053 _474_.D a_50660_20452# 0.05972f
C9054 _455_.Q a_23332_26344# 0.12434f
C9055 _424_.B1 a_49764_26724# 0.04213f
C9056 _411_.A2 _412_.A1 1.81472f
C9057 a_32904_28776# uo_out[7] 0.00106f
C9058 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.03721f
C9059 _325_.A2 a_43400_18909# 0.04763f
C9060 a_58500_26344# a_58364_25112# 0.00154f
C9061 _290_.ZN a_34404_31048# 0.0027f
C9062 _281_.ZN _474_.Q 0.12141f
C9063 a_44364_17272# VPWR 0.29448f
C9064 a_67124_10664# a_67012_9476# 0.02666f
C9065 a_65332_10664# a_65308_9432# 0.0016f
C9066 _358_.A3 a_34155_25273# 0.01073f
C9067 a_4940_12135# a_4964_11044# 0.0016f
C9068 a_28572_1159# a_28932_1256# 0.08717f
C9069 a_55900_12568# a_55812_11044# 0.00151f
C9070 a_58476_12135# a_58836_12232# 0.08707f
C9071 a_4852_12232# a_5300_12232# 0.01328f
C9072 a_61276_1592# VPWR 0.29679f
C9073 _346_.A2 a_22352_25987# 0.00815f
C9074 a_21092_1636# a_21540_1636# 0.01328f
C9075 a_17508_1636# a_17596_1592# 0.28563f
C9076 _452_.Q a_40468_16936# 0.00426f
C9077 a_59332_29816# VPWR 0.76405f
C9078 a_41012_23208# VPWR 0.00695f
C9079 _448_.Q a_39475_21236# 0.00422f
C9080 a_17036_21543# VPWR 0.29679f
C9081 _304_.B a_50068_27508# 0.03083f
C9082 a_48420_2824# VPWR 0.20348f
C9083 a_62396_11000# a_62508_10567# 0.02634f
C9084 _251_.A1 a_62308_27912# 0.00155f
C9085 a_22748_23111# a_22660_23208# 0.28563f
C9086 a_17396_24776# a_17844_24776# 0.01328f
C9087 a_54108_21543# VPWR 0.31907f
C9088 a_60404_28292# a_60852_28292# 0.01328f
C9089 a_51332_9476# VPWR 0.20677f
C9090 _242_.Z a_59260_26680# 0.00273f
C9091 a_54108_14136# VPWR 0.31389f
C9092 _325_.A1 a_39780_22805# 0.00107f
C9093 a_58948_2824# a_58948_1636# 0.05841f
C9094 a_24564_31048# VPWR 0.20774f
C9095 a_32964_18504# a_33412_18504# 0.01328f
C9096 _311_.Z a_37084_21543# 0.02744f
C9097 a_39548_15704# a_39996_15704# 0.01288f
C9098 a_55476_12232# VPWR 0.20622f
C9099 a_43492_15748# a_43580_15704# 0.28563f
C9100 _304_.B _424_.B2 0.00439f
C9101 _435_.A3 _434_.ZN 0.45181f
C9102 a_34716_20937# a_35060_20569# 0.00275f
C9103 a_49112_29885# a_49600_30180# 0.8399f
C9104 a_38676_20452# a_38764_20408# 0.28563f
C9105 a_28903_24776# VPWR 0.50869f
C9106 a_28124_30600# _340_.A2 0.00932f
C9107 a_61188_20072# VPWR 0.15132f
C9108 a_53100_16839# a_53124_15748# 0.0016f
C9109 a_32740_21640# a_32716_20408# 0.0016f
C9110 _305_.A2 _304_.ZN 0.00366f
C9111 a_8636_2727# a_8996_2824# 0.08717f
C9112 _395_.A2 a_50792_26344# 0.02578f
C9113 a_50436_15748# VPWR 0.24967f
C9114 _325_.A2 _448_.D 0.1406f
C9115 a_49540_9476# a_49628_9432# 0.28563f
C9116 _442_.ZN a_40580_26344# 0.00671f
C9117 _461_.D a_32476_29167# 0.22071f
C9118 a_57604_14180# a_57244_14136# 0.08663f
C9119 _459_.CLK _454_.D 0.08209f
C9120 _452_.CLK a_38752_26344# 0.00128f
C9121 a_62508_21976# vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I 0.00473f
C9122 _300_.A2 _319_.A3 0.00107f
C9123 _412_.A1 _399_.ZN 0.04094f
C9124 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN 0.14067f
C9125 a_58588_2727# a_59036_2727# 0.0131f
C9126 a_46628_12612# a_47076_12612# 0.01328f
C9127 a_57940_20452# VPWR 0.15775f
C9128 a_36100_26344# VPWR 0.20348f
C9129 a_2276_20072# a_2724_20072# 0.01328f
C9130 a_1828_12232# a_1828_11044# 0.05841f
C9131 a_11324_1159# VPWR 0.34493f
C9132 a_39996_1159# a_39908_1256# 0.28563f
C9133 a_932_3204# a_1020_3160# 0.28563f
C9134 _383_.ZN VPWR 0.42824f
C9135 a_5300_21640# VPWR 0.21406f
C9136 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I a_67996_21976# 0.01016f
C9137 a_47388_17272# a_47836_17272# 0.01288f
C9138 a_51332_17316# a_51420_17272# 0.28563f
C9139 _473_.Q _416_.A2 0.60331f
C9140 a_50068_27508# VPWR 0.89223f
C9141 _350_.A2 _370_.ZN 0.64202f
C9142 a_44700_1592# a_44700_1159# 0.05841f
C9143 a_67324_1592# a_67772_1592# 0.01222f
C9144 a_59372_10567# a_59820_10567# 0.01288f
C9145 a_45372_10567# a_45732_10664# 0.08717f
C9146 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I 0.00129f
C9147 a_5636_2824# a_5500_1592# 0.00154f
C9148 a_35292_30951# a_35740_30951# 0.01222f
C9149 _459_.CLK a_28036_26724# 0.00637f
C9150 a_21316_23208# a_21764_23208# 0.01328f
C9151 a_33276_23111# a_33636_23208# 0.08663f
C9152 a_63852_23111# VPWR 0.29679f
C9153 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN a_54824_22045# 0.00173f
C9154 a_5300_26344# a_5388_24679# 0.0027f
C9155 a_2812_23544# VPWR 0.30213f
C9156 a_33152_22091# a_34032_22505# 0.00306f
C9157 a_62308_9476# VPWR 0.20595f
C9158 a_4604_3160# VPWR 0.32824f
C9159 a_15692_21543# a_15604_21640# 0.28563f
C9160 a_2812_6296# VPWR 0.30213f
C9161 a_1916_13703# VPWR 0.297f
C9162 a_3620_29480# a_3620_28292# 0.05841f
C9163 a_27900_21543# a_28348_21543# 0.01288f
C9164 _325_.A1 a_39796_22504# 0.42892f
C9165 a_58911_30644# a_59163_30644# 0.00184f
C9166 a_54804_26724# a_54892_26680# 0.28563f
C9167 a_43003_28409# _330_.A1 0.00192f
C9168 _452_.CLK a_33948_18840# 0.00252f
C9169 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN _248_.B1 0.33812f
C9170 _424_.A2 a_47776_20893# 0.00107f
C9171 a_36996_25156# VPWR 0.20348f
C9172 a_46852_15748# a_46492_15704# 0.08707f
C9173 a_5052_11000# VPWR 0.33516f
C9174 _395_.A2 _281_.ZN 0.10306f
C9175 _435_.ZN a_39536_23588# 0.0063f
C9176 _424_.B2 VPWR 0.55211f
C9177 a_59396_2824# a_59844_2824# 0.01328f
C9178 a_9635_30644# a_9668_29860# 0.02559f
C9179 a_66540_19975# a_66452_20072# 0.28563f
C9180 _474_.CLK a_54444_18407# 0.00239f
C9181 _237_.A1 a_60285_30600# 0.03951f
C9182 _324_.C a_48384_26724# 0.00104f
C9183 _459_.CLK a_41228_27815# 0.00112f
C9184 a_31708_18840# VPWR 0.29679f
C9185 _359_.B a_37844_29860# 0.00114f
C9186 a_14796_26247# VPWR 0.30073f
C9187 _226_.ZN a_42154_21236# 0.00108f
C9188 a_20060_2727# a_19972_2824# 0.28563f
C9189 _281_.ZN a_46984_23588# 0.16593f
C9190 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.6831f
C9191 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN 0.00552f
C9192 a_37968_31048# uo_out[1] 0.00163f
C9193 _304_.B a_44744_26355# 0.04242f
C9194 _424_.A2 _395_.A3 0.02532f
C9195 a_54780_9432# a_55228_9432# 0.0131f
C9196 a_1380_31048# a_1828_31048# 0.01328f
C9197 a_65444_14180# a_65892_14180# 0.01328f
C9198 _459_.Q a_32292_26344# 0.02411f
C9199 _475_.D _416_.A2 0.01024f
C9200 a_62308_14180# a_61948_14136# 0.08707f
C9201 _474_.Q a_50660_20452# 0.01888f
C9202 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN 0.30261f
C9203 a_52452_24072# _384_.A1 0.00505f
C9204 _424_.ZN a_52944_19759# 0.00134f
C9205 _397_.A1 a_48596_28292# 0.01821f
C9206 _337_.A3 a_25124_28776# 0.25548f
C9207 _290_.ZN _362_.B 0.654f
C9208 a_62420_13800# a_62396_12568# 0.0016f
C9209 a_29716_31048# uio_out[0] 0.00101f
C9210 a_33724_1159# VPWR 0.30128f
C9211 _474_.CLK vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I 0.04707f
C9212 a_50972_1159# a_51332_1256# 0.08717f
C9213 a_50100_12232# a_50212_11044# 0.02666f
C9214 a_66228_12232# a_66676_12232# 0.01328f
C9215 a_27228_1592# a_27676_1592# 0.01288f
C9216 a_31172_1636# a_31260_1592# 0.28563f
C9217 a_45060_31048# a_45012_29816# 0.00125f
C9218 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN 0.63963f
C9219 a_36636_21543# VPWR 0.31201f
C9220 a_63404_23544# VPWR 0.2963f
C9221 _267_.A1 a_55140_28292# 0.01095f
C9222 a_58500_26344# clk 0.002f
C9223 a_32592_25227# a_34396_24679# 0.00456f
C9224 a_33148_25641# a_33164_24679# 0.0019f
C9225 a_56460_10567# a_56372_10664# 0.28563f
C9226 _264_.B hold1.Z 0.00221f
C9227 hold2.I _260_.ZN 0.88921f
C9228 a_3708_21976# VPWR 0.33374f
C9229 _402_.A1 a_43492_27912# 0.00625f
C9230 _279_.Z a_48321_23208# 0.03193f
C9231 a_25684_23588# VPWR 0.20947f
C9232 a_39796_22504# _327_.A2 0.00243f
C9233 a_51240_23340# VPWR 0.53621f
C9234 a_26556_21543# a_26916_21640# 0.08707f
C9235 a_63404_13703# VPWR 0.31556f
C9236 a_2276_18884# a_1916_18840# 0.08717f
C9237 a_13788_2727# VPWR 0.31143f
C9238 _467_.D a_16500_28292# 0.03726f
C9239 a_4068_18884# a_4516_18884# 0.01328f
C9240 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN 0.6364f
C9241 _355_.C a_22996_28292# 0.0302f
C9242 _459_.CLK a_32848_29123# 0.01308f
C9243 a_58500_11044# VPWR 0.21691f
C9244 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I a_58836_17316# 0.00409f
C9245 a_53212_15704# a_53660_15704# 0.012f
C9246 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I a_63964_19975# 0.00305f
C9247 _371_.A3 a_28036_26724# 0.00521f
C9248 a_64772_15748# a_64860_15704# 0.28563f
C9249 _330_.A1 a_35492_20072# 0.01625f
C9250 a_3260_27815# VPWR 0.30487f
C9251 a_36548_26344# a_36548_25156# 0.05841f
C9252 a_58476_20408# vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN 0.001f
C9253 _438_.A2 a_37532_25112# 0.00269f
C9254 _373_.ZN _371_.A2 0.02733f
C9255 a_30812_2727# a_31396_2824# 0.01675f
C9256 a_64860_3160# a_64996_2824# 0.00168f
C9257 a_65084_30951# vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.00525f
C9258 _421_.A1 a_47297_25596# 0.06473f
C9259 a_44744_26355# VPWR 1.10271f
C9260 a_48888_19243# a_48172_18840# 0.00367f
C9261 a_4964_23588# a_5052_23544# 0.28563f
C9262 a_60516_9476# a_60604_9432# 0.28563f
C9263 a_4068_7908# a_4156_7864# 0.28563f
C9264 a_4964_6340# a_5052_6296# 0.28563f
C9265 _325_.A2 a_39684_20072# 0.00869f
C9266 _316_.ZN a_34160_20523# 0.00369f
C9267 a_20308_20452# a_19948_20408# 0.08717f
C9268 a_3260_30951# a_3620_31048# 0.08717f
C9269 a_57244_27815# _241_.Z 0.00532f
C9270 a_58911_30644# ui_in[3] 0.01221f
C9271 a_25436_1592# a_25572_1256# 0.00168f
C9272 a_7292_1592# VPWR 0.3289f
C9273 a_56708_12612# a_56796_12568# 0.28563f
C9274 _459_.CLK a_17932_25112# 0.00189f
C9275 _393_.A1 a_46198_27060# 0.00147f
C9276 _324_.C _435_.A3 0.47014f
C9277 _302_.Z a_42982_21730# 0.01705f
C9278 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_62508_23111# 0.00207f
C9279 a_24004_24776# a_23980_23544# 0.0016f
C9280 a_62396_1159# a_62308_1256# 0.28563f
C9281 a_61612_20408# VPWR 0.31431f
C9282 a_56124_1159# VPWR 0.3289f
C9283 a_45696_20072# a_47552_19715# 0.02307f
C9284 _416_.A2 a_47252_18884# 0.00415f
C9285 a_57044_12232# a_57156_11044# 0.02666f
C9286 a_53236_12232# a_53212_11000# 0.0016f
C9287 a_34532_1636# a_34172_1592# 0.08707f
C9288 a_34155_25273# a_34400_25641# 0.00232f
C9289 a_64860_18840# VPWR 0.30145f
C9290 _416_.A1 a_42161_24776# 0.00963f
C9291 _441_.ZN a_39536_23588# 0.00526f
C9292 a_44476_27815# _330_.A1 0.03789f
C9293 _452_.CLK a_36300_23544# 0.00135f
C9294 a_53236_10664# a_53684_10664# 0.01328f
C9295 a_67212_10567# a_67572_10664# 0.08717f
C9296 _467_.D a_17396_27912# 0.00242f
C9297 a_22300_1159# a_22748_1159# 0.0131f
C9298 _229_.I a_63313_28776# 0.00452f
C9299 _304_.B _260_.ZN 0.74699f
C9300 _370_.B VPWR 0.56352f
C9301 _355_.C a_24304_29480# 0.01262f
C9302 a_31484_26680# a_30724_26020# 0.02977f
C9303 a_26580_22020# VPWR 0.2131f
C9304 vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I 0.15767f
C9305 _393_.ZN _384_.ZN 0.00515f
C9306 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I 0.00267f
C9307 a_33860_18884# a_33500_18840# 0.08717f
C9308 _384_.A3 a_51332_24372# 0.05296f
C9309 a_24900_21640# a_25348_21640# 0.01328f
C9310 a_36188_2727# VPWR 0.31143f
C9311 a_52228_2824# a_52316_1159# 0.0027f
C9312 a_57492_13800# VPWR 0.21191f
C9313 _459_.D a_30476_23544# 0.00193f
C9314 a_1380_15368# a_1828_15368# 0.01328f
C9315 a_12804_29860# VPWR 0.20614f
C9316 a_55252_26724# VPWR 0.2078f
C9317 _350_.A2 a_31068_28292# 0.02879f
C9318 a_65084_11000# VPWR 0.32163f
C9319 a_3260_15271# a_3172_15368# 0.28563f
C9320 a_21964_21976# a_21852_21543# 0.02634f
C9321 a_23644_23111# VPWR 0.31547f
C9322 a_4940_15271# a_5388_15271# 0.01222f
C9323 _247_.ZN a_59380_27508# 0.00886f
C9324 _336_.A1 _358_.A2 0.0052f
C9325 a_66652_17272# a_66564_15748# 0.00151f
C9326 a_53996_26680# a_54444_26680# 0.01255f
C9327 a_42236_2727# a_42148_2824# 0.28563f
C9328 _294_.A2 a_34084_28776# 0.02004f
C9329 a_63764_23208# a_64212_23208# 0.01328f
C9330 _285_.Z a_39748_29480# 0.00348f
C9331 a_62532_17316# a_62980_17316# 0.01328f
C9332 _260_.A1 a_41642_25156# 0.00145f
C9333 _249_.A2 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN 0.43867f
C9334 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I _248_.B1 0.16858f
C9335 _397_.A2 _412_.A1 0.0385f
C9336 a_64076_16839# a_64436_16936# 0.08717f
C9337 _281_.ZN _427_.A2 0.07018f
C9338 a_65756_9432# a_66204_9432# 0.0131f
C9339 a_67100_7864# a_67548_7864# 0.0131f
C9340 a_18740_23588# a_18828_23544# 0.28563f
C9341 a_23108_1256# a_23780_1256# 0.00347f
C9342 a_3620_25156# a_3708_25112# 0.28563f
C9343 a_14796_23544# a_15244_23544# 0.01288f
C9344 a_1468_4295# a_1916_4295# 0.0131f
C9345 a_64860_4728# a_64860_4295# 0.05841f
C9346 _281_.ZN a_51196_21543# 0.09788f
C9347 _416_.A1 a_50996_28292# 0.00578f
C9348 a_66428_14136# a_66316_13703# 0.02634f
C9349 a_2364_2727# a_2812_2727# 0.0131f
C9350 a_52428_13703# a_52876_13703# 0.01288f
C9351 a_34644_16936# a_34620_15271# 0.00134f
C9352 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I a_60940_15704# 0.00708f
C9353 a_18268_30951# a_18180_31048# 0.28563f
C9354 a_13788_29383# a_14236_29383# 0.0131f
C9355 _350_.A1 a_33956_31048# 0.00164f
C9356 _452_.CLK a_35540_18504# 0.00594f
C9357 a_21092_1636# VPWR 0.2085f
C9358 a_50300_12568# a_50188_12135# 0.02634f
C9359 a_68020_20452# a_67884_19975# 0.00168f
C9360 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I 0.62955f
C9361 a_5276_30951# a_5724_30951# 0.01255f
C9362 _274_.A3 a_53412_29480# 0.00127f
C9363 _474_.CLK a_52024_20083# 0.02647f
C9364 _324_.C _399_.A2 0.00286f
C9365 _459_.CLK a_31844_26344# 0.02067f
C9366 a_60404_28292# VPWR 0.20334f
C9367 a_63068_15271# a_62980_15368# 0.28563f
C9368 a_41028_1636# a_41476_1636# 0.01328f
C9369 a_32964_18504# VPWR 0.20348f
C9370 a_51556_11044# a_51644_11000# 0.28563f
C9371 a_47612_11000# a_48060_11000# 0.01288f
C9372 a_38676_16936# a_39124_16936# 0.01328f
C9373 a_55788_24679# a_56236_24679# 0.012f
C9374 _336_.A1 _355_.ZN 0.05797f
C9375 _284_.B a_47636_25940# 1.5187f
C9376 a_64860_15704# a_64996_15368# 0.00168f
C9377 a_1380_26724# a_1020_26680# 0.08717f
C9378 a_3172_26724# a_3620_26724# 0.01328f
C9379 a_32848_29123# uo_out[7] 0.00588f
C9380 a_49112_29885# VPWR 1.14825f
C9381 _260_.ZN VPWR 0.98764f
C9382 _324_.C a_55588_28292# 0.0019f
C9383 _379_.A2 a_22100_29480# 0.00218f
C9384 a_61689_29860# VPWR 0.00601f
C9385 _355_.C _371_.A2 0.06923f
C9386 a_49852_30951# a_50436_30689# 0.01958f
C9387 a_35728_29480# a_36116_29167# 0.00393f
C9388 a_39796_27912# a_39536_26795# 0.00187f
C9389 a_37291_29535# a_37576_29535# 0.00277f
C9390 a_46628_12612# VPWR 0.20348f
C9391 a_58588_2727# VPWR 0.31968f
C9392 _393_.A1 a_46580_28292# 0.01426f
C9393 a_65308_18407# a_65220_18504# 0.28563f
C9394 a_15156_26344# a_15604_26344# 0.01328f
C9395 a_3172_2824# a_3620_2824# 0.01328f
C9396 a_1020_29383# a_1380_29480# 0.08717f
C9397 a_2276_20072# VPWR 0.20634f
C9398 a_58500_26344# a_58948_26344# 0.01328f
C9399 _346_.B a_21540_28292# 0.00758f
C9400 a_59372_10567# VPWR 0.31389f
C9401 a_37744_20452# _323_.A3 0.00186f
C9402 a_39324_15271# a_39684_15368# 0.08717f
C9403 a_28908_21976# a_28796_21543# 0.02634f
C9404 a_35292_30951# VPWR 0.32508f
C9405 a_21316_23208# VPWR 0.20595f
C9406 _304_.A1 _302_.Z 0.05832f
C9407 _255_.I ui_in[2] 0.00185f
C9408 _427_.ZN a_55452_21543# 0.01131f
C9409 _330_.A1 a_37408_23208# 0.003f
C9410 _399_.ZN _473_.Q 0.00262f
C9411 _409_.ZN a_50276_27912# 0.01541f
C9412 a_2812_28248# a_3260_28248# 0.0131f
C9413 _250_.A2 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN 0.1051f
C9414 a_53212_2727# a_53572_2824# 0.08717f
C9415 _304_.B a_53996_26680# 0.00469f
C9416 a_19276_23544# a_19188_22020# 0.00151f
C9417 _360_.ZN VPWR 0.36736f
C9418 _419_.Z a_51428_20452# 0.00627f
C9419 a_30724_16936# a_30724_15748# 0.05841f
C9420 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I 0.00144f
C9421 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I 0.64143f
C9422 a_20980_25156# a_21428_25156# 0.01328f
C9423 a_22548_23588# a_22636_23544# 0.28563f
C9424 a_17396_25156# a_17484_25112# 0.28563f
C9425 a_1380_31048# VPWR 0.20348f
C9426 a_63292_14136# a_63316_13800# 0.00172f
C9427 _397_.Z _475_.Q 0.0029f
C9428 a_49740_13703# a_49652_13800# 0.28563f
C9429 a_31284_20452# a_30924_20408# 0.08717f
C9430 a_32628_20452# a_33076_20452# 0.01328f
C9431 a_22188_30951# a_22636_30951# 0.01255f
C9432 a_36060_19369# a_36404_19001# 0.00275f
C9433 a_58063_30644# _270_.A2 0.0434f
C9434 a_57120_31048# _272_.B1 0.02409f
C9435 a_36524_16839# a_36436_16936# 0.28563f
C9436 a_57156_27912# VPWR 0.20495f
C9437 a_63740_11000# a_63652_9476# 0.00151f
C9438 _384_.ZN a_50084_24328# 0.00192f
C9439 a_27228_1592# VPWR 0.36633f
C9440 _284_.B a_46156_25112# 0.0134f
C9441 a_66876_12568# a_67324_12568# 0.01288f
C9442 a_57244_12568# a_57132_12135# 0.02634f
C9443 _460_.Q a_33520_25597# 0.01058f
C9444 a_4068_1636# a_4516_1636# 0.01328f
C9445 a_4964_25156# a_4940_24679# 0.00172f
C9446 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN a_60416_25156# 0.00237f
C9447 _371_.A2 a_27908_27912# 0.00613f
C9448 a_57492_12232# a_57580_10567# 0.00151f
C9449 a_1468_11000# a_1468_10567# 0.05841f
C9450 a_54916_11044# a_54556_11000# 0.08707f
C9451 _397_.A1 _400_.ZN 0.05752f
C9452 _350_.A1 _359_.B 0.20838f
C9453 a_44700_1159# a_45148_1159# 0.0131f
C9454 a_3620_27912# a_3620_26724# 0.05841f
C9455 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN a_65556_23588# 0.0273f
C9456 a_44300_19001# VPWR 0.00246f
C9457 a_62532_18884# a_62980_18884# 0.01328f
C9458 a_21652_20452# VPWR 0.21296f
C9459 a_60292_12612# VPWR 0.21323f
C9460 a_1828_15748# a_2276_15748# 0.01328f
C9461 _245_.Z a_59828_26724# 0.0036f
C9462 _355_.C a_22996_25156# 0.00618f
C9463 a_10428_2727# a_10564_1636# 0.00154f
C9464 a_48644_15368# a_49092_15368# 0.01328f
C9465 a_12444_29383# a_12356_29480# 0.28563f
C9466 _251_.A1 _268_.A1 0.01229f
C9467 a_24864_29931# _349_.A4 0.02667f
C9468 a_16588_28248# a_16588_27815# 0.05841f
C9469 a_53236_10664# VPWR 0.20614f
C9470 a_50748_15271# a_50660_15368# 0.28563f
C9471 _424_.A2 _427_.B1 0.00369f
C9472 a_1468_7431# a_1828_7528# 0.08717f
C9473 a_52764_27815# a_53124_27912# 0.0869f
C9474 a_3260_4295# a_3620_4392# 0.08717f
C9475 a_2364_5863# a_2724_5960# 0.08717f
C9476 _294_.A2 a_31080_29977# 0.00118f
C9477 a_44340_26183# a_45128_26031# 0.02112f
C9478 _381_.Z _411_.A2 0.06486f
C9479 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I a_66540_19975# 0.00105f
C9480 a_52092_15271# a_52540_15271# 0.0131f
C9481 a_1380_15368# VPWR 0.20348f
C9482 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I 0.00229f
C9483 _416_.A1 a_40220_26247# 0.00525f
C9484 a_64636_2727# a_64548_2824# 0.28563f
C9485 a_15692_21976# a_16140_21976# 0.01288f
C9486 a_19636_22020# a_19724_21976# 0.28563f
C9487 a_55788_25112# clk 0.00706f
C9488 a_4940_15271# VPWR 0.31945f
C9489 a_23084_23544# a_22996_22020# 0.00151f
C9490 a_4604_17272# a_4516_15748# 0.0027f
C9491 _330_.A1 _412_.A1 1.22281f
C9492 a_42982_21730# a_43814_21236# 0.10659f
C9493 a_33500_16839# a_33948_16839# 0.0131f
C9494 a_53996_26680# VPWR 0.33401f
C9495 a_48956_30951# a_48868_31048# 0.28563f
C9496 a_62532_17316# VPWR 0.20348f
C9497 a_30052_23208# a_30140_21543# 0.0027f
C9498 a_28556_29167# VPWR 0.39696f
C9499 a_67100_7864# VPWR 0.29679f
C9500 a_23108_1256# VPWR 0.20968f
C9501 a_29716_23588# a_30388_23588# 0.00347f
C9502 _325_.A2 a_38644_19368# 0.01553f
C9503 a_45508_1256# a_45956_1256# 0.01328f
C9504 a_41056_30669# _304_.B 0.4008f
C9505 a_1468_4295# VPWR 0.29679f
C9506 a_57244_14136# a_57156_12612# 0.00151f
C9507 a_46180_13800# a_46628_13800# 0.01328f
C9508 a_13788_29383# VPWR 0.29679f
C9509 a_24764_2727# a_25212_2727# 0.0131f
C9510 a_60268_13703# a_60628_13800# 0.08707f
C9511 a_5276_30951# VPWR 0.31143f
C9512 a_43232_29480# a_45088_29123# 0.02307f
C9513 a_47052_16839# a_47412_16936# 0.08707f
C9514 _480_.Q a_44795_29535# 0.00145f
C9515 _470_.D a_44864_27165# 0.05052f
C9516 a_52340_10664# a_52228_9476# 0.02666f
C9517 a_50548_10664# a_50524_9432# 0.0016f
C9518 a_38676_16936# VPWR 0.20637f
C9519 a_41028_1636# VPWR 0.21092f
C9520 a_6172_1159# a_6084_1256# 0.28563f
C9521 a_64188_12568# a_64300_12135# 0.02634f
C9522 a_54108_12568# a_54132_12232# 0.00172f
C9523 a_55788_24679# VPWR 0.29679f
C9524 _260_.A2 a_41642_25156# 0.0312f
C9525 _252_.B a_59828_26724# 0.00497f
C9526 a_18828_25112# a_18716_24679# 0.02634f
C9527 _230_.I _258_.I 0.00448f
C9528 a_1916_29816# a_2364_29816# 0.01288f
C9529 a_5860_29860# a_5948_29816# 0.28563f
C9530 _416_.A1 _402_.B 0.00605f
C9531 a_32068_17316# a_32516_17316# 0.01328f
C9532 a_4604_15704# a_4516_14180# 0.0027f
C9533 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN a_67772_21543# 0.00168f
C9534 _311_.Z VPWR 0.85753f
C9535 a_49852_30951# VPWR 0.34212f
C9536 a_61412_11044# a_61860_11044# 0.01328f
C9537 a_41048_17341# a_42484_16936# 0.00116f
C9538 a_52004_11044# a_51980_10567# 0.00172f
C9539 a_48060_11000# a_48060_10567# 0.05841f
C9540 a_61724_15271# a_61860_14180# 0.00154f
C9541 vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I 0.70581f
C9542 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN 0.00197f
C9543 a_61412_17316# VPWR 0.15832f
C9544 a_51108_1636# a_51196_1592# 0.28563f
C9545 a_54692_1636# a_55140_1636# 0.01328f
C9546 a_3172_2824# VPWR 0.20993f
C9547 _384_.A3 a_51668_23340# 0.00476f
C9548 a_31620_20072# a_31620_18884# 0.05841f
C9549 a_3260_23111# a_3708_23111# 0.0131f
C9550 _452_.CLK _358_.A3 0.52665f
C9551 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN 0.03922f
C9552 a_62844_27815# vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN 0.00558f
C9553 _459_.CLK a_19164_26247# 0.00915f
C9554 a_50860_18407# a_51220_18504# 0.08717f
C9555 _346_.ZN a_20844_26680# 0.03601f
C9556 a_44612_2824# a_44612_1636# 0.05841f
C9557 a_40804_2824# a_40668_1592# 0.00154f
C9558 a_52564_18504# a_52652_16839# 0.00151f
C9559 a_49316_18504# VPWR 0.21855f
C9560 a_20980_25156# VPWR 0.20792f
C9561 _452_.D a_41048_17341# 0.28621f
C9562 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I 0.00152f
C9563 a_3620_27912# a_4068_27912# 0.01328f
C9564 _296_.ZN uo_out[0] 1.90653f
C9565 a_22188_30951# VPWR 0.31143f
C9566 a_32628_20452# VPWR 0.20665f
C9567 a_57120_31048# VPWR 0.01432f
C9568 a_66876_12568# VPWR 0.31547f
C9569 _475_.D a_46252_19759# 0.00278f
C9570 a_38652_15704# a_38788_15368# 0.00168f
C9571 _248_.B1 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN 0.00323f
C9572 a_25572_2824# a_26020_2824# 0.01328f
C9573 _416_.A2 _416_.ZN 0.12128f
C9574 a_25796_27912# a_26468_27912# 0.00347f
C9575 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN _250_.B 0.00835f
C9576 _437_.A1 _304_.A1 0.07804f
C9577 _284_.ZN a_43564_27209# 0.05288f
C9578 _272_.B1 a_58116_30344# 0.00197f
C9579 _424_.A1 a_53884_20408# 0.00498f
C9580 _424_.B1 a_51108_21640# 0.01222f
C9581 a_1828_15748# VPWR 0.20348f
C9582 a_48644_15368# VPWR 0.21038f
C9583 _402_.A1 a_43736_25896# 0.24221f
C9584 _281_.A1 _419_.Z 0.00185f
C9585 _279_.Z a_47689_25156# 0.00303f
C9586 _352_.A2 a_28891_25273# 0.0039f
C9587 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN 0.09574f
C9588 a_22996_22020# a_22636_21976# 0.08707f
C9589 _268_.A2 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.02994f
C9590 a_52092_15271# VPWR 0.32932f
C9591 a_46628_14180# a_47076_14180# 0.01328f
C9592 a_34396_17272# a_34308_15748# 0.0027f
C9593 _304_.B a_41099_26841# 0.0458f
C9594 a_33500_16839# VPWR 0.30042f
C9595 a_22636_30951# a_22996_31048# 0.08663f
C9596 a_45508_1256# VPWR 0.20348f
C9597 a_41056_30669# VPWR 0.48044f
C9598 a_61052_14136# a_60964_12612# 0.00151f
C9599 a_3620_13800# a_3620_12612# 0.05841f
C9600 _274_.A1 _267_.A1 0.06632f
C9601 _246_.B2 a_59572_29076# 0.02278f
C9602 a_22064_27912# a_23420_26247# 0.00113f
C9603 _454_.D a_22352_25987# 0.00101f
C9604 a_16948_23208# a_16948_22020# 0.05841f
C9605 a_32068_17316# VPWR 0.20348f
C9606 a_54692_1636# VPWR 0.20348f
C9607 a_17148_1159# a_17508_1256# 0.08717f
C9608 _395_.A3 a_49988_21236# 0.00132f
C9609 a_52540_12568# a_52452_11044# 0.00151f
C9610 a_62844_27815# VPWR 0.32561f
C9611 a_61164_12135# a_61612_12135# 0.01288f
C9612 a_10204_1592# a_10652_1592# 0.01288f
C9613 a_14148_1636# a_14236_1592# 0.28563f
C9614 a_10340_29480# a_10788_29480# 0.01328f
C9615 a_47164_12135# a_47524_12232# 0.08717f
C9616 a_30924_23544# a_31036_23111# 0.02634f
C9617 a_33483_29535# uo_out[4] 0.00133f
C9618 a_58164_16936# vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I 0.00155f
C9619 a_9220_29860# a_8860_29816# 0.08707f
C9620 _336_.Z a_30240_24776# 0.00274f
C9621 a_47524_31048# a_47972_31048# 0.01328f
C9622 a_54916_15368# a_54916_14180# 0.05841f
C9623 a_58948_11044# a_58924_10567# 0.00172f
C9624 a_55004_11000# a_55116_10567# 0.02634f
C9625 _459_.CLK a_20844_26680# 0.00836f
C9626 a_25572_2824# VPWR 0.21094f
C9627 a_30364_1592# a_30364_1159# 0.05841f
C9628 _459_.CLK a_16588_27815# 0.0079f
C9629 a_2364_23111# a_2276_23208# 0.28563f
C9630 a_23644_24679# a_24092_24679# 0.01288f
C9631 a_15244_24679# a_15156_24776# 0.28563f
C9632 a_2276_9096# a_2724_9096# 0.01328f
C9633 _248_.B1 VPWR 1.11993f
C9634 a_67100_1159# a_67548_1159# 0.01222f
C9635 _455_.Q a_20396_27815# 0.00111f
C9636 a_31708_19975# a_32156_19975# 0.0131f
C9637 a_3172_7528# a_3620_7528# 0.01328f
C9638 _304_.B _407_.ZN 0.07332f
C9639 a_4068_5960# a_4852_5960# 0.00276f
C9640 a_46628_14180# VPWR 0.20952f
C9641 a_2364_18407# a_2724_18504# 0.08717f
C9642 a_33052_18407# a_33500_18407# 0.0131f
C9643 _287_.A2 a_30724_26020# 0.00118f
C9644 a_54804_25156# a_55252_25156# 0.01328f
C9645 _330_.A2 a_39264_18147# 0.01618f
C9646 a_61164_12135# VPWR 0.31547f
C9647 a_10340_29480# VPWR 0.20722f
C9648 a_36188_15704# a_36636_15704# 0.01288f
C9649 a_26160_27165# _352_.ZN 0.00854f
C9650 _383_.A2 _411_.A2 0.00114f
C9651 _242_.Z _243_.ZN 0.13817f
C9652 a_47524_31048# VPWR 0.20875f
C9653 _419_.Z a_47271_21640# 0.04102f
C9654 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN VPWR 1.39693f
C9655 a_23644_24679# VPWR 0.32277f
C9656 a_51332_15748# a_51196_15271# 0.00168f
C9657 a_47388_15704# a_47388_15271# 0.05841f
C9658 a_3172_7528# VPWR 0.20993f
C9659 a_5300_4392# VPWR 0.21488f
C9660 a_54804_25156# VPWR 0.20622f
C9661 a_36188_15704# VPWR 0.3289f
C9662 _424_.A2 _422_.ZN 0.04742f
C9663 _246_.B2 _257_.B 0.06286f
C9664 a_52204_18407# a_52652_18407# 0.0131f
C9665 _402_.A1 _417_.A2 0.00447f
C9666 a_29356_21976# a_29804_21976# 0.012f
C9667 _430_.ZN _434_.ZN 0.11514f
C9668 _230_.I a_62148_29505# 0.01998f
C9669 VPWR uio_oe[2] 0.08163f
C9670 a_41099_26841# VPWR 0.36602f
C9671 a_66788_15368# a_66788_14180# 0.05841f
C9672 _474_.D a_50212_20452# 0.01235f
C9673 _245_.I1 a_64212_23588# 0.0021f
C9674 a_52204_18407# VPWR 0.31838f
C9675 a_23084_28248# _454_.Q 0.03132f
C9676 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN VPWR 0.75187f
C9677 a_67908_1256# VPWR 0.20924f
C9678 _279_.Z _399_.A1 0.02203f
C9679 _284_.A2 _448_.Q 0.01877f
C9680 _226_.ZN a_40668_20408# 0.00726f
C9681 _452_.CLK _324_.B 0.20943f
C9682 a_51892_13800# a_52004_12612# 0.02666f
C9683 a_47164_2727# a_47612_2727# 0.0131f
C9684 a_58500_21640# vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.00229f
C9685 _223_.ZN uo_out[6] 0.05834f
C9686 a_48060_18407# a_48196_17316# 0.00154f
C9687 a_24004_23208# a_23892_22020# 0.02666f
C9688 a_28572_1159# a_28484_1256# 0.28563f
C9689 _358_.A3 a_34448_25597# 0.02373f
C9690 a_60828_1592# VPWR 0.29679f
C9691 a_58476_12135# a_58388_12232# 0.28563f
C9692 a_17508_1636# a_17148_1592# 0.08707f
C9693 _346_.A2 a_22059_26399# 0.00872f
C9694 a_15580_29816# a_16028_29816# 0.012f
C9695 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I clk 0.0658f
C9696 _452_.Q a_40020_16936# 0.00112f
C9697 a_58116_30344# VPWR 0.81902f
C9698 a_16588_21543# VPWR 0.29679f
C9699 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I _241_.Z 0.00727f
C9700 _281_.A1 _424_.A1 0.05435f
C9701 a_65892_11044# a_65868_10567# 0.00172f
C9702 a_48060_10567# a_48508_10567# 0.0131f
C9703 _251_.A1 a_59036_26247# 0.0028f
C9704 a_60828_1592# a_61276_1592# 0.01288f
C9705 a_47972_2824# VPWR 0.20348f
C9706 a_932_23208# a_1380_23208# 0.01328f
C9707 a_22300_23111# a_22660_23208# 0.08707f
C9708 hold1.Z a_44038_21236# 0.2378f
C9709 a_53660_21543# VPWR 0.33173f
C9710 a_22996_31048# VPWR 0.21171f
C9711 a_50884_9476# VPWR 0.2131f
C9712 _407_.ZN VPWR 0.48451f
C9713 a_16588_21543# a_17036_21543# 0.0131f
C9714 _419_.A4 clk 0.00212f
C9715 a_53660_14136# VPWR 0.31389f
C9716 _242_.Z a_58140_26680# 0.05801f
C9717 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN a_64100_27912# 0.05499f
C9718 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN 0.86967f
C9719 a_55028_12232# VPWR 0.20622f
C9720 a_43492_15748# a_43132_15704# 0.08707f
C9721 a_6308_29860# a_6172_29383# 0.00168f
C9722 a_47972_2824# a_48420_2824# 0.01328f
C9723 a_2364_29816# a_2364_29383# 0.05841f
C9724 a_28679_24776# VPWR 0.00667f
C9725 a_38676_20452# a_38316_20408# 0.08674f
C9726 _474_.D a_51240_19624# 0.0206f
C9727 a_27668_31048# _340_.A2 0.00936f
C9728 a_8636_2727# a_8548_2824# 0.28563f
C9729 a_49988_15748# VPWR 0.21606f
C9730 _474_.CLK _251_.A1 0.04382f
C9731 _448_.D a_36076_18407# 0.00413f
C9732 _442_.ZN a_40132_26344# 0.03112f
C9733 a_53660_21543# a_54108_21543# 0.01255f
C9734 _324_.C _411_.A2 0.087f
C9735 a_49540_9476# a_49180_9432# 0.08717f
C9736 a_50884_9476# a_51332_9476# 0.01328f
C9737 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN _249_.A2 0.03478f
C9738 _461_.D a_32848_29123# 0.00472f
C9739 a_53660_14136# a_54108_14136# 0.0131f
C9740 a_57156_14180# a_57244_14136# 0.28563f
C9741 _459_.CLK a_22064_27912# 0.07646f
C9742 a_35204_31048# a_35652_31048# 0.01328f
C9743 _452_.CLK a_37892_26344# 0.00546f
C9744 vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I VPWR 0.95416f
C9745 a_58836_18884# vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN 0.00413f
C9746 a_11100_1592# a_11236_1256# 0.00168f
C9747 a_58836_13800# a_58948_12612# 0.02666f
C9748 a_55028_13800# a_55004_12568# 0.0016f
C9749 _417_.Z a_49896_18909# 0.00117f
C9750 a_2276_24776# a_2276_23588# 0.05841f
C9751 a_30948_23208# a_30836_22020# 0.02666f
C9752 _355_.C a_22636_29383# 0.00625f
C9753 a_35652_26344# VPWR 0.20348f
C9754 a_10876_1159# VPWR 0.33578f
C9755 a_39548_1159# a_39908_1256# 0.08717f
C9756 a_932_6340# a_1380_6340# 0.01328f
C9757 a_55028_12232# a_55476_12232# 0.01328f
C9758 a_31844_26344# a_31820_25112# 0.0016f
C9759 a_23868_1592# a_24452_1636# 0.01675f
C9760 a_39796_22504# VPWR 1.3342f
C9761 a_4852_21640# VPWR 0.22733f
C9762 a_64100_27912# VPWR 0.1979f
C9763 a_51332_17316# a_50972_17272# 0.08707f
C9764 _350_.A2 a_29232_29931# 0.07439f
C9765 _473_.Q a_47860_21640# 0.01236f
C9766 _325_.A1 _304_.ZN 0.00341f
C9767 a_45372_10567# a_45284_10664# 0.28563f
C9768 _287_.A2 _337_.ZN 0.03127f
C9769 _290_.ZN _359_.B 0.754f
C9770 _287_.A1 _365_.ZN 0.02241f
C9771 _334_.A1 _296_.ZN 0.03805f
C9772 a_33276_23111# a_33188_23208# 0.28563f
C9773 a_63404_23111# VPWR 0.29679f
C9774 _459_.CLK a_27588_26724# 0.03028f
C9775 a_33152_22091# a_33540_22505# 0.00393f
C9776 _316_.ZN a_34715_22137# 0.00511f
C9777 _337_.A3 _336_.A1 0.07865f
C9778 a_2364_6296# VPWR 0.30029f
C9779 a_2364_23544# VPWR 0.30029f
C9780 a_61860_9476# VPWR 0.20595f
C9781 a_54420_21976# a_54824_22045# 0.41635f
C9782 _252_.ZN vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN 0.00128f
C9783 a_1468_13703# VPWR 0.29679f
C9784 a_15244_21543# a_15604_21640# 0.08717f
C9785 a_4156_3160# VPWR 0.30552f
C9786 a_54804_26724# a_54444_26680# 0.0869f
C9787 _251_.A1 _247_.ZN 0.00107f
C9788 a_43296_28733# _330_.A1 0.00211f
C9789 _350_.A2 _335_.ZN 0.4479f
C9790 _424_.A2 a_46476_20937# 0.0066f
C9791 _424_.B2 a_52204_18407# 0.02248f
C9792 a_4604_11000# VPWR 0.33016f
C9793 a_46404_15748# a_46492_15704# 0.28563f
C9794 _435_.ZN a_39332_23588# 0.00183f
C9795 _441_.ZN _438_.ZN 0.00326f
C9796 a_49988_15748# a_50436_15748# 0.01328f
C9797 a_36548_25156# VPWR 0.20348f
C9798 a_47768_20569# VPWR 0.00204f
C9799 a_66092_19975# a_66452_20072# 0.0869f
C9800 _397_.A2 _381_.Z 0.32803f
C9801 _275_.A2 a_51791_30644# 0.00258f
C9802 _331_.ZN _452_.D 0.10149f
C9803 _474_.CLK a_53996_18407# 0.00616f
C9804 a_31260_18840# VPWR 0.29679f
C9805 a_5388_26247# VPWR 0.35526f
C9806 a_67741_30600# ena 0.47748f
C9807 a_19388_2727# a_19972_2824# 0.01675f
C9808 _359_.B a_37396_29860# 0.0015f
C9809 _452_.Q _305_.A2 0.19709f
C9810 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I 0.65511f
C9811 _416_.A1 a_46352_22021# 0.00379f
C9812 a_37386_31048# uo_out[1] 0.00107f
C9813 _267_.A2 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN 0.02905f
C9814 _462_.D uo_out[3] 0.00681f
C9815 _324_.C _399_.ZN 1.64482f
C9816 a_1468_9432# a_1468_8999# 0.05841f
C9817 _416_.A1 _441_.A2 0.00202f
C9818 _475_.D a_47860_21640# 0.0016f
C9819 a_61860_14180# a_61948_14136# 0.28563f
C9820 a_51196_14136# a_51084_13703# 0.02634f
C9821 a_27564_21976# a_27476_20452# 0.00151f
C9822 _379_.Z uio_out[7] 0.24551f
C9823 _474_.Q a_50212_20452# 0.02438f
C9824 _459_.Q a_31844_26344# 0.00437f
C9825 a_52452_24072# a_52660_24072# 0.00334f
C9826 _250_.ZN a_60916_29612# 0.00177f
C9827 a_65780_13800# a_65892_12612# 0.02666f
C9828 a_49404_12568# a_49852_12568# 0.01288f
C9829 _438_.ZN a_39873_21236# 0.00631f
C9830 _474_.CLK a_55452_21543# 0.04081f
C9831 a_50972_1159# a_50884_1256# 0.28563f
C9832 _402_.ZN _284_.B 0.06024f
C9833 a_19972_24776# a_20084_23588# 0.02666f
C9834 a_33276_1159# VPWR 0.29975f
C9835 a_59820_12135# a_59844_11044# 0.0016f
C9836 a_31172_1636# a_30812_1592# 0.08707f
C9837 a_35652_26344# a_36100_26344# 0.01328f
C9838 a_35816_21192# VPWR 0.30379f
C9839 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I 0.00848f
C9840 a_62284_23544# VPWR 0.33401f
C9841 _267_.A1 a_52891_28776# 0.00943f
C9842 a_10876_1159# a_11324_1159# 0.0131f
C9843 a_56012_10567# a_56372_10664# 0.08663f
C9844 a_2276_10664# a_2724_10664# 0.01328f
C9845 a_3260_21976# VPWR 0.30487f
C9846 _355_.C a_25524_26344# 0.00165f
C9847 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN 0.10165f
C9848 _402_.A1 a_43044_27912# 0.00546f
C9849 a_36544_24419# a_37179_24831# 0.02112f
C9850 a_35616_24776# a_37472_24419# 0.02307f
C9851 a_31844_23208# a_32292_23208# 0.01328f
C9852 a_54780_18840# a_54804_18504# 0.00172f
C9853 _229_.I vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I 0.13999f
C9854 a_39796_22504# a_40452_22504# 0.01436f
C9855 _424_.B1 _417_.A2 0.8727f
C9856 _352_.ZN a_27172_24328# 0.02866f
C9857 a_25236_23588# VPWR 0.20614f
C9858 a_932_9096# VPWR 0.22176f
C9859 a_4852_21640# a_5300_21640# 0.01328f
C9860 a_26556_21543# a_26468_21640# 0.28563f
C9861 _467_.D a_16052_28292# 0.00857f
C9862 a_62956_13703# VPWR 0.31556f
C9863 a_1828_18884# a_1916_18840# 0.28563f
C9864 a_13340_2727# VPWR 0.31143f
C9865 a_40804_2824# a_40892_1159# 0.0027f
C9866 _419_.A4 _416_.A3 0.40202f
C9867 _459_.CLK a_31920_29480# 0.0721f
C9868 _355_.C a_22548_28292# 0.02058f
C9869 _324_.B a_43668_19668# 0.13536f
C9870 a_67237_31198# VPWR 0.00423f
C9871 _304_.B a_54804_26724# 0.00502f
C9872 a_49852_30951# a_49112_29885# 0.00101f
C9873 a_49404_30951# a_49600_30180# 0.00105f
C9874 a_58052_11044# VPWR 0.2284f
C9875 _371_.A3 a_27588_26724# 0.01448f
C9876 a_20756_26724# VPWR 0.20799f
C9877 _474_.Q a_51240_19624# 0.00555f
C9878 a_64772_15748# a_64412_15704# 0.08717f
C9879 a_67460_15748# a_67908_15748# 0.01328f
C9880 a_2812_27815# VPWR 0.30213f
C9881 _416_.A3 a_46940_17272# 0.00118f
C9882 _330_.A1 a_34644_20072# 0.00356f
C9883 a_63616_31128# vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.01938f
C9884 a_63404_23111# a_63852_23111# 0.0131f
C9885 a_30812_2727# a_30724_2824# 0.28563f
C9886 a_48084_18884# a_48172_18840# 0.28563f
C9887 a_4964_23588# a_4604_23544# 0.08674f
C9888 a_2364_23544# a_2812_23544# 0.0131f
C9889 a_59932_9432# a_60604_9432# 0.00544f
C9890 a_11684_1256# a_12356_1256# 0.00347f
C9891 _384_.ZN _397_.Z 0.00401f
C9892 a_61860_9476# a_62308_9476# 0.01328f
C9893 a_4068_7908# a_3708_7864# 0.08717f
C9894 a_1468_7864# a_1916_7864# 0.0131f
C9895 a_2364_6296# a_2812_6296# 0.0131f
C9896 a_4964_6340# a_4604_6296# 0.08674f
C9897 a_17732_31048# a_18180_31048# 0.01328f
C9898 _325_.A2 a_39236_20072# 0.00875f
C9899 rst_n clk 0.02969f
C9900 a_58924_14136# a_58924_13703# 0.05841f
C9901 a_3260_4728# a_3708_4728# 0.0131f
C9902 a_4156_3160# a_4604_3160# 0.01222f
C9903 a_1468_13703# a_1916_13703# 0.0131f
C9904 a_19860_20452# a_19948_20408# 0.28563f
C9905 a_2364_29383# a_2812_29383# 0.0131f
C9906 a_58687_31220# ui_in[3] 0.01058f
C9907 a_3260_30951# a_3172_31048# 0.28563f
C9908 a_6844_1592# VPWR 0.3289f
C9909 a_56708_12612# a_56348_12568# 0.08707f
C9910 _459_.CLK a_17484_25112# 0.00189f
C9911 a_59284_13800# a_59372_12135# 0.00151f
C9912 a_3260_12568# a_3260_12135# 0.05841f
C9913 _302_.Z a_42778_21812# 0.01919f
C9914 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_62060_23111# 0.009f
C9915 _330_.A1 _317_.A2 0.63624f
C9916 _416_.A2 a_47028_18884# 0.01232f
C9917 a_61164_20408# VPWR 0.31512f
C9918 a_55676_1159# VPWR 0.32824f
C9919 _416_.ZN a_46252_19759# 0.25445f
C9920 a_45696_20072# a_47259_20127# 0.41635f
C9921 a_4604_11000# a_5052_11000# 0.01222f
C9922 a_66764_12135# a_66788_11044# 0.0016f
C9923 a_61948_1159# a_62308_1256# 0.08717f
C9924 a_2276_16936# a_2724_16936# 0.01328f
C9925 a_34084_1636# a_34172_1592# 0.28563f
C9926 a_37668_1636# a_38116_1636# 0.01328f
C9927 a_36548_25156# a_36996_25156# 0.01328f
C9928 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN a_67772_24679# 0.00396f
C9929 a_64412_18840# VPWR 0.29986f
C9930 _441_.ZN a_39332_23588# 0.0015f
C9931 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN clk 0.04025f
C9932 _454_.Q a_25796_27912# 0.0021f
C9933 a_40692_27912# a_41140_27912# 0.01328f
C9934 _474_.Q _475_.Q 1.13539f
C9935 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN _245_.I1 0.98343f
C9936 a_44028_27815# _330_.A1 0.00843f
C9937 a_44476_27815# a_44388_27912# 0.28563f
C9938 a_62532_1636# a_62396_1159# 0.00168f
C9939 a_58588_1592# a_58588_1159# 0.05841f
C9940 a_67212_10567# a_67124_10664# 0.28563f
C9941 _467_.D a_16948_27912# 0.02026f
C9942 _244_.Z _245_.I1 0.00139f
C9943 a_32516_18504# a_32516_17316# 0.05841f
C9944 a_32240_31048# VPWR 0.6615f
C9945 _287_.A2 a_30795_29977# 0.0437f
C9946 a_26132_22020# VPWR 0.21332f
C9947 _397_.A2 _383_.A2 0.19387f
C9948 a_57044_13800# VPWR 0.23066f
C9949 a_31260_18840# a_31708_18840# 0.0131f
C9950 a_35740_2727# VPWR 0.31143f
C9951 a_33412_18884# a_33500_18840# 0.28563f
C9952 _284_.ZN _416_.A1 0.1727f
C9953 _427_.B1 _478_.D 0.77434f
C9954 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN a_56484_29480# 0.00767f
C9955 a_12356_29860# VPWR 0.20804f
C9956 a_54804_26724# VPWR 0.20698f
C9957 a_63092_16936# a_62980_15748# 0.02666f
C9958 _350_.A2 a_30596_28292# 0.01126f
C9959 _334_.A1 _335_.ZN 1.62203f
C9960 _381_.Z _330_.A1 0.02065f
C9961 a_64636_11000# VPWR 0.33474f
C9962 a_2812_15271# a_3172_15368# 0.08717f
C9963 vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN a_64860_26247# 0.0053f
C9964 ui_in[1] ui_in[0] 0.07726f
C9965 a_63404_23544# a_63404_23111# 0.05841f
C9966 a_23196_23111# VPWR 0.31547f
C9967 _247_.ZN a_58020_27508# 0.00785f
C9968 _349_.A4 _455_.Q 0.01944f
C9969 _378_.I VPWR 0.9863f
C9970 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I 0.00324f
C9971 _285_.Z a_39300_29480# 0.00162f
C9972 a_41788_2727# a_42148_2824# 0.08717f
C9973 a_28000_29480# a_29856_29123# 0.02307f
C9974 a_28928_29123# a_29563_29535# 0.02112f
C9975 a_64076_16839# a_63988_16936# 0.28563f
C9976 _260_.A1 a_40468_25157# 0.11045f
C9977 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN a_67772_24679# 0.04806f
C9978 _281_.ZN a_51332_24072# 0.03104f
C9979 a_18740_23588# a_18380_23544# 0.08707f
C9980 a_62172_18407# a_62620_18407# 0.0131f
C9981 a_67460_9476# a_67548_9432# 0.28563f
C9982 a_3620_25156# a_3260_25112# 0.08717f
C9983 a_61164_20408# a_61188_20072# 0.00172f
C9984 a_1020_25112# a_1468_25112# 0.0131f
C9985 a_66900_20072# a_67012_18884# 0.02666f
C9986 a_55452_14136# a_55476_13800# 0.00172f
C9987 _381_.A2 clk 0.00561f
C9988 a_25100_20408# a_25548_20408# 0.0131f
C9989 a_17820_30951# a_18180_31048# 0.0869f
C9990 _350_.A1 a_33508_31048# 0.00169f
C9991 a_67548_17272# a_67436_16839# 0.02634f
C9992 a_20644_1636# VPWR 0.2085f
C9993 a_58140_11000# a_58052_9476# 0.00151f
C9994 a_63204_12612# a_63652_12612# 0.01328f
C9995 _274_.A3 a_52964_29480# 0.00134f
C9996 _417_.A2 _218_.ZN 0.10204f
C9997 a_62620_15271# a_62980_15368# 0.08717f
C9998 a_32516_18504# VPWR 0.20348f
C9999 a_51556_11044# a_51196_11000# 0.08707f
C10000 a_9220_1636# a_9084_1159# 0.00168f
C10001 a_63764_12232# a_63652_11044# 0.02666f
C10002 _272_.B1 _274_.A2 0.04776f
C10003 _336_.A1 a_27328_25227# 0.04379f
C10004 hold1.Z a_44162_24120# 0.0486f
C10005 _330_.A1 _434_.ZN 0.19343f
C10006 a_932_26724# a_1020_26680# 0.28563f
C10007 a_63764_10664# a_64212_10664# 0.01328f
C10008 a_31920_29480# uo_out[7] 0.01124f
C10009 a_67884_18407# a_67908_17316# 0.0016f
C10010 a_33276_1159# a_33724_1159# 0.0131f
C10011 a_41476_24776# VPWR 0.171f
C10012 a_30276_2824# a_30276_1636# 0.05841f
C10013 a_26468_2824# a_26332_1592# 0.00154f
C10014 a_25796_24776# a_25884_23111# 0.00151f
C10015 _324_.C a_55140_28292# 0.00196f
C10016 a_65072_29860# VPWR 1.0503f
C10017 _379_.A2 a_21652_29480# 0.00424f
C10018 _355_.C a_26954_28776# 0.00229f
C10019 a_40132_26344# _441_.ZN 0.01462f
C10020 a_46180_12612# VPWR 0.20348f
C10021 a_58140_2727# VPWR 0.35834f
C10022 a_63204_2824# a_63292_1159# 0.0027f
C10023 a_35816_21192# a_36636_21543# 0.00481f
C10024 _470_.Q _404_.A1 0.89263f
C10025 a_64860_18407# a_65220_18504# 0.08663f
C10026 _460_.Q _223_.ZN 0.00554f
C10027 a_1020_29383# a_932_29480# 0.28563f
C10028 a_1828_20072# VPWR 0.20348f
C10029 a_37220_15368# a_37668_15368# 0.01328f
C10030 _346_.B a_19328_28733# 0.03616f
C10031 _399_.ZN _281_.A1 0.00106f
C10032 a_1020_15704# a_1020_15271# 0.05841f
C10033 a_58924_10567# VPWR 0.31389f
C10034 a_39324_15271# a_39236_15368# 0.28563f
C10035 a_20868_23208# VPWR 0.20595f
C10036 a_60401_30300# ui_in[2] 0.00481f
C10037 _304_.B _274_.A2 0.04278f
C10038 a_40668_15271# a_41116_15271# 0.0131f
C10039 _397_.A2 _324_.C 0.18863f
C10040 a_4964_28292# a_5052_28248# 0.28563f
C10041 _330_.A1 a_36772_23208# 0.00754f
C10042 _288_.ZN uo_out[2] 1.91482f
C10043 _427_.ZN a_55004_21543# 0.01267f
C10044 a_58687_31220# _267_.A2 0.00754f
C10045 a_3260_21976# a_3708_21976# 0.0131f
C10046 a_53212_2727# a_53124_2824# 0.28563f
C10047 a_64860_17272# a_65308_17272# 0.0131f
C10048 a_32380_26247# VPWR 0.32953f
C10049 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN a_58500_21640# 0.00636f
C10050 a_19076_23208# a_19164_21543# 0.00151f
C10051 a_25236_23588# a_25684_23588# 0.01328f
C10052 a_21964_23544# a_22636_23544# 0.00544f
C10053 a_17396_25156# a_17036_25112# 0.08707f
C10054 a_932_31048# VPWR 0.22176f
C10055 a_34084_1256# a_34532_1256# 0.01328f
C10056 a_3708_18840# a_3708_18407# 0.05841f
C10057 _435_.A3 _432_.ZN 0.01334f
C10058 a_30836_20452# a_30924_20408# 0.28563f
C10059 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN 0.00136f
C10060 a_49292_13703# a_49652_13800# 0.08707f
C10061 a_62956_13703# a_63404_13703# 0.01288f
C10062 a_13340_2727# a_13788_2727# 0.0131f
C10063 _438_.A2 _444_.D 0.07857f
C10064 _317_.A2 a_35723_20569# 0.0138f
C10065 a_36076_16839# a_36436_16936# 0.08707f
C10066 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN 0.02372f
C10067 a_53324_10567# a_53348_9476# 0.0016f
C10068 a_66787_30600# vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN 0.03008f
C10069 a_26780_1592# VPWR 0.339f
C10070 _460_.Q a_32592_25227# 0.00124f
C10071 a_17820_30951# a_18268_30951# 0.01255f
C10072 _284_.B a_46068_25156# 0.01f
C10073 _350_.A2 _223_.I 0.08758f
C10074 a_2364_25112# a_2364_24679# 0.05841f
C10075 a_67741_30600# a_67861_31220# 0.00165f
C10076 _473_.Q a_47483_20569# 0.00633f
C10077 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN a_60064_25156# 0.00179f
C10078 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN 0.00707f
C10079 a_49204_16936# a_49652_16936# 0.01328f
C10080 a_43804_1592# a_44252_1592# 0.01288f
C10081 a_54468_11044# a_54556_11000# 0.28563f
C10082 a_58052_11044# a_58500_11044# 0.01328f
C10083 a_5052_9432# a_4964_7908# 0.00151f
C10084 a_43344_19001# VPWR 0.00204f
C10085 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN 0.002f
C10086 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.00549f
C10087 a_2812_27815# a_3260_27815# 0.0131f
C10088 a_4604_29816# a_4516_28292# 0.0027f
C10089 a_21204_20452# VPWR 0.20677f
C10090 a_59844_12612# VPWR 0.20703f
C10091 _388_.B _397_.A1 0.00776f
C10092 a_14148_2824# a_14596_2824# 0.01328f
C10093 a_11772_29383# a_12356_29480# 0.01675f
C10094 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN VPWR 0.74446f
C10095 a_52788_10664# VPWR 0.20614f
C10096 vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN 0.00365f
C10097 a_36996_15748# a_36860_15271# 0.00168f
C10098 a_33052_15704# a_33052_15271# 0.05841f
C10099 a_54444_26680# a_54356_25156# 0.00151f
C10100 a_50300_15271# a_50660_15368# 0.08717f
C10101 a_2364_5863# a_2276_5960# 0.28563f
C10102 a_1468_7431# a_1380_7528# 0.28563f
C10103 a_52764_27815# a_52676_27912# 0.28563f
C10104 a_3260_4295# a_3172_4392# 0.28563f
C10105 a_1828_21640# a_1828_20452# 0.05841f
C10106 a_37084_26680# a_37532_26680# 0.01255f
C10107 _274_.A2 VPWR 0.31925f
C10108 _389_.ZN a_47924_28292# 0.00183f
C10109 _223_.I a_31516_28292# 0.00214f
C10110 a_932_15368# VPWR 0.22176f
C10111 a_55340_25112# clk 0.00335f
C10112 a_19636_22020# a_19276_21976# 0.08707f
C10113 a_64188_2727# a_64548_2824# 0.08717f
C10114 _416_.A1 a_39772_26247# 0.00549f
C10115 a_4156_15271# VPWR 0.3269f
C10116 a_48508_30951# a_48868_31048# 0.08717f
C10117 a_42778_21812# a_43814_21236# 0.00389f
C10118 a_60740_26724# VPWR 0.1524f
C10119 a_13788_29383# uio_oe[2] 0.0027f
C10120 a_28928_29123# VPWR 0.18818f
C10121 a_62084_17316# VPWR 0.22423f
C10122 a_29716_23588# a_29804_23544# 0.28563f
C10123 _325_.A2 a_39268_18840# 0.02834f
C10124 a_1020_4295# VPWR 0.30073f
C10125 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_57916_25112# 0.00221f
C10126 a_22660_1256# VPWR 0.20348f
C10127 a_66652_7864# VPWR 0.29679f
C10128 a_60268_13703# a_60180_13800# 0.28563f
C10129 a_13340_29383# VPWR 0.29679f
C10130 a_4828_30951# VPWR 0.31605f
C10131 a_40644_17272# a_40992_17433# 0.00277f
C10132 a_43232_29480# a_44795_29535# 0.41635f
C10133 a_47052_16839# a_46964_16936# 0.28563f
C10134 _470_.D a_43564_27209# 0.22603f
C10135 _480_.Q a_43788_29167# 0.24835f
C10136 a_65196_23544# vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN 0.00223f
C10137 _474_.CLK _409_.ZN 0.04799f
C10138 a_38228_16936# VPWR 0.20932f
C10139 a_40580_1636# VPWR 0.2085f
C10140 a_50188_12135# a_50636_12135# 0.01288f
C10141 a_5724_1159# a_6084_1256# 0.08717f
C10142 a_55340_24679# VPWR 0.29679f
C10143 a_67684_12612# a_67660_12135# 0.00172f
C10144 a_6844_1592# a_7292_1592# 0.01288f
C10145 _260_.A2 a_40468_25157# 0.00383f
C10146 a_5860_29860# a_5500_29816# 0.08707f
C10147 a_4604_20408# a_4516_18884# 0.0027f
C10148 _384_.ZN _284_.B 0.01847f
C10149 a_49404_30951# VPWR 0.31266f
C10150 a_68020_12232# a_68108_10567# 0.0027f
C10151 a_2724_2824# VPWR 0.20782f
C10152 a_51108_1636# a_50748_1592# 0.08707f
C10153 a_34980_22895# VPWR 0.31741f
C10154 _384_.A3 a_51428_23340# 0.00743f
C10155 _303_.ZN a_39684_20452# 0.00315f
C10156 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN a_64884_26724# 0.0126f
C10157 a_49180_15271# a_49316_14180# 0.00154f
C10158 a_3260_24679# a_3708_24679# 0.0131f
C10159 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I clk 0.0019f
C10160 _459_.CLK a_18716_26247# 0.01008f
C10161 a_50860_18407# a_50772_18504# 0.28563f
C10162 a_61164_20408# a_61612_20408# 0.01222f
C10163 a_55676_1159# a_56124_1159# 0.0131f
C10164 _325_.A1 _328_.A2 0.46163f
C10165 a_48868_18504# VPWR 0.21169f
C10166 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I a_56348_15271# 0.00151f
C10167 _441_.A3 a_40332_21543# 0.00154f
C10168 a_20532_25156# VPWR 0.20348f
C10169 a_64412_18840# a_64860_18840# 0.0131f
C10170 _352_.A2 a_28012_24679# 0.01116f
C10171 _397_.A4 _281_.ZN 0.7451f
C10172 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN a_59172_22020# 0.07299f
C10173 vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN 0.0982f
C10174 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN a_64860_19975# 0.00168f
C10175 a_17932_27815# a_17844_27912# 0.28563f
C10176 a_32180_20452# VPWR 0.20595f
C10177 a_21740_30951# VPWR 0.31143f
C10178 _343_.A2 _454_.Q 0.34566f
C10179 a_56260_31048# VPWR 0.21382f
C10180 _336_.Z VPWR 1.39286f
C10181 a_66428_12568# VPWR 0.32136f
C10182 a_32964_15748# a_33412_15748# 0.01328f
C10183 _416_.A2 a_45696_20072# 0.07375f
C10184 _475_.D a_46624_19715# 0.00263f
C10185 _470_.Q a_48384_26724# 0.0093f
C10186 _435_.A3 _260_.A1 0.2073f
C10187 a_19948_26680# uio_out[7] 0.00488f
C10188 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN a_63952_29480# 0.00393f
C10189 _398_.C _421_.A1 0.0235f
C10190 _447_.Q _324_.B 0.07631f
C10191 _324_.C _330_.A1 0.88849f
C10192 a_26556_21543# a_26580_20452# 0.0016f
C10193 _272_.B1 a_57500_30344# 0.00128f
C10194 a_1380_15748# VPWR 0.20348f
C10195 a_48196_15368# VPWR 0.20952f
C10196 a_47297_25596# a_47689_25156# 0.00762f
C10197 _352_.A2 a_29184_25597# 0.03093f
C10198 a_32240_31048# _370_.B 0.08934f
C10199 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_62844_27815# 0.02542f
C10200 a_22548_22020# a_22636_21976# 0.28563f
C10201 a_26132_22020# a_26580_22020# 0.01328f
C10202 a_44364_16839# a_44812_16839# 0.01288f
C10203 a_51644_15271# VPWR 0.32932f
C10204 _304_.B a_41392_27165# 0.05526f
C10205 a_33052_16839# VPWR 0.29736f
C10206 a_22636_30951# a_22548_31048# 0.28563f
C10207 a_45060_1256# VPWR 0.20348f
C10208 a_56484_1256# a_56932_1256# 0.01328f
C10209 a_57044_13800# a_57492_13800# 0.01328f
C10210 a_35740_2727# a_36188_2727# 0.0131f
C10211 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN 0.00571f
C10212 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN _248_.B1 0.25267f
C10213 a_40040_17675# a_40556_16839# 0.00138f
C10214 _454_.D a_22059_26399# 0.00177f
C10215 a_31620_17316# VPWR 0.20348f
C10216 a_59284_10664# a_59396_9476# 0.02666f
C10217 a_17148_1159# a_17060_1256# 0.28563f
C10218 a_47164_12135# a_47076_12232# 0.28563f
C10219 a_61052_12568# a_61076_12232# 0.00172f
C10220 a_54244_1636# VPWR 0.20348f
C10221 a_62396_27815# VPWR 0.31228f
C10222 _475_.Q a_51196_21543# 0.02873f
C10223 a_14148_1636# a_13788_1592# 0.08707f
C10224 a_66900_20072# a_66988_18407# 0.00151f
C10225 a_54804_26724# a_55252_26724# 0.01328f
C10226 a_12356_29860# a_12804_29860# 0.01328f
C10227 a_8772_29860# a_8860_29816# 0.28563f
C10228 a_57380_16936# vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I 0.03006f
C10229 a_34844_17272# a_35292_17272# 0.01288f
C10230 _336_.Z a_28903_24776# 0.10588f
C10231 a_48284_17272# a_48308_16936# 0.00172f
C10232 uio_out[5] uio_out[4] 0.1308f
C10233 _223_.I _334_.A1 0.18237f
C10234 a_25124_2824# VPWR 0.20815f
C10235 a_57604_1636# a_58052_1636# 0.01328f
C10236 _459_.CLK a_20396_26680# 0.01456f
C10237 a_64636_11000# a_65084_11000# 0.01288f
C10238 _301_.A1 _302_.Z 0.25493f
C10239 _334_.A1 _443_.D 0.00769f
C10240 _459_.CLK a_16140_27815# 0.00525f
C10241 a_1916_23111# a_2276_23208# 0.08717f
C10242 a_23196_23111# a_23644_23111# 0.01288f
C10243 _327_.A2 _328_.A2 0.64767f
C10244 a_14796_24679# a_15156_24776# 0.08717f
C10245 _234_.ZN a_40692_27912# 0.10639f
C10246 a_46180_14180# VPWR 0.20948f
C10247 a_6980_2824# a_7068_1159# 0.0027f
C10248 a_2364_18407# a_2276_18504# 0.28563f
C10249 VPWR uio_out[0] 0.05439f
C10250 a_33376_23659# a_34939_23705# 0.41635f
C10251 _330_.A2 a_38971_18559# 0.0588f
C10252 a_29232_29931# _370_.ZN 0.24439f
C10253 a_9892_29480# VPWR 0.20536f
C10254 a_60716_12135# VPWR 0.33016f
C10255 a_24316_2727# a_24452_1636# 0.00154f
C10256 a_36548_2824# a_36996_2824# 0.01328f
C10257 _274_.A3 _274_.A1 0.24459f
C10258 a_42796_23981# a_43246_24163# 0.00184f
C10259 a_47076_31048# VPWR 0.20348f
C10260 _474_.CLK a_55340_26680# 0.00457f
C10261 _229_.I _247_.B 0.00601f
C10262 _334_.A1 a_34260_29860# 0.00282f
C10263 vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN a_64972_26680# 0.0053f
C10264 a_58340_29860# VPWR 0.007f
C10265 a_23196_24679# VPWR 0.31589f
C10266 _452_.CLK a_38506_26724# 0.00269f
C10267 a_2724_7528# VPWR 0.20782f
C10268 a_35224_23705# VPWR 0.00235f
C10269 a_4852_4392# VPWR 0.22748f
C10270 a_45708_16839# a_45732_15748# 0.0016f
C10271 a_54356_25156# VPWR 0.20595f
C10272 a_35740_15704# VPWR 0.3289f
C10273 _424_.A2 a_51108_21640# 0.01372f
C10274 a_3708_9432# a_4156_9432# 0.0131f
C10275 a_38616_24328# _434_.ZN 0.00148f
C10276 a_4828_29383# a_4964_28292# 0.00154f
C10277 a_49404_14136# a_49852_14136# 0.01288f
C10278 a_51756_18407# VPWR 0.32205f
C10279 a_62980_15368# a_62844_14136# 0.00154f
C10280 a_41392_27165# VPWR 0.53259f
C10281 a_54892_16839# VPWR 0.32015f
C10282 _279_.Z VPWR 1.10458f
C10283 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN a_62508_21976# 0.00875f
C10284 a_67460_1256# VPWR 0.20348f
C10285 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN 0.13615f
C10286 _337_.A3 a_27676_26247# 0.02887f
C10287 _304_.B _304_.ZN 0.43323f
C10288 a_44632_30206# vgaringosc.workerclkbuff_notouch_.I 0.03351f
C10289 _346_.ZN a_21268_27912# 0.01477f
C10290 _334_.A1 a_32508_30644# 0.00117f
C10291 a_66676_10664# a_66564_9476# 0.02666f
C10292 a_64884_10664# a_64860_9432# 0.0016f
C10293 a_38842_17316# VPWR 0.01466f
C10294 _358_.A3 a_33148_25641# 0.01059f
C10295 a_60380_1592# VPWR 0.29679f
C10296 a_28124_1159# a_28484_1256# 0.08717f
C10297 a_17060_1636# a_17148_1592# 0.28563f
C10298 a_20644_1636# a_21092_1636# 0.01328f
C10299 a_55452_12568# a_55364_11044# 0.00151f
C10300 _346_.A2 a_21052_26031# 0.00291f
C10301 a_4068_12232# a_4852_12232# 0.00276f
C10302 a_58028_12135# a_58388_12232# 0.08707f
C10303 a_55956_25940# clk 0.00156f
C10304 a_16140_21543# VPWR 0.29679f
C10305 a_61948_11000# a_62060_10567# 0.02634f
C10306 a_47524_2824# VPWR 0.20839f
C10307 a_22300_23111# a_22212_23208# 0.28563f
C10308 a_16948_24776# a_17396_24776# 0.01328f
C10309 hold1.Z a_43814_21236# 0.01277f
C10310 a_25884_24679# a_25796_24776# 0.28563f
C10311 a_50436_9476# VPWR 0.25076f
C10312 _218_.ZN a_50644_21640# 0.00197f
C10313 a_58500_2824# a_58500_1636# 0.05841f
C10314 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN a_62756_27912# 0.00568f
C10315 a_50704_27912# VPWR 0.00825f
C10316 a_22548_31048# VPWR 0.20688f
C10317 a_53212_14136# VPWR 0.3185f
C10318 a_32516_18504# a_32964_18504# 0.01328f
C10319 _275_.ZN a_51665_30344# 0.00356f
C10320 _311_.Z a_35816_21192# 0.00124f
C10321 _294_.A2 a_35140_26680# 0.00181f
C10322 a_54580_12232# VPWR 0.20622f
C10323 a_43044_15748# a_43132_15704# 0.28563f
C10324 a_39100_15704# a_39548_15704# 0.01288f
C10325 a_38228_20452# a_38316_20408# 0.28563f
C10326 _248_.B1 a_64100_27912# 0.00151f
C10327 _467_.D a_17786_29480# 0.02598f
C10328 a_27004_30951# _340_.A2 0.00458f
C10329 a_52652_16839# a_52676_15748# 0.0016f
C10330 a_32292_21640# a_32268_20408# 0.0016f
C10331 a_7964_2727# a_8548_2824# 0.01675f
C10332 _417_.A2 a_51877_21236# 0.00137f
C10333 a_49540_15748# VPWR 0.21104f
C10334 a_24952_29032# _454_.Q 0.00714f
C10335 _474_.CLK a_56348_30951# 0.04414f
C10336 _384_.A3 a_49828_22020# 0.01909f
C10337 _442_.ZN a_39684_26344# 0.02111f
C10338 a_49092_9476# a_49180_9432# 0.28563f
C10339 _461_.D a_31920_29480# 0.24637f
C10340 _435_.A3 _260_.A2 0.03179f
C10341 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I 0.63235f
C10342 _452_.CLK a_37444_26344# 0.00546f
C10343 a_4156_14136# a_4156_13703# 0.05841f
C10344 a_57156_14180# a_56796_14136# 0.08674f
C10345 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I clk 0.00166f
C10346 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_64100_27912# 0.01676f
C10347 a_45484_28248# _400_.ZN 0.00887f
C10348 _258_.I _272_.A2 0.09941f
C10349 _384_.A1 _427_.B2 0.00964f
C10350 a_46180_12612# a_46628_12612# 0.01328f
C10351 a_58140_2727# a_58588_2727# 0.0131f
C10352 _304_.ZN VPWR 2.02478f
C10353 a_56932_23208# vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.00205f
C10354 a_35204_26344# VPWR 0.16518f
C10355 _355_.C a_22188_29383# 0.00613f
C10356 a_39548_1159# a_39460_1256# 0.28563f
C10357 _274_.A1 _324_.C 0.01042f
C10358 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN 0.10254f
C10359 a_10428_1159# VPWR 0.3335f
C10360 a_1828_20072# a_2276_20072# 0.01328f
C10361 a_4068_9096# a_4068_7908# 0.05841f
C10362 a_1380_12232# a_1380_11044# 0.05841f
C10363 _384_.ZN _474_.Q 0.06379f
C10364 a_4068_21640# VPWR 0.22146f
C10365 a_50884_17316# a_50972_17272# 0.28563f
C10366 a_46940_17272# a_47388_17272# 0.01288f
C10367 _230_.I vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.03205f
C10368 _409_.ZN _393_.A3 0.11095f
C10369 a_62756_27912# VPWR 0.20835f
C10370 _437_.A1 _301_.A1 0.00573f
C10371 _340_.A2 a_25252_30345# 0.0014f
C10372 a_58924_10567# a_59372_10567# 0.01288f
C10373 a_44252_1592# a_44252_1159# 0.05841f
C10374 a_66876_1592# a_67324_1592# 0.01222f
C10375 a_5188_2824# a_5052_1592# 0.00154f
C10376 a_36960_27912# a_37348_27599# 0.00393f
C10377 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN a_58028_13703# 0.00189f
C10378 a_20868_23208# a_21316_23208# 0.01328f
C10379 _459_.CLK a_27140_26724# 0.02059f
C10380 a_62956_23111# VPWR 0.31163f
C10381 a_32828_23111# a_33188_23208# 0.08707f
C10382 a_61412_9476# VPWR 0.20595f
C10383 a_33152_22091# a_34715_22137# 0.41635f
C10384 a_1916_23544# VPWR 0.297f
C10385 a_54040_22366# _427_.ZN 0.01687f
C10386 a_27452_21543# a_27900_21543# 0.01288f
C10387 a_15244_21543# a_15156_21640# 0.28563f
C10388 a_3172_29480# a_3172_28292# 0.05841f
C10389 a_4852_26344# a_4940_24679# 0.00151f
C10390 a_1916_6296# VPWR 0.297f
C10391 a_1020_13703# VPWR 0.30073f
C10392 a_3708_3160# VPWR 0.33374f
C10393 a_59955_30600# a_60405_31198# 0.00209f
C10394 a_54356_26724# a_54444_26680# 0.28563f
C10395 a_41996_28777# _330_.A1 0.0021f
C10396 _474_.CLK vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN 0.00134f
C10397 _424_.A2 a_46848_20893# 0.00775f
C10398 a_21740_29383# uio_out[5] 0.0012f
C10399 a_36100_25156# VPWR 0.20348f
C10400 a_4156_11000# VPWR 0.30552f
C10401 a_45820_15704# a_46492_15704# 0.00544f
C10402 a_58948_2824# a_59396_2824# 0.01328f
C10403 a_46820_20569# VPWR 0.00246f
C10404 _393_.ZN _404_.A1 0.01005f
C10405 a_9084_30951# a_9220_29860# 0.00154f
C10406 a_66092_19975# a_66004_20072# 0.28563f
C10407 _331_.ZN a_41776_18504# 0.01553f
C10408 _474_.CLK a_53548_18407# 0.00711f
C10409 a_30812_18840# VPWR 0.30073f
C10410 a_50704_27912# a_50068_27508# 0.02745f
C10411 _304_.A1 _312_.ZN 1.40839f
C10412 a_67117_30600# ena 0.07449f
C10413 a_4940_26247# VPWR 0.31945f
C10414 _359_.B a_36948_29860# 0.00249f
C10415 a_19388_2727# a_19300_2824# 0.28563f
C10416 a_32380_26247# _360_.ZN 0.06386f
C10417 _452_.Q a_42084_24072# 0.00127f
C10418 a_36288_31048# uo_out[3] 0.00254f
C10419 _334_.A1 a_37584_29123# 0.33867f
C10420 a_54332_9432# a_54780_9432# 0.0131f
C10421 a_56036_9476# a_56708_9476# 0.00347f
C10422 _304_.B a_44340_26183# 0.05089f
C10423 a_932_31048# a_1380_31048# 0.01328f
C10424 a_64996_14180# a_65444_14180# 0.01328f
C10425 a_61860_14180# a_61500_14136# 0.08707f
C10426 a_47271_21640# a_47860_21640# 0.08978f
C10427 _474_.Q a_49068_20408# 0.28468f
C10428 _330_.A1 a_38852_18884# 0.00233f
C10429 _250_.ZN a_60656_29612# 0.00468f
C10430 _455_.Q a_25124_28776# 0.07533f
C10431 _452_.CLK _319_.A3 0.05163f
C10432 a_61972_13800# a_61948_12568# 0.0016f
C10433 _268_.A1 _267_.ZN 0.13719f
C10434 _438_.ZN a_39669_21236# 0.00263f
C10435 a_6308_29860# uio_oe[7] 0.00193f
C10436 _433_.ZN a_41440_23208# 0.00218f
C10437 _325_.A2 a_43664_17317# 0.10898f
C10438 a_32828_1159# VPWR 0.29679f
C10439 a_50524_1159# a_50884_1256# 0.08717f
C10440 _474_.CLK a_55004_21543# 0.03075f
C10441 a_26780_1592# a_27228_1592# 0.01288f
C10442 a_30724_1636# a_30812_1592# 0.28563f
C10443 a_65780_12232# a_66228_12232# 0.01328f
C10444 a_49652_12232# a_49764_11044# 0.02666f
C10445 a_35268_21640# VPWR 0.00734f
C10446 _268_.A1 _390_.ZN 0.0017f
C10447 a_39772_26247# _431_.A3 0.00236f
C10448 _452_.Q a_41216_23208# 0.01348f
C10449 a_61836_23544# VPWR 0.33492f
C10450 a_56012_10567# a_55924_10664# 0.28563f
C10451 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN a_53212_27815# 0.0036f
C10452 _452_.Q _325_.A1 0.33462f
C10453 _355_.C a_25300_26344# 0.01623f
C10454 a_2812_21976# VPWR 0.30213f
C10455 _402_.A1 a_42596_27912# 0.00222f
C10456 a_35616_24776# a_37179_24831# 0.41635f
C10457 a_36544_24419# a_36172_24463# 0.10745f
C10458 _251_.A1 _251_.ZN 0.68375f
C10459 a_65756_23111# vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN 0.05734f
C10460 a_67548_8999# VPWR 0.32135f
C10461 a_3620_18884# a_4068_18884# 0.01328f
C10462 _352_.ZN a_25884_24679# 0.01516f
C10463 a_24788_23588# VPWR 0.20597f
C10464 a_1828_18884# a_1468_18840# 0.08717f
C10465 a_25884_21543# a_26468_21640# 0.01675f
C10466 a_12892_2727# VPWR 0.31143f
C10467 a_16612_29480# a_16500_28292# 0.02666f
C10468 a_62508_13703# VPWR 0.31556f
C10469 _383_.A2 _393_.A1 0.52018f
C10470 _467_.D a_15604_28292# 0.0036f
C10471 _355_.C a_21628_28248# 0.03576f
C10472 _438_.A2 _436_.ZN 0.00182f
C10473 a_51084_28248# _408_.ZN 0.00958f
C10474 _443_.D a_37532_26680# 0.01201f
C10475 a_67741_30600# VPWR 0.77946f
C10476 _304_.B a_54356_26724# 0.00449f
C10477 a_52764_15704# a_53212_15704# 0.01288f
C10478 a_57604_11044# VPWR 0.21273f
C10479 _359_.B _373_.ZN 0.01548f
C10480 _459_.CLK _379_.Z 0.01907f
C10481 a_20308_26724# VPWR 0.20348f
C10482 _255_.I _247_.ZN 0.00511f
C10483 _474_.Q a_48776_20204# 0.41502f
C10484 _462_.D a_36284_29167# 0.21102f
C10485 a_36100_26344# a_36100_25156# 0.05841f
C10486 a_64324_15748# a_64412_15704# 0.28563f
C10487 a_2364_27815# VPWR 0.30029f
C10488 a_30364_2727# a_30724_2824# 0.08717f
C10489 a_64412_3160# a_64548_2824# 0.00168f
C10490 a_48084_18884# a_47724_18840# 0.08674f
C10491 a_44340_26183# VPWR 0.35524f
C10492 _416_.A1 _470_.D 0.04293f
C10493 _325_.A2 a_38788_20072# 0.00876f
C10494 a_4516_23588# a_4604_23544# 0.28563f
C10495 a_3620_7908# a_3708_7864# 0.28563f
C10496 a_4516_6340# a_4604_6296# 0.28563f
C10497 a_7540_31048# a_7516_29383# 0.00134f
C10498 _448_.Q a_38576_22504# 0.04584f
C10499 a_19860_20452# a_19500_20408# 0.08717f
C10500 a_21204_20452# a_21652_20452# 0.01328f
C10501 a_2812_30951# a_3172_31048# 0.08717f
C10502 a_6396_1592# VPWR 0.3289f
C10503 a_24988_1592# a_25124_1256# 0.00168f
C10504 a_59844_12612# a_60292_12612# 0.01328f
C10505 _459_.CLK a_17036_25112# 0.00171f
C10506 a_56260_12612# a_56348_12568# 0.28563f
C10507 _330_.A1 a_36148_21976# 0.09159f
C10508 _419_.A4 _284_.A2 0.02554f
C10509 _402_.A1 _395_.A1 0.17953f
C10510 a_23556_24776# a_23532_23544# 0.0016f
C10511 _324_.B _421_.B 0.09309f
C10512 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_61612_23111# 0.05915f
C10513 a_55228_1159# VPWR 0.29679f
C10514 _371_.ZN _337_.A3 0.02851f
C10515 a_61948_1159# a_61860_1256# 0.28563f
C10516 _416_.ZN a_46624_19715# 0.04642f
C10517 a_45696_20072# a_46252_19759# 0.8399f
C10518 a_63964_18840# VPWR 0.29679f
C10519 a_34084_1636# a_33724_1592# 0.08707f
C10520 a_44028_27815# a_44388_27912# 0.08674f
C10521 a_43580_27815# _330_.A1 0.00424f
C10522 a_52408_19759# _424_.ZN 0.02083f
C10523 _467_.D a_16500_27912# 0.04646f
C10524 _452_.Q _327_.A2 0.58892f
C10525 a_52788_10664# a_53236_10664# 0.01328f
C10526 a_66764_10567# a_67124_10664# 0.08717f
C10527 a_21852_1159# a_22300_1159# 0.0131f
C10528 a_51791_30644# VPWR 0.6978f
C10529 a_25684_22020# VPWR 0.20903f
C10530 _355_.C a_22996_29480# 0.00148f
C10531 _258_.I _228_.ZN 0.02963f
C10532 _272_.A2 _255_.ZN 0.09259f
C10533 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN _231_.I 0.00102f
C10534 a_24452_21640# a_24900_21640# 0.01328f
C10535 a_33412_18884# a_33052_18840# 0.08717f
C10536 a_56372_13800# VPWR 0.21291f
C10537 _424_.A2 _417_.A2 0.64545f
C10538 a_35292_2727# VPWR 0.32369f
C10539 a_51780_2824# a_51868_1159# 0.0027f
C10540 a_40038_28720# _234_.ZN 0.81603f
C10541 a_932_15368# a_1380_15368# 0.01328f
C10542 a_54356_26724# VPWR 0.20348f
C10543 _459_.CLK uo_out[6] 0.05329f
C10544 a_11908_29860# VPWR 0.21787f
C10545 a_64188_11000# VPWR 0.31526f
C10546 a_2812_15271# a_2724_15368# 0.28563f
C10547 a_21516_21976# a_21404_21543# 0.02634f
C10548 _350_.A2 a_29575_28293# 0.02906f
C10549 a_22748_23111# VPWR 0.31547f
C10550 _459_.CLK a_28054_30196# 0.02643f
C10551 a_4156_15271# a_4940_15271# 0.00443f
C10552 _349_.A4 a_24392_28248# 0.00619f
C10553 a_66204_17272# a_66116_15748# 0.00151f
C10554 a_63316_23208# a_63764_23208# 0.01328f
C10555 a_41788_2727# a_41700_2824# 0.28563f
C10556 a_62084_17316# a_62532_17316# 0.01328f
C10557 a_28000_29480# a_29563_29535# 0.41635f
C10558 a_5052_23544# a_4964_22020# 0.00151f
C10559 a_28928_29123# a_28556_29167# 0.10745f
C10560 a_63628_16839# a_63988_16936# 0.08717f
C10561 _281_.ZN a_50940_24072# 0.00103f
C10562 a_65308_9432# a_65756_9432# 0.0131f
C10563 a_67460_9476# a_67100_9432# 0.08717f
C10564 a_66652_7864# a_67100_7864# 0.0131f
C10565 a_18292_23588# a_18380_23544# 0.28563f
C10566 a_22660_1256# a_23108_1256# 0.01328f
C10567 a_3172_25156# a_3260_25112# 0.28563f
C10568 a_67548_6296# a_67996_6296# 0.012f
C10569 a_64412_4728# a_64412_4295# 0.05841f
C10570 a_1020_4295# a_1468_4295# 0.0131f
C10571 a_65980_14136# a_65868_13703# 0.02634f
C10572 a_51980_13703# a_52428_13703# 0.01288f
C10573 a_1916_2727# a_2364_2727# 0.0131f
C10574 a_17820_30951# a_17732_31048# 0.28563f
C10575 a_41028_26344# a_41476_26344# 0.01328f
C10576 a_13340_29383# a_13788_29383# 0.0131f
C10577 _350_.A1 a_33060_31048# 0.00164f
C10578 a_20196_1636# VPWR 0.2085f
C10579 a_49852_12568# a_49740_12135# 0.02634f
C10580 a_4828_30951# a_5276_30951# 0.01255f
C10581 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I 0.08744f
C10582 _474_.CLK a_51620_19911# 0.0036f
C10583 _435_.A3 _311_.A2 0.00439f
C10584 a_17596_29816# _467_.D 0.0059f
C10585 a_47164_11000# a_47612_11000# 0.01288f
C10586 a_51108_11044# a_51196_11000# 0.28563f
C10587 a_62620_15271# a_62532_15368# 0.28563f
C10588 a_61412_17316# a_62084_17316# 0.00347f
C10589 a_38228_16936# a_38676_16936# 0.01328f
C10590 a_40580_1636# a_41028_1636# 0.01328f
C10591 a_32068_18504# VPWR 0.20348f
C10592 a_55340_24679# a_55788_24679# 0.01222f
C10593 _336_.A2 _355_.ZN 0.31224f
C10594 hold1.Z a_43750_23544# 0.06579f
C10595 a_51576_25896# a_52360_26355# 0.02307f
C10596 a_2724_26724# a_3172_26724# 0.01328f
C10597 _355_.C _359_.B 0.01923f
C10598 a_40973_24776# VPWR 0.00669f
C10599 _355_.C a_26750_28776# 0.00395f
C10600 a_39684_26344# _441_.ZN 0.00283f
C10601 a_36284_29167# a_36628_29535# 0.00275f
C10602 VPWR ui_in[2] 0.42839f
C10603 _403_.ZN a_45169_27509# 0.00488f
C10604 _274_.ZN a_52756_29076# 0.27543f
C10605 a_60516_26344# vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN 0.00104f
C10606 a_49404_30951# a_49852_30951# 0.0131f
C10607 a_57468_2727# VPWR 0.34658f
C10608 a_34980_22895# _311_.Z 0.22162f
C10609 a_45732_12612# VPWR 0.20348f
C10610 a_2724_2824# a_3172_2824# 0.01328f
C10611 a_14708_26344# a_15156_26344# 0.01328f
C10612 a_64860_18407# a_64772_18504# 0.28563f
C10613 _346_.B a_19035_28409# 0.00284f
C10614 a_1380_20072# VPWR 0.20348f
C10615 _438_.A2 _439_.ZN 0.08702f
C10616 a_28460_21976# a_28348_21543# 0.02634f
C10617 a_58476_10567# VPWR 0.32775f
C10618 _459_.CLK a_28891_25273# 0.02467f
C10619 a_38876_15271# a_39236_15368# 0.08717f
C10620 _287_.A1 VPWR 3.81081f
C10621 a_20420_23208# VPWR 0.20595f
C10622 a_29856_29123# _337_.ZN 0.02693f
C10623 vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN VPWR 0.76999f
C10624 _275_.A2 _268_.A1 0.52624f
C10625 _330_.A1 a_36288_23208# 0.01818f
C10626 _427_.ZN a_54556_21543# 0.01268f
C10627 a_54824_22045# vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I 0.00474f
C10628 a_4964_28292# a_4604_28248# 0.08674f
C10629 a_2364_28248# a_2812_28248# 0.0131f
C10630 a_52764_2727# a_53124_2824# 0.08717f
C10631 a_40668_20408# _325_.A2 0.00346f
C10632 a_18828_23544# a_18740_22020# 0.00151f
C10633 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN a_55364_21640# 0.00467f
C10634 a_31932_26247# VPWR 0.31599f
C10635 a_48868_18504# a_49316_18504# 0.01328f
C10636 _397_.A1 _402_.A1 0.11427f
C10637 a_20532_25156# a_20980_25156# 0.01328f
C10638 _350_.A2 _363_.Z 0.00342f
C10639 a_16948_25156# a_17036_25112# 0.28563f
C10640 a_49292_13703# a_49204_13800# 0.28563f
C10641 a_62844_14136# a_62868_13800# 0.00172f
C10642 a_32180_20452# a_32628_20452# 0.01328f
C10643 _352_.A2 _351_.A2 0.43329f
C10644 a_30836_20452# a_30476_20408# 0.08717f
C10645 _436_.B _325_.A1 0.00482f
C10646 a_37980_26247# _444_.D 0.00453f
C10647 a_21740_30951# a_22188_30951# 0.01255f
C10648 a_36076_16839# a_35988_16936# 0.28563f
C10649 _317_.A2 a_36016_20893# 0.0499f
C10650 a_51108_21640# a_49988_21236# 0.07589f
C10651 _373_.A2 _459_.CLK 0.52317f
C10652 a_63292_11000# a_63204_9476# 0.00151f
C10653 a_26332_1592# VPWR 0.33528f
C10654 a_3620_1636# a_4068_1636# 0.01328f
C10655 _352_.A2 a_29680_26724# 0.00948f
C10656 a_66428_12568# a_66876_12568# 0.01288f
C10657 _304_.B _328_.A2 0.00335f
C10658 _473_.Q a_47776_20893# 0.08726f
C10659 a_54468_11044# a_54108_11000# 0.08707f
C10660 a_57044_12232# a_57132_10567# 0.00151f
C10661 a_1020_11000# a_1020_10567# 0.05841f
C10662 a_47300_1636# a_47972_1636# 0.00347f
C10663 _324_.B a_47524_22021# 0.0244f
C10664 _474_.CLK _267_.ZN 0.00898f
C10665 a_49492_18840# a_49404_18407# 0.02951f
C10666 _474_.CLK vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.0323f
C10667 _246_.B2 a_59620_27208# 0.4116f
C10668 a_44252_1159# a_44700_1159# 0.0131f
C10669 _334_.A1 a_38584_28292# 0.00609f
C10670 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN a_64660_23588# 0.00102f
C10671 uo_out[7] uo_out[6] 0.12464f
C10672 a_3172_27912# a_3172_26724# 0.05841f
C10673 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I 0.05458f
C10674 a_48888_19243# VPWR 0.70085f
C10675 a_62084_18884# a_62532_18884# 0.01328f
C10676 a_51048_26680# _284_.A2 0.21683f
C10677 _260_.ZN _304_.ZN 0.17743f
C10678 _455_.D a_21052_26031# 0.2178f
C10679 _474_.CLK _390_.ZN 0.0053f
C10680 a_20756_20452# VPWR 0.20677f
C10681 _293_.A2 VPWR 1.05901f
C10682 a_28054_30196# uo_out[7] 0.0034f
C10683 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I a_61836_25515# 0.00366f
C10684 a_59396_12612# VPWR 0.20703f
C10685 a_1380_15748# a_1828_15748# 0.01328f
C10686 a_9980_2727# a_10116_1636# 0.00154f
C10687 a_11772_29383# a_11684_29480# 0.28563f
C10688 a_48196_15368# a_48644_15368# 0.01328f
C10689 _441_.B VPWR 1.06224f
C10690 _397_.A4 a_47636_25940# 0.00131f
C10691 a_58924_17272# vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I 0.00171f
C10692 a_16140_28248# a_16140_27815# 0.05841f
C10693 a_24864_29931# a_25744_30345# 0.00306f
C10694 a_1020_7431# a_1380_7528# 0.08717f
C10695 a_52340_10664# VPWR 0.20641f
C10696 a_50300_15271# a_50212_15368# 0.28563f
C10697 a_1916_5863# a_2276_5960# 0.08717f
C10698 a_52316_27815# a_52676_27912# 0.0869f
C10699 _244_.Z a_61836_26680# 0.00142f
C10700 a_4940_16839# a_4964_15748# 0.0016f
C10701 a_2812_4295# a_3172_4392# 0.08717f
C10702 _389_.ZN a_47700_28292# 0.0063f
C10703 a_44340_26183# a_44744_26355# 0.41635f
C10704 _470_.Q _411_.A2 0.08852f
C10705 _395_.A1 _424_.B1 0.14768f
C10706 a_51644_15271# a_52092_15271# 0.0131f
C10707 a_67772_15271# VPWR 0.34901f
C10708 a_19188_22020# a_19276_21976# 0.28563f
C10709 a_54892_25112# clk 0.00335f
C10710 _416_.A1 a_39324_26247# 0.00977f
C10711 a_15244_21976# a_15692_21976# 0.01288f
C10712 a_64188_2727# a_64100_2824# 0.28563f
C10713 a_3708_15271# VPWR 0.33374f
C10714 a_33052_16839# a_33500_16839# 0.0131f
C10715 a_48508_30951# a_48420_31048# 0.28563f
C10716 a_22636_23544# a_22548_22020# 0.00151f
C10717 a_42982_21730# a_43214_21812# 0.00212f
C10718 a_61500_17272# VPWR 0.34556f
C10719 a_28000_29480# VPWR 1.10142f
C10720 a_45060_1256# a_45508_1256# 0.01328f
C10721 _255_.ZN _228_.ZN 0.04437f
C10722 a_29604_23208# a_29692_21543# 0.00151f
C10723 a_22212_1256# VPWR 0.20348f
C10724 a_28820_24072# a_29804_23544# 0.00505f
C10725 a_67996_4728# VPWR 0.35142f
C10726 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_55788_25112# 0.02408f
C10727 a_66204_7864# VPWR 0.31657f
C10728 _325_.A2 a_37312_19369# 0.00111f
C10729 a_59820_13703# a_60180_13800# 0.08707f
C10730 a_56796_14136# a_56708_12612# 0.0027f
C10731 a_45732_13800# a_46180_13800# 0.01328f
C10732 a_24316_2727# a_24764_2727# 0.0131f
C10733 a_12892_29383# VPWR 0.29679f
C10734 a_4156_30951# VPWR 0.34855f
C10735 a_43232_29480# a_43788_29167# 0.8399f
C10736 _470_.D a_43936_27165# 0.023f
C10737 _480_.Q a_44160_29123# 0.01542f
C10738 a_46604_16839# a_46964_16936# 0.08707f
C10739 _474_.CLK a_49496_30345# 0.00923f
C10740 a_5724_1159# a_5636_1256# 0.28563f
C10741 a_51892_10664# a_51780_9476# 0.02666f
C10742 a_50100_10664# a_50076_9432# 0.0016f
C10743 a_40132_1636# VPWR 0.22925f
C10744 a_37780_16936# VPWR 0.2061f
C10745 a_63740_12568# a_63852_12135# 0.02634f
C10746 a_54892_24679# VPWR 0.29679f
C10747 uo_out[0] uo_out[3] 0.12785f
C10748 a_53660_12568# a_53684_12232# 0.00172f
C10749 _328_.A2 VPWR 0.54653f
C10750 a_5412_29860# a_5500_29816# 0.28563f
C10751 a_1468_29816# a_1916_29816# 0.01288f
C10752 a_31620_17316# a_32068_17316# 0.01328f
C10753 a_51556_11044# a_51532_10567# 0.00172f
C10754 a_47612_11000# a_47612_10567# 0.05841f
C10755 a_48956_30951# VPWR 0.3122f
C10756 a_61276_15271# a_61412_14180# 0.00154f
C10757 a_60964_11044# a_61412_11044# 0.01328f
C10758 a_2276_2824# VPWR 0.20634f
C10759 a_34586_23208# VPWR 0.01598f
C10760 a_50660_1636# a_50748_1592# 0.28563f
C10761 a_54244_1636# a_54692_1636# 0.01328f
C10762 a_62396_27815# a_62844_27815# 0.012f
C10763 _352_.A2 a_28756_25940# 0.00289f
C10764 a_31172_20072# a_31172_18884# 0.05841f
C10765 a_2812_23111# a_3260_23111# 0.0131f
C10766 a_11012_29860# uio_oe[4] 0.0033f
C10767 a_50412_18407# a_50772_18504# 0.08717f
C10768 _459_.CLK a_17932_26247# 0.00821f
C10769 a_52116_18504# a_52204_16839# 0.00151f
C10770 _251_.A1 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I 0.00277f
C10771 a_68108_20408# a_67908_18884# 0.00119f
C10772 a_40356_2824# a_40220_1592# 0.00154f
C10773 a_44164_2824# a_44164_1636# 0.05841f
C10774 a_48420_18504# VPWR 0.20897f
C10775 _352_.A2 a_27172_24328# 0.4988f
C10776 a_20084_25156# VPWR 0.20593f
C10777 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN a_64412_19975# 0.00479f
C10778 _432_.ZN _441_.A3 0.09375f
C10779 a_31732_20452# VPWR 0.20595f
C10780 a_3172_27912# a_3620_27912# 0.01328f
C10781 a_17484_27815# a_17844_27912# 0.08717f
C10782 _343_.A2 a_23084_28248# 0.00108f
C10783 a_21292_30951# VPWR 0.31267f
C10784 a_65980_12568# VPWR 0.36289f
C10785 a_25124_2824# a_25572_2824# 0.01328f
C10786 _412_.B2 a_51332_24372# 0.37631f
C10787 _284_.A2 _381_.A2 0.41401f
C10788 _395_.A2 a_51576_25896# 0.00644f
C10789 _284_.ZN a_43008_26795# 0.04213f
C10790 _324_.C a_44388_27912# 0.05966f
C10791 _267_.A2 a_52764_27815# 0.00123f
C10792 _300_.A2 VPWR 0.68288f
C10793 _304_.B a_53908_25156# 0.00225f
C10794 a_932_15748# VPWR 0.22176f
C10795 _355_.C uio_out[4] 0.00548f
C10796 _474_.CLK a_48580_27508# 0.0017f
C10797 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I uio_in[0] 0.0262f
C10798 _476_.Q _419_.Z 1.25694f
C10799 a_47748_15368# VPWR 0.20952f
C10800 _352_.A2 a_27884_25641# 0.00905f
C10801 a_21964_21976# a_22636_21976# 0.00544f
C10802 _474_.CLK a_54040_22366# 0.00439f
C10803 a_51196_15271# VPWR 0.32932f
C10804 _373_.A2 uo_out[7] 0.00575f
C10805 a_46180_14180# a_46628_14180# 0.01328f
C10806 a_32604_16839# VPWR 0.29679f
C10807 a_22188_30951# a_22548_31048# 0.0869f
C10808 a_44612_1256# VPWR 0.20348f
C10809 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN a_66228_20452# 0.02061f
C10810 a_67117_30600# vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I 0.00245f
C10811 a_3172_13800# a_3172_12612# 0.05841f
C10812 _334_.A1 _363_.Z 2.1771f
C10813 a_40040_17675# a_40108_16839# 0.03137f
C10814 a_31172_17316# VPWR 0.20348f
C10815 a_16500_23208# a_16500_22020# 0.05841f
C10816 a_53796_1636# VPWR 0.20874f
C10817 a_16700_1159# a_17060_1256# 0.08717f
C10818 a_46716_12135# a_47076_12232# 0.08717f
C10819 a_9892_29480# a_10340_29480# 0.01328f
C10820 a_60716_12135# a_61164_12135# 0.01288f
C10821 a_52092_12568# a_52004_11044# 0.00151f
C10822 a_9756_1592# a_10204_1592# 0.01288f
C10823 a_13700_1636# a_13788_1592# 0.28563f
C10824 a_61948_27815# VPWR 0.32915f
C10825 a_30476_23544# a_30588_23111# 0.02634f
C10826 a_8188_29816# a_8860_29816# 0.00544f
C10827 a_59955_30600# _270_.A2 0.00518f
C10828 a_54468_15368# a_54468_14180# 0.05841f
C10829 a_47076_31048# a_47524_31048# 0.01328f
C10830 a_58500_11044# a_58476_10567# 0.00172f
C10831 a_54556_11000# a_54668_10567# 0.02634f
C10832 a_29916_1592# a_29916_1159# 0.05841f
C10833 _459_.CLK a_19948_26680# 0.02236f
C10834 a_24676_2824# VPWR 0.20815f
C10835 _301_.A1 a_39172_22504# 0.00136f
C10836 a_63764_23208# vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I 0.00438f
C10837 _334_.A1 a_36960_27912# 0.01039f
C10838 _459_.CLK a_15692_27815# 0.00105f
C10839 a_14796_24679# a_14708_24776# 0.28563f
C10840 a_23196_24679# a_23644_24679# 0.01288f
C10841 a_1916_23111# a_1828_23208# 0.28563f
C10842 _438_.A2 _303_.ZN 0.75229f
C10843 a_31260_19975# a_31708_19975# 0.0131f
C10844 a_2724_7528# a_3172_7528# 0.01328f
C10845 a_66652_1159# a_67100_1159# 0.01255f
C10846 _350_.A2 _371_.A2 0.05256f
C10847 a_1828_9096# a_2276_9096# 0.01328f
C10848 _230_.I ui_in[1] 0.04344f
C10849 a_45732_14180# VPWR 0.20812f
C10850 a_3620_5960# a_4068_5960# 0.01328f
C10851 _395_.A1 _218_.ZN 0.19878f
C10852 a_1916_18407# a_2276_18504# 0.08717f
C10853 a_32604_18407# a_33052_18407# 0.0131f
C10854 a_4852_4392# a_5300_4392# 0.01328f
C10855 a_4940_4295# a_4964_3204# 0.0016f
C10856 a_33376_23659# a_35232_24029# 0.02307f
C10857 _313_.ZN a_33932_24073# 0.22517f
C10858 _390_.ZN _398_.C 0.18164f
C10859 _452_.CLK _305_.A2 0.17215f
C10860 vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN VPWR 0.7068f
C10861 a_54356_25156# a_54804_25156# 0.01328f
C10862 _252_.ZN _250_.ZN 0.28962f
C10863 a_39268_18840# a_39264_18147# 0.00551f
C10864 a_60268_12135# VPWR 0.31389f
C10865 a_35740_15704# a_36188_15704# 0.01288f
C10866 _397_.A1 _424_.B1 0.07092f
C10867 a_9444_29480# VPWR 0.20348f
C10868 a_46628_31048# VPWR 0.22451f
C10869 _334_.A1 a_33812_29860# 0.00351f
C10870 a_61297_30300# VPWR 0.49238f
C10871 vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN a_63180_26680# 0.05355f
C10872 _474_.CLK a_54892_26680# 0.00768f
C10873 a_50884_15748# a_50748_15271# 0.00168f
C10874 a_46940_15704# a_46940_15271# 0.05841f
C10875 a_22748_24679# VPWR 0.31592f
C10876 _285_.Z _437_.A1 0.34488f
C10877 a_2276_7528# VPWR 0.20634f
C10878 a_34276_23705# VPWR 0.00267f
C10879 a_4068_4392# VPWR 0.22146f
C10880 _251_.A1 _237_.A1 0.18358f
C10881 a_53908_25156# VPWR 0.2249f
C10882 a_35292_15704# VPWR 0.33596f
C10883 a_41392_27165# a_41099_26841# 0.49319f
C10884 a_51756_18407# a_52204_18407# 0.0131f
C10885 _474_.CLK vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN 0.00412f
C10886 a_58116_30344# a_58340_29860# 0.01342f
C10887 a_28908_21976# a_29356_21976# 0.01288f
C10888 a_66340_15368# a_66340_14180# 0.05841f
C10889 a_40092_27209# VPWR 0.39697f
C10890 a_54892_16839# vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN 0.00597f
C10891 _452_.CLK a_45260_17272# 0.00375f
C10892 a_51308_18407# VPWR 0.32117f
C10893 _324_.C a_44786_24120# 0.00895f
C10894 a_22636_28248# a_23084_28248# 0.01222f
C10895 a_22996_28292# _454_.Q 0.00461f
C10896 a_47297_25596# VPWR 0.48613f
C10897 a_54444_16839# VPWR 0.32732f
C10898 a_67460_1256# a_67908_1256# 0.01328f
C10899 _275_.A2 _474_.CLK 0.0839f
C10900 _337_.A3 a_27228_26247# 0.0016f
C10901 _397_.A1 _386_.ZN 0.03867f
C10902 a_67012_1256# VPWR 0.20348f
C10903 a_46716_2727# a_47164_2727# 0.0131f
C10904 a_43828_29860# vgaringosc.workerclkbuff_notouch_.I 0.05224f
C10905 a_47612_18407# a_47748_17316# 0.00154f
C10906 a_51444_13800# a_51556_12612# 0.02666f
C10907 a_67572_13800# a_68020_13800# 0.01328f
C10908 _325_.A2 a_42996_18840# 0.00914f
C10909 _287_.A1 _370_.B 0.06246f
C10910 _260_.A1 _441_.A3 0.00656f
C10911 _459_.CLK _460_.Q 0.0991f
C10912 a_23556_23208# a_23444_22020# 0.02666f
C10913 _358_.A3 a_33520_25597# 0.00899f
C10914 a_59932_1592# VPWR 0.29679f
C10915 a_28124_1159# a_28036_1256# 0.28563f
C10916 a_58028_12135# a_57940_12232# 0.28563f
C10917 _346_.A2 a_21424_25987# 0.00421f
C10918 a_17060_1636# a_16700_1592# 0.08707f
C10919 _304_.B _412_.ZN 0.05562f
C10920 a_15132_29816# a_15580_29816# 0.01288f
C10921 a_15692_21543# VPWR 0.29679f
C10922 _476_.Q _424_.A1 1.42846f
C10923 vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I 0.0101f
C10924 a_47076_2824# VPWR 0.20815f
C10925 a_65444_11044# a_65420_10567# 0.00172f
C10926 a_47612_10567# a_48060_10567# 0.0131f
C10927 a_60380_1592# a_60828_1592# 0.01288f
C10928 _300_.ZN a_39772_20408# 0.00655f
C10929 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 1.25234f
C10930 a_25436_24679# a_25796_24776# 0.08663f
C10931 a_21852_23111# a_22212_23208# 0.08707f
C10932 a_49988_9476# VPWR 0.21421f
C10933 a_62844_27815# a_62756_27912# 0.28563f
C10934 a_50276_27912# VPWR 0.00477f
C10935 a_22100_31048# VPWR 0.20773f
C10936 a_16140_21543# a_16588_21543# 0.0131f
C10937 a_60180_14180# VPWR 0.20924f
C10938 _324_.B _325_.B 0.30621f
C10939 _313_.ZN a_33708_22505# 0.00429f
C10940 a_60909_30600# _246_.B2 0.00349f
C10941 _294_.A2 a_34532_27208# 0.00138f
C10942 a_1916_29816# a_1916_29383# 0.05841f
C10943 a_5860_29860# a_5724_29383# 0.00168f
C10944 a_54132_12232# VPWR 0.20622f
C10945 a_43044_15748# a_42684_15704# 0.08707f
C10946 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I a_56708_15368# 0.00134f
C10947 a_47524_2824# a_47972_2824# 0.01328f
C10948 uo_out[0] uio_in[7] 0.01021f
C10949 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I clk 0.00389f
C10950 _323_.A3 _448_.D 0.03555f
C10951 _390_.ZN _393_.A3 0.00285f
C10952 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN 0.69544f
C10953 a_50384_19204# a_50796_19001# 0.00275f
C10954 a_26548_24372# VPWR 0.01232f
C10955 a_26556_30951# _340_.A2 0.01477f
C10956 _447_.Q _319_.A3 0.01949f
C10957 _417_.A2 a_49988_21236# 0.02232f
C10958 a_7964_2727# a_7876_2824# 0.28563f
C10959 a_49092_15748# VPWR 0.20929f
C10960 _412_.A1 a_49764_26724# 0.42641f
C10961 a_48508_9432# a_49180_9432# 0.00544f
C10962 a_50436_9476# a_50884_9476# 0.01328f
C10963 _442_.ZN a_39236_26344# 0.00675f
C10964 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I a_59260_21976# 0.00529f
C10965 a_59172_22020# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I 0.01673f
C10966 a_53212_14136# a_53660_14136# 0.0131f
C10967 a_56708_14180# a_56796_14136# 0.28563f
C10968 a_22548_31048# a_22996_31048# 0.01328f
C10969 _452_.CLK a_36996_26344# 0.00546f
C10970 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN 0.07373f
C10971 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_62756_27912# 0.01178f
C10972 _437_.A1 a_37444_26724# 0.00228f
C10973 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN a_57828_25156# 0.04011f
C10974 _334_.A1 uo_out[3] 0.0047f
C10975 a_10652_1592# a_10788_1256# 0.00168f
C10976 vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN a_54780_18840# 0.01934f
C10977 a_54580_13800# a_54556_12568# 0.0016f
C10978 a_58388_13800# a_58500_12612# 0.02666f
C10979 a_56484_23208# vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.002f
C10980 _304_.B _452_.Q 0.12913f
C10981 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN 0.63083f
C10982 a_34308_26344# VPWR 0.67167f
C10983 _355_.C a_21740_29383# 0.00621f
C10984 a_30500_23208# a_30388_22020# 0.02666f
C10985 a_1828_24776# a_1828_23588# 0.05841f
C10986 a_4852_7528# a_4964_6340# 0.02666f
C10987 a_52428_12135# a_52452_11044# 0.0016f
C10988 a_9980_1159# VPWR 0.33193f
C10989 a_39100_1159# a_39460_1256# 0.08717f
C10990 a_54580_12232# a_55028_12232# 0.01328f
C10991 a_23420_1592# a_23868_1592# 0.012f
C10992 _412_.ZN VPWR 0.30801f
C10993 a_3620_21640# VPWR 0.22347f
C10994 _334_.A1 a_35660_27508# 0.06942f
C10995 _437_.A1 a_37408_23208# 0.00108f
C10996 a_50884_17316# a_50524_17272# 0.08707f
C10997 a_62308_27912# VPWR 0.20622f
C10998 _340_.A2 a_28054_30196# 0.01469f
C10999 a_5388_10567# a_5300_10664# 0.28563f
C11000 _395_.A1 _407_.A1 0.00486f
C11001 _370_.B a_28000_29480# 0.01033f
C11002 _459_.Q uo_out[6] 0.00831f
C11003 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN a_57580_13703# 0.00144f
C11004 a_32828_23111# a_32740_23208# 0.28563f
C11005 a_62508_23111# VPWR 0.32937f
C11006 _337_.A3 _336_.A2 1.33637f
C11007 a_1468_23544# VPWR 0.29679f
C11008 _316_.ZN a_33708_22505# 0.23272f
C11009 a_33152_22091# a_35008_22461# 0.02307f
C11010 a_60964_9476# VPWR 0.20595f
C11011 a_67772_14136# VPWR 0.33516f
C11012 a_3260_3160# VPWR 0.30487f
C11013 a_14796_21543# a_15156_21640# 0.08717f
C11014 _427_.A2 a_51540_23588# 0.01325f
C11015 a_1468_6296# VPWR 0.29679f
C11016 a_54356_26724# a_53996_26680# 0.0869f
C11017 _267_.A2 _258_.I 1.30848f
C11018 a_43296_28733# a_43940_27912# 0.00172f
C11019 _474_.CLK a_55700_25156# 0.02564f
C11020 a_16164_31048# a_16028_29816# 0.00154f
C11021 _424_.A2 a_45920_20523# 0.02404f
C11022 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN 0.7984f
C11023 _285_.Z a_37844_29860# 0.00166f
C11024 a_35652_25156# VPWR 0.17189f
C11025 a_49540_15748# a_49988_15748# 0.01328f
C11026 a_3708_11000# VPWR 0.33374f
C11027 _346_.A2 _351_.ZN 0.00447f
C11028 a_65308_19975# a_66004_20072# 0.01227f
C11029 _402_.B _324_.B 0.08089f
C11030 _251_.A1 _242_.Z 0.04712f
C11031 _397_.A2 _470_.Q 1.0899f
C11032 _474_.CLK a_53100_18407# 0.00721f
C11033 _331_.ZN a_41572_18504# 0.00759f
C11034 a_34308_18884# VPWR 0.21975f
C11035 _304_.A1 a_33636_23208# 0.00395f
C11036 a_50276_27912# a_50068_27508# 0.01565f
C11037 _359_.B a_36500_29860# 0.00553f
C11038 a_4156_26247# VPWR 0.3269f
C11039 a_18940_2727# a_19300_2824# 0.08717f
C11040 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_64972_26680# 0.03562f
C11041 _432_.ZN _226_.ZN 0.00982f
C11042 a_35652_31048# uo_out[3] 0.00345f
C11043 _454_.Q _371_.A2 1.32562f
C11044 a_1020_9432# a_1020_8999# 0.05841f
C11045 a_56036_9476# a_56124_9432# 0.28563f
C11046 _334_.A1 a_37291_29535# 0.02108f
C11047 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I a_65668_27912# 0.00205f
C11048 _370_.ZN a_29575_28293# 0.07669f
C11049 a_27116_21976# a_27028_20452# 0.00151f
C11050 _460_.Q uo_out[7] 0.04552f
C11051 a_4604_20408# a_5052_20408# 0.01222f
C11052 a_53660_17272# a_53572_15748# 0.00151f
C11053 _461_.D uo_out[6] 0.01868f
C11054 a_61412_14180# a_61500_14136# 0.28563f
C11055 a_50748_14136# a_50636_13703# 0.02634f
C11056 a_24392_28248# a_25124_28776# 0.02695f
C11057 a_48956_12568# a_49404_12568# 0.01288f
C11058 a_65332_13800# a_65444_12612# 0.02666f
C11059 _438_.ZN a_39475_21236# 0.00201f
C11060 _452_.Q VPWR 3.28463f
C11061 a_19524_24776# a_19636_23588# 0.02666f
C11062 a_32380_1159# VPWR 0.29679f
C11063 _432_.ZN _300_.ZN 0.0935f
C11064 _433_.ZN _325_.A1 0.67597f
C11065 _474_.CLK a_54556_21543# 0.00855f
C11066 a_50524_1159# a_50436_1256# 0.28563f
C11067 a_30724_1636# a_30364_1592# 0.08707f
C11068 a_59372_12135# a_59396_11044# 0.0016f
C11069 _359_.B _462_.D 0.96164f
C11070 a_39324_26247# _431_.A3 0.01333f
C11071 _330_.A1 _260_.A1 0.00197f
C11072 a_35044_21640# VPWR 0.0251f
C11073 a_35204_26344# a_35652_26344# 0.01328f
C11074 _302_.Z a_42168_22504# 1.37932f
C11075 _452_.Q a_41012_23208# 0.00595f
C11076 a_1828_10664# a_2276_10664# 0.01328f
C11077 a_55564_10567# a_55924_10664# 0.08707f
C11078 a_10428_1159# a_10876_1159# 0.0131f
C11079 _355_.C a_24228_26344# 0.01738f
C11080 a_48964_20204# VPWR 0.00964f
C11081 _260_.A2 _441_.A3 0.12864f
C11082 a_2364_21976# VPWR 0.30029f
C11083 a_54332_18840# a_54356_18504# 0.00172f
C11084 a_31396_23208# a_31844_23208# 0.01328f
C11085 a_35616_24776# a_36172_24463# 0.8399f
C11086 _402_.A1 a_42148_27912# 0.00468f
C11087 a_24340_23588# VPWR 0.20631f
C11088 a_67100_8999# VPWR 0.29679f
C11089 a_40356_2824# a_40444_1159# 0.0027f
C11090 a_4068_21640# a_4852_21640# 0.00276f
C11091 a_25884_21543# a_25796_21640# 0.28563f
C11092 _467_.D a_15156_28292# 0.00187f
C11093 _383_.A2 a_47525_29480# 0.00403f
C11094 _397_.A1 _386_.A4 1.02296f
C11095 a_62060_13703# VPWR 0.31556f
C11096 a_1380_18884# a_1468_18840# 0.28563f
C11097 a_12444_2727# VPWR 0.31605f
C11098 _260_.ZN _328_.A2 0.00164f
C11099 _324_.C _395_.A3 0.02316f
C11100 a_67117_30600# VPWR 0.5739f
C11101 _304_.B a_53908_26724# 0.00497f
C11102 a_36960_27912# a_37532_26680# 0.00105f
C11103 _443_.D a_37084_26680# 0.00194f
C11104 a_57156_11044# VPWR 0.21061f
C11105 _459_.CLK a_17148_29383# 0.04961f
C11106 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN a_54692_26344# 0.005f
C11107 a_27004_27815# a_27140_26724# 0.00154f
C11108 a_19860_26724# VPWR 0.16504f
C11109 _461_.D uo_out[5] 0.00133f
C11110 _373_.A2 _340_.A2 0.11653f
C11111 _462_.D a_36656_29123# 0.00472f
C11112 _474_.Q a_47552_19715# 0.00472f
C11113 a_67012_15748# a_67460_15748# 0.01328f
C11114 a_64324_15748# a_63964_15704# 0.08717f
C11115 a_1916_27815# VPWR 0.297f
C11116 a_62956_23111# a_63404_23111# 0.0131f
C11117 a_30364_2727# a_30276_2824# 0.28563f
C11118 a_41264_30669# uo_out[3] 0.00117f
C11119 _388_.B a_41708_30644# 0.02944f
C11120 a_47636_18884# a_47724_18840# 0.28563f
C11121 _416_.A1 a_44961_27912# 0.01392f
C11122 _268_.A2 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I 0.04381f
C11123 _252_.B vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN 0.0147f
C11124 _378_.ZN VPWR 0.47224f
C11125 a_61412_9476# a_61860_9476# 0.01328f
C11126 a_1916_23544# a_2364_23544# 0.0131f
C11127 a_4516_23588# a_4156_23544# 0.08674f
C11128 a_11236_1256# a_11684_1256# 0.01328f
C11129 a_4516_6340# a_4156_6296# 0.08674f
C11130 a_1020_7864# a_1468_7864# 0.0131f
C11131 a_3620_7908# a_3260_7864# 0.08717f
C11132 a_1916_6296# a_2364_6296# 0.0131f
C11133 a_17284_31048# a_17732_31048# 0.01328f
C11134 a_2812_4728# a_3260_4728# 0.0131f
C11135 a_1020_13703# a_1468_13703# 0.0131f
C11136 a_3708_3160# a_4156_3160# 0.0131f
C11137 a_19412_20452# a_19500_20408# 0.28563f
C11138 _230_.I _324_.C 0.12478f
C11139 a_1916_29383# a_2364_29383# 0.0131f
C11140 a_2812_30951# a_2724_31048# 0.28563f
C11141 a_5948_1592# VPWR 0.3289f
C11142 a_2812_12568# a_2812_12135# 0.05841f
C11143 _459_.Q a_33612_24679# 0.00334f
C11144 a_56260_12612# a_55900_12568# 0.08707f
C11145 _459_.CLK a_16588_25112# 0.00189f
C11146 a_58836_13800# a_58924_12135# 0.00151f
C11147 _433_.ZN _327_.A2 0.10165f
C11148 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_61164_23111# 0.05629f
C11149 _355_.ZN a_28348_23111# 0.00279f
C11150 a_61276_1159# a_61860_1256# 0.01675f
C11151 a_45696_20072# a_46624_19715# 1.16391f
C11152 a_54780_1159# VPWR 0.29679f
C11153 a_66316_12135# a_66340_11044# 0.0016f
C11154 a_63516_18840# VPWR 0.29679f
C11155 a_56372_12232# a_56260_11044# 0.02666f
C11156 a_1828_16936# a_2276_16936# 0.01328f
C11157 a_33636_1636# a_33724_1592# 0.28563f
C11158 a_37220_1636# a_37668_1636# 0.01328f
C11159 a_4156_11000# a_4604_11000# 0.01222f
C11160 a_36100_25156# a_36548_25156# 0.01328f
C11161 _346_.A2 a_21044_27508# 0.51116f
C11162 a_43132_27815# _330_.A1 0.00502f
C11163 a_44028_27815# a_43940_27912# 0.28563f
C11164 a_52512_19715# _424_.ZN 0.24727f
C11165 _311_.A2 _430_.ZN 0.15141f
C11166 _467_.D a_16052_27912# 0.00857f
C11167 a_66764_10567# a_66676_10664# 0.28563f
C11168 a_32068_18504# a_32068_17316# 0.05841f
C11169 a_62084_1636# a_61948_1159# 0.00168f
C11170 a_58140_1592# a_58140_1159# 0.05841f
C11171 _384_.ZN a_49405_22805# 0.0024f
C11172 a_25236_22020# VPWR 0.20614f
C11173 _223_.I a_29232_29931# 0.00113f
C11174 _355_.C a_22548_29480# 0.00646f
C11175 _350_.A2 _294_.ZN 0.05041f
C11176 _260_.A1 _226_.ZN 1.23708f
C11177 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN a_57580_23544# 0.00717f
C11178 _416_.A1 _480_.Q 0.03126f
C11179 a_32964_18884# a_33052_18840# 0.28563f
C11180 a_34620_2727# VPWR 0.35448f
C11181 a_30812_18840# a_31260_18840# 0.0131f
C11182 a_4940_26247# a_5388_26247# 0.01222f
C11183 a_55924_13800# VPWR 0.20622f
C11184 _379_.A2 a_18400_28733# 0.00632f
C11185 a_11460_29860# VPWR 0.22977f
C11186 a_53908_26724# VPWR 0.23143f
C11187 a_55340_25112# a_55788_25112# 0.012f
C11188 a_63740_11000# VPWR 0.31389f
C11189 _350_.A2 a_29351_28293# 0.00115f
C11190 _470_.Q _330_.A1 0.52378f
C11191 a_62644_16936# a_62532_15748# 0.02666f
C11192 a_2364_15271# a_2724_15368# 0.08717f
C11193 a_22300_23111# VPWR 0.33016f
C11194 _386_.ZN _389_.ZN 0.04774f
C11195 _335_.ZN _443_.D 0.00119f
C11196 a_20379_29977# a_20664_29977# 0.00277f
C11197 _459_.CLK a_26427_29977# 0.00275f
C11198 _304_.B _436_.B 0.26929f
C11199 _474_.CLK vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN 0.00172f
C11200 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _274_.ZN 0.07855f
C11201 a_41340_2727# a_41700_2824# 0.08717f
C11202 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I 0.01777f
C11203 _261_.ZN _325_.A1 0.31082f
C11204 _260_.A1 _300_.ZN 0.16746f
C11205 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN 0.04782f
C11206 _242_.Z a_58020_27508# 0.46923f
C11207 a_28000_29480# a_28556_29167# 0.8399f
C11208 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN 0.01427f
C11209 _416_.A1 uio_in[0] 0.03094f
C11210 a_63628_16839# a_63540_16936# 0.28563f
C11211 a_67012_9476# a_67100_9432# 0.28563f
C11212 a_61724_18407# a_62172_18407# 0.0131f
C11213 a_18292_23588# a_17932_23544# 0.08707f
C11214 a_3172_25156# a_2812_25112# 0.08717f
C11215 a_66452_20072# a_66564_18884# 0.02666f
C11216 a_55004_14136# a_55028_13800# 0.00172f
C11217 a_24652_20408# a_25100_20408# 0.0131f
C11218 _267_.A2 _255_.ZN 0.0352f
C11219 a_17372_30951# a_17732_31048# 0.0869f
C11220 uio_out[3] uio_out[4] 0.06758f
C11221 _324_.C a_44038_21236# 0.0012f
C11222 a_67100_17272# a_66988_16839# 0.02634f
C11223 a_57692_11000# a_57604_9476# 0.00151f
C11224 a_62756_12612# a_63204_12612# 0.01328f
C11225 a_19748_1636# VPWR 0.2159f
C11226 a_61297_30300# a_61689_29860# 0.00762f
C11227 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN a_64324_29860# 0.01046f
C11228 a_60852_15748# a_61300_15748# 0.01328f
C11229 a_17148_29816# _467_.D 0.00312f
C11230 a_33612_24679# _313_.ZN 0.00193f
C11231 a_61412_17316# a_61500_17272# 0.28563f
C11232 a_62172_15271# a_62532_15368# 0.08717f
C11233 a_63316_12232# a_63204_11044# 0.02666f
C11234 a_8772_1636# a_8636_1159# 0.00168f
C11235 a_31620_18504# VPWR 0.20348f
C11236 a_51108_11044# a_50748_11000# 0.08707f
C11237 a_56260_31048# _274_.A2 0.00397f
C11238 _336_.A2 a_27328_25227# 0.04941f
C11239 hold1.Z a_43126_24119# 0.03894f
C11240 _312_.ZN _301_.A1 0.0011f
C11241 _427_.ZN VPWR 0.54384f
C11242 a_63316_10664# a_63764_10664# 0.01328f
C11243 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN _267_.A1 0.0421f
C11244 _419_.A4 _381_.A2 0.03785f
C11245 a_32828_1159# a_33276_1159# 0.0131f
C11246 a_40357_24776# VPWR 0.51924f
C11247 a_29828_2824# a_29828_1636# 0.05841f
C11248 a_26020_2824# a_25884_1592# 0.00154f
C11249 a_67436_18407# a_67460_17316# 0.0016f
C11250 _448_.Q _438_.ZN 0.21091f
C11251 a_25348_24776# a_25436_23111# 0.00151f
C11252 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I a_60852_15748# 0.00193f
C11253 _355_.C a_26556_28776# 0.00163f
C11254 _365_.ZN _452_.CLK 0.01761f
C11255 a_62756_2824# a_62844_1159# 0.0027f
C11256 a_45284_12612# VPWR 0.22176f
C11257 a_57020_2727# VPWR 0.31581f
C11258 a_64412_18407# a_64772_18504# 0.08717f
C11259 a_36772_15368# a_37220_15368# 0.01328f
C11260 a_932_20072# VPWR 0.22176f
C11261 a_61836_23544# a_62284_23544# 0.01222f
C11262 a_58028_10567# VPWR 0.33765f
C11263 a_38876_15271# a_38788_15368# 0.28563f
C11264 _459_.CLK a_29184_25597# 0.0365f
C11265 a_19972_23208# VPWR 0.20631f
C11266 a_58700_16839# vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I 0.00573f
C11267 _251_.A1 vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN 0.00578f
C11268 _436_.B VPWR 1.17897f
C11269 a_40220_15271# a_40668_15271# 0.0131f
C11270 _427_.ZN a_54108_21543# 0.01268f
C11271 _330_.A1 a_36084_23208# 0.00141f
C11272 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.00102f
C11273 a_4516_28292# a_4604_28248# 0.28563f
C11274 _324_.C _325_.A2 0.04971f
C11275 a_40220_20408# _325_.A2 0.00231f
C11276 a_2812_21976# a_3260_21976# 0.0131f
C11277 a_52764_2727# a_52676_2824# 0.28563f
C11278 a_64412_17272# a_64860_17272# 0.0131f
C11279 a_30724_26020# VPWR 0.77617f
C11280 a_18628_23208# a_18716_21543# 0.00151f
C11281 a_33636_1256# a_34084_1256# 0.01328f
C11282 a_16948_25156# a_16588_25112# 0.08707f
C11283 a_4940_19975# a_4964_18884# 0.0016f
C11284 a_24788_23588# a_25236_23588# 0.01328f
C11285 a_3260_18840# a_3260_18407# 0.05841f
C11286 a_12892_2727# a_13340_2727# 0.0131f
C11287 a_62508_13703# a_62956_13703# 0.01288f
C11288 a_48508_13703# a_49204_13800# 0.01227f
C11289 a_30388_20452# a_30476_20408# 0.28563f
C11290 VPWR uio_out[6] 1.23078f
C11291 a_37532_26247# _444_.D 0.00453f
C11292 a_35628_16839# a_35988_16936# 0.08707f
C11293 _317_.A2 a_34716_20937# 0.00141f
C11294 a_50644_21640# a_49988_21236# 0.01565f
C11295 a_52876_10567# a_52900_9476# 0.0016f
C11296 a_25884_1592# VPWR 0.33312f
C11297 a_60292_12612# a_60268_12135# 0.00172f
C11298 a_56348_12568# a_56460_12135# 0.02634f
C11299 _352_.A2 a_28596_26725# 0.13115f
C11300 _350_.A1 _285_.Z 0.05001f
C11301 a_17372_30951# a_17820_30951# 0.01255f
C11302 a_1916_25112# a_1916_24679# 0.05841f
C11303 a_67348_18504# a_67796_18504# 0.01328f
C11304 a_57604_11044# a_58052_11044# 0.01328f
C11305 a_54020_11044# a_54108_11000# 0.28563f
C11306 a_48756_16936# a_49204_16936# 0.01328f
C11307 _330_.A1 a_37892_17316# 0.0044f
C11308 a_47300_1636# a_47388_1592# 0.28563f
C11309 a_43356_1592# a_43804_1592# 0.01288f
C11310 a_15580_1592# a_15580_1159# 0.05841f
C11311 _324_.B a_46352_22021# 0.02687f
C11312 _395_.A3 _281_.A1 1.10134f
C11313 _474_.CLK a_49740_29383# 0.00696f
C11314 _352_.A2 _358_.A3 0.00576f
C11315 _371_.A1 _355_.B 0.01678f
C11316 a_17803_26841# a_17168_27165# 0.02112f
C11317 a_18096_27165# a_16240_26795# 0.02366f
C11318 a_20308_26724# a_20756_26724# 0.01328f
C11319 _231_.I VPWR 0.80044f
C11320 _435_.ZN _304_.A1 0.00307f
C11321 _246_.B2 a_59260_26680# 0.04903f
C11322 a_4604_9432# a_4516_7908# 0.0027f
C11323 _230_.I _252_.ZN 0.03793f
C11324 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I 0.65551f
C11325 a_56484_29480# vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I 0.00445f
C11326 a_48084_18884# VPWR 0.20771f
C11327 _346_.B _346_.ZN 0.01765f
C11328 _455_.D a_21424_25987# 0.0069f
C11329 a_20308_20452# VPWR 0.20677f
C11330 a_2364_27815# a_2812_27815# 0.0131f
C11331 _474_.CLK a_48141_29480# 0.0015f
C11332 a_50084_24328# _399_.ZN 0.00172f
C11333 a_37968_31048# VPWR 0.01424f
C11334 _304_.B _268_.A1 0.09942f
C11335 _334_.A1 _294_.ZN 0.24277f
C11336 a_58948_12612# VPWR 0.20703f
C11337 a_13700_2824# a_14148_2824# 0.01328f
C11338 a_11324_29383# a_11684_29480# 0.08717f
C11339 _397_.Z _399_.A2 0.77658f
C11340 a_38584_28292# a_39256_28292# 0.00488f
C11341 a_36548_15748# a_36412_15271# 0.00168f
C11342 a_32604_15704# a_32604_15271# 0.05841f
C11343 a_51892_10664# VPWR 0.20641f
C11344 _474_.Q a_49764_23588# 0.00155f
C11345 a_52316_27815# a_52228_27912# 0.28563f
C11346 a_49852_15271# a_50212_15368# 0.08717f
C11347 _370_.ZN _371_.A2 0.00504f
C11348 a_1380_21640# a_1380_20452# 0.05841f
C11349 a_2812_4295# a_2724_4392# 0.28563f
C11350 a_1916_5863# a_1828_5960# 0.28563f
C11351 a_36636_26680# a_37084_26680# 0.01255f
C11352 _251_.A1 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I 0.07801f
C11353 _260_.A2 _226_.ZN 0.00444f
C11354 _389_.ZN a_47476_28292# 0.0063f
C11355 a_67324_15271# VPWR 0.32932f
C11356 _441_.B a_39780_22805# 0.00359f
C11357 _475_.D a_46476_20937# 0.22486f
C11358 a_63740_2727# a_64100_2824# 0.08717f
C11359 _256_.A2 _258_.I 0.00219f
C11360 a_54444_25112# clk 0.00335f
C11361 a_19188_22020# a_18828_21976# 0.08707f
C11362 _421_.A1 _421_.B 0.45397f
C11363 a_3260_15271# VPWR 0.30487f
C11364 a_48060_30951# a_48420_31048# 0.08717f
C11365 a_67236_15368# a_67684_15368# 0.01328f
C11366 _459_.Q _460_.Q 2.03964f
C11367 a_26970_29480# VPWR 0.01637f
C11368 _274_.A2 a_57500_30344# 0.00136f
C11369 a_65756_7864# VPWR 0.31505f
C11370 a_21764_1256# VPWR 0.20348f
C11371 a_28820_24072# a_29028_24072# 0.00334f
C11372 a_22636_25112# a_23084_25112# 0.01222f
C11373 _397_.A1 a_46794_25156# 0.00124f
C11374 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I 0.04475f
C11375 _249_.A2 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I 0.02533f
C11376 a_67548_4728# VPWR 0.29679f
C11377 a_59820_13703# a_59732_13800# 0.28563f
C11378 a_12444_29383# VPWR 0.30141f
C11379 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN a_56260_15368# 0.0015f
C11380 a_3708_30951# VPWR 0.34839f
C11381 a_46604_16839# a_46516_16936# 0.28563f
C11382 _470_.D a_43008_26795# 0.27272f
C11383 a_43232_29480# a_44160_29123# 1.16391f
C11384 _474_.CLK a_49600_30180# 0.02246f
C11385 a_37332_16936# VPWR 0.2061f
C11386 a_39548_1592# VPWR 0.32517f
C11387 a_5276_1159# a_5636_1256# 0.08717f
C11388 _260_.A2 _300_.ZN 0.00118f
C11389 a_67236_12612# a_67212_12135# 0.00172f
C11390 a_54444_24679# VPWR 0.29679f
C11391 a_6396_1592# a_6844_1592# 0.01288f
C11392 _388_.B uo_out[0] 0.00772f
C11393 a_49740_12135# a_50188_12135# 0.01288f
C11394 a_21876_25156# a_21852_24679# 0.00172f
C11395 a_17932_25112# a_17932_24679# 0.05841f
C11396 _386_.A4 _389_.ZN 0.31711f
C11397 a_5412_29860# a_5052_29816# 0.08707f
C11398 a_33708_22505# a_33724_21543# 0.0019f
C11399 _447_.Q _305_.A2 0.52099f
C11400 a_67572_12232# a_67660_10567# 0.00151f
C11401 a_48508_30951# VPWR 0.31143f
C11402 a_50660_1636# a_50300_1592# 0.08707f
C11403 a_1828_2824# VPWR 0.20348f
C11404 _384_.A3 a_50420_23233# 0.00133f
C11405 _459_.CLK _346_.B 0.01421f
C11406 a_48732_15271# a_48868_14180# 0.00154f
C11407 _424_.ZN a_53348_18884# 0.00456f
C11408 _243_.ZN a_59172_27912# 0.10906f
C11409 _459_.CLK a_17484_26247# 0.0081f
C11410 a_2812_24679# a_3260_24679# 0.0131f
C11411 a_42896_18504# a_43776_18191# 0.00306f
C11412 a_55228_1159# a_55676_1159# 0.0131f
C11413 a_50412_18407# a_50324_18504# 0.28563f
C11414 _448_.Q a_37744_20452# 0.00373f
C11415 a_41776_20072# _450_.D 0.00621f
C11416 _325_.A1 _327_.Z 0.00349f
C11417 a_47972_18504# VPWR 0.20897f
C11418 a_63964_18840# a_64412_18840# 0.0131f
C11419 _352_.A2 a_25884_24679# 0.01249f
C11420 a_19636_25156# VPWR 0.21729f
C11421 a_17484_27815# a_17396_27912# 0.28563f
C11422 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN 0.03998f
C11423 _452_.Q _260_.ZN 0.08381f
C11424 a_20250_31048# VPWR 0.01454f
C11425 a_31284_20452# VPWR 0.20595f
C11426 _268_.A1 VPWR 1.25532f
C11427 a_65532_12568# VPWR 0.32412f
C11428 a_32516_15748# a_32964_15748# 0.01328f
C11429 a_34160_20523# a_35040_20937# 0.00306f
C11430 _381_.Z a_49764_26724# 0.05981f
C11431 _395_.A2 a_50120_26476# 0.00968f
C11432 _324_.C a_43940_27912# 0.01173f
C11433 a_35000_22137# VPWR 0.0037f
C11434 _337_.ZN VPWR 1.63829f
C11435 _393_.ZN _397_.A2 0.01596f
C11436 a_67796_16936# VPWR 0.21165f
C11437 a_47300_15368# VPWR 0.20952f
C11438 _474_.CLK a_48376_27508# 0.00513f
C11439 _352_.A2 a_28256_25597# 0.05026f
C11440 a_25684_22020# a_26132_22020# 0.01328f
C11441 a_28672_31048# uo_out[7] 0.00109f
C11442 a_50748_15271# VPWR 0.33868f
C11443 a_43916_16839# a_44364_16839# 0.01288f
C11444 a_32156_16839# VPWR 0.29679f
C11445 a_56036_1256# a_56484_1256# 0.01328f
C11446 a_44164_1256# VPWR 0.20348f
C11447 a_22188_30951# a_22100_31048# 0.28563f
C11448 a_35292_2727# a_35740_2727# 0.0131f
C11449 _441_.ZN _304_.A1 0.03804f
C11450 a_56372_13800# a_57044_13800# 0.00347f
C11451 a_39324_17272# a_39212_16839# 0.02634f
C11452 _355_.C _459_.D 0.54889f
C11453 a_30724_17316# VPWR 0.22176f
C11454 a_58836_10664# a_58948_9476# 0.02666f
C11455 a_53348_1636# VPWR 0.2085f
C11456 a_16700_1159# a_16612_1256# 0.28563f
C11457 a_46716_12135# a_46628_12232# 0.28563f
C11458 a_13700_1636# a_13340_1592# 0.08707f
C11459 a_61500_27815# VPWR 0.33095f
C11460 a_58911_30644# _270_.A2 0.26477f
C11461 a_66452_20072# a_66540_18407# 0.00151f
C11462 a_54356_26724# a_54804_26724# 0.01328f
C11463 a_11908_29860# a_12356_29860# 0.01328f
C11464 a_34396_17272# a_34844_17272# 0.01288f
C11465 a_64188_11000# a_64636_11000# 0.01288f
C11466 a_47836_17272# a_47860_16936# 0.00172f
C11467 a_24228_2824# VPWR 0.20812f
C11468 a_57156_1636# a_57604_1636# 0.01328f
C11469 a_63316_23208# vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I 0.0404f
C11470 _301_.A1 a_38968_22504# 0.00243f
C11471 _448_.Q a_43192_22504# 0.00106f
C11472 a_22748_23111# a_23196_23111# 0.01288f
C11473 a_1468_23111# a_1828_23208# 0.08717f
C11474 _327_.A2 _327_.Z 0.13472f
C11475 _350_.A1 _371_.A1 0.09656f
C11476 _343_.A2 a_24952_29032# 0.22375f
C11477 a_6532_2824# a_6620_1159# 0.0027f
C11478 a_45284_14180# VPWR 0.22176f
C11479 _281_.ZN a_51332_24372# 0.00297f
C11480 a_1916_18407# a_1828_18504# 0.28563f
C11481 _313_.ZN a_34304_24029# 0.01194f
C11482 a_33376_23659# a_33932_24073# 0.8399f
C11483 a_60276_29032# _250_.ZN 0.47448f
C11484 _247_.ZN _238_.I 0.07197f
C11485 _384_.ZN _397_.A4 0.02463f
C11486 a_59820_12135# VPWR 0.31389f
C11487 a_8996_29480# VPWR 0.20348f
C11488 _330_.A2 a_38336_18147# 0.0044f
C11489 a_36100_2824# a_36548_2824# 0.01328f
C11490 _431_.A3 a_39781_24372# 0.00449f
C11491 a_45956_31048# VPWR 0.21215f
C11492 _474_.CLK a_54444_26680# 0.02252f
C11493 a_59620_27208# a_60276_26724# 0.01565f
C11494 a_22300_24679# VPWR 0.33026f
C11495 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_61524_23208# 0.00284f
C11496 a_1828_7528# VPWR 0.20348f
C11497 a_3620_4392# VPWR 0.22347f
C11498 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN 0.00159f
C11499 a_45260_16839# a_45284_15748# 0.0016f
C11500 _330_.A1 _311_.A2 2.13901f
C11501 a_34844_15704# VPWR 0.37398f
C11502 _400_.ZN _284_.A2 0.02853f
C11503 a_3260_9432# a_3708_9432# 0.0131f
C11504 _435_.A3 _284_.B 0.01673f
C11505 _330_.A1 a_37067_19001# 0.01042f
C11506 _474_.CLK a_56236_24679# 0.00799f
C11507 a_62532_15368# a_62396_14136# 0.00154f
C11508 a_48956_14136# a_49404_14136# 0.01288f
C11509 a_50860_18407# VPWR 0.32097f
C11510 a_40464_27165# VPWR 0.18808f
C11511 a_22996_28292# a_23084_28248# 0.28563f
C11512 _452_.CLK a_44812_17272# 0.00613f
C11513 _245_.I1 a_62196_23588# 0.00142f
C11514 _264_.B _432_.ZN 0.01382f
C11515 a_53996_16839# VPWR 0.33016f
C11516 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I 0.74042f
C11517 a_66564_1256# VPWR 0.20631f
C11518 _421_.A1 a_47524_22021# 0.03076f
C11519 _452_.CLK _325_.A1 0.14277f
C11520 _325_.A2 a_38852_18884# 0.00215f
C11521 _304_.B a_41564_26247# 0.05037f
C11522 a_27676_1159# a_28036_1256# 0.08717f
C11523 _358_.A3 a_32592_25227# 0.02476f
C11524 a_66228_10664# a_66116_9476# 0.02666f
C11525 a_59484_1592# VPWR 0.29679f
C11526 a_3620_12232# a_4068_12232# 0.01328f
C11527 a_57580_12135# a_57940_12232# 0.08707f
C11528 a_16612_1636# a_16700_1592# 0.28563f
C11529 a_20196_1636# a_20644_1636# 0.01328f
C11530 _346_.A2 a_20496_26344# 0.00715f
C11531 a_55004_12568# a_54916_11044# 0.00151f
C11532 a_15244_21543# VPWR 0.29679f
C11533 a_61500_11000# a_61612_10567# 0.02634f
C11534 _474_.CLK _272_.B1 0.40317f
C11535 a_46628_2824# VPWR 0.22891f
C11536 a_62868_23208# vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN 0.00137f
C11537 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_56516_26344# 0.07359f
C11538 a_54780_26247# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.0367f
C11539 a_55956_25940# vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I 0.01773f
C11540 a_21852_23111# a_21764_23208# 0.28563f
C11541 _245_.I1 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN 0.00998f
C11542 a_16500_24776# a_16948_24776# 0.01328f
C11543 a_25436_24679# a_25348_24776# 0.28563f
C11544 a_49540_9476# VPWR 0.21186f
C11545 a_21652_31048# VPWR 0.20348f
C11546 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I 0.03855f
C11547 a_62396_27815# a_62756_27912# 0.08663f
C11548 a_59732_14180# VPWR 0.20821f
C11549 a_58052_2824# a_58052_1636# 0.05841f
C11550 _313_.ZN a_34080_22461# 0.00368f
C11551 a_32068_18504# a_32516_18504# 0.01328f
C11552 a_21044_27508# _455_.D 0.00828f
C11553 _294_.A2 a_34348_27208# 0.00105f
C11554 a_38652_15704# a_39100_15704# 0.01288f
C11555 a_53684_12232# VPWR 0.20622f
C11556 a_42596_15748# a_42684_15704# 0.28563f
C11557 _397_.A1 _424_.A2 0.0972f
C11558 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I a_56260_15368# 0.00277f
C11559 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN a_58924_18840# 0.00133f
C11560 a_27924_24776# VPWR 0.16935f
C11561 a_26108_30951# _340_.A2 0.01795f
C11562 _304_.B _474_.CLK 0.44396f
C11563 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN 0.02161f
C11564 a_52204_16839# a_52228_15748# 0.0016f
C11565 a_7516_2727# a_7876_2824# 0.08717f
C11566 _447_.Q a_37532_21543# 0.04158f
C11567 a_31844_21640# a_31820_20408# 0.0016f
C11568 a_48644_15748# VPWR 0.2068f
C11569 _437_.A1 _434_.ZN 0.04419f
C11570 a_34732_19975# a_34644_20072# 0.28563f
C11571 a_30795_29977# VPWR 0.37382f
C11572 _237_.A1 _255_.I 0.40618f
C11573 _274_.ZN _416_.A1 0.06191f
C11574 a_59172_22020# a_59260_21976# 0.28563f
C11575 input9.Z ui_in[4] 0.00133f
C11576 a_56708_14180# a_56348_14136# 0.08674f
C11577 a_3708_14136# a_3708_13703# 0.05841f
C11578 _452_.CLK a_36548_26344# 0.00656f
C11579 a_57468_2727# a_58140_2727# 0.00544f
C11580 _452_.CLK _327_.A2 0.52555f
C11581 _417_.Z a_49492_18840# 0.00248f
C11582 a_45732_12612# a_46180_12612# 0.01328f
C11583 a_54892_18407# vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN 0.00203f
C11584 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN a_53660_17272# 0.00869f
C11585 _304_.A1 _437_.ZN 0.03054f
C11586 _427_.B1 _281_.A1 0.0237f
C11587 a_41564_26247# VPWR 0.35218f
C11588 a_3620_9096# a_3620_7908# 0.05841f
C11589 a_9532_1159# VPWR 0.3289f
C11590 a_39100_1159# a_39012_1256# 0.28563f
C11591 a_1380_20072# a_1828_20072# 0.01328f
C11592 a_932_12232# a_932_11044# 0.05841f
C11593 a_31484_30951# uo_out[6] 0.00812f
C11594 a_59036_26247# VPWR 0.33176f
C11595 a_3172_21640# VPWR 0.20993f
C11596 _352_.A2 a_27476_23588# 0.02154f
C11597 a_61860_27912# VPWR 0.20622f
C11598 a_50436_17316# a_50524_17272# 0.28563f
C11599 a_46492_17272# a_46940_17272# 0.01288f
C11600 _340_.A2 a_26427_29977# 0.02245f
C11601 _311_.A2 _300_.ZN 0.04557f
C11602 a_4940_10567# a_5300_10664# 0.08674f
C11603 a_43804_1592# a_43804_1159# 0.05841f
C11604 a_66428_1592# a_66876_1592# 0.0131f
C11605 a_58476_10567# a_58924_10567# 0.01288f
C11606 a_4740_2824# a_4604_1592# 0.00154f
C11607 a_29804_30951# uo_out[6] 0.00233f
C11608 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN 0.63948f
C11609 a_32380_23111# a_32740_23208# 0.08707f
C11610 a_62060_23111# VPWR 0.3289f
C11611 a_20420_23208# a_20868_23208# 0.01328f
C11612 _452_.CLK a_37444_25156# 0.002f
C11613 _459_.CLK a_26160_27165# 0.00127f
C11614 _337_.A3 a_28036_26724# 0.01913f
C11615 a_33152_22091# a_33708_22505# 0.8399f
C11616 _316_.ZN a_34080_22461# 0.01766f
C11617 a_1020_6296# VPWR 0.30073f
C11618 a_60516_9476# VPWR 0.22752f
C11619 a_1020_23544# VPWR 0.30073f
C11620 a_27004_21543# a_27452_21543# 0.01288f
C11621 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN 0.02667f
C11622 a_14796_21543# a_14708_21640# 0.28563f
C11623 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I 0.00117f
C11624 a_51332_24072# a_51540_23588# 0.01751f
C11625 a_64996_2824# a_64996_1636# 0.05841f
C11626 a_2724_29480# a_2724_28292# 0.05841f
C11627 a_2812_3160# VPWR 0.30213f
C11628 a_67324_14136# VPWR 0.31547f
C11629 a_53908_26724# a_53996_26680# 0.28563f
C11630 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I VPWR 0.70858f
C11631 _474_.CLK a_55252_25156# 0.02104f
C11632 _260_.A1 _264_.B 0.29231f
C11633 a_3260_11000# VPWR 0.30487f
C11634 _287_.A1 a_32380_26247# 0.00231f
C11635 a_62560_25112# vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN 0.00466f
C11636 a_34155_25273# VPWR 0.38712f
C11637 _346_.A2 a_24304_26795# 0.00609f
C11638 a_51240_20452# VPWR 0.3154f
C11639 a_58500_2824# a_58948_2824# 0.01328f
C11640 a_28891_25273# a_29176_25273# 0.00277f
C11641 _324_.C a_49764_26724# 0.03936f
C11642 _474_.CLK a_52652_18407# 0.00706f
C11643 _474_.CLK VPWR 7.69724f
C11644 _419_.Z _474_.D 0.03293f
C11645 a_3708_26247# VPWR 0.33374f
C11646 a_33860_18884# VPWR 0.20799f
C11647 _294_.A2 a_31844_26344# 0.00265f
C11648 _359_.B a_35818_29860# 0.00222f
C11649 a_18940_2727# a_18852_2824# 0.28563f
C11650 _335_.ZN a_38584_28292# 0.0062f
C11651 a_31932_26247# a_32380_26247# 0.01222f
C11652 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_63180_26680# 0.01931f
C11653 _304_.B _265_.ZN 0.22218f
C11654 _251_.A1 a_62503_28293# 0.10506f
C11655 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN a_58588_21543# 0.00486f
C11656 _334_.A1 a_36284_29167# 0.01187f
C11657 _433_.ZN VPWR 0.48262f
C11658 a_56036_9476# a_55676_9432# 0.08717f
C11659 a_53884_9432# a_54332_9432# 0.0131f
C11660 a_67908_22020# a_67996_21976# 0.28563f
C11661 a_31484_30951# uo_out[5] 0.00309f
C11662 a_61412_14180# a_61052_14136# 0.08707f
C11663 a_64548_14180# a_64996_14180# 0.01328f
C11664 a_37584_29123# _443_.D 0.00176f
C11665 a_67117_30600# _248_.B1 0.0017f
C11666 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN a_61164_23111# 0.00306f
C11667 _250_.ZN a_62564_29032# 0.00111f
C11668 a_24392_28248# a_24780_28776# 0.00334f
C11669 _334_.A1 _362_.B 3.1106f
C11670 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN 0.0056f
C11671 a_52452_12612# a_53124_12612# 0.00347f
C11672 a_61524_13800# a_61500_12568# 0.0016f
C11673 _424_.A1 a_54916_21640# 0.00104f
C11674 _474_.CLK a_54108_21543# 0.00443f
C11675 a_49852_1159# a_50436_1256# 0.01675f
C11676 _370_.B _337_.ZN 0.07906f
C11677 _402_.ZN a_46100_26399# 0.00179f
C11678 a_31932_1159# VPWR 0.32982f
C11679 a_49204_12232# a_49316_11044# 0.02666f
C11680 a_65332_12232# a_65780_12232# 0.01328f
C11681 a_30276_1636# a_30364_1592# 0.28563f
C11682 a_26332_1592# a_26780_1592# 0.01288f
C11683 a_34308_21640# VPWR 0.23143f
C11684 _281_.ZN a_51668_23340# 0.00357f
C11685 a_55564_10567# a_55476_10664# 0.28563f
C11686 _319_.A3 _319_.A2 0.78408f
C11687 a_15492_2824# a_15492_1636# 0.05841f
C11688 a_11684_2824# a_11548_1592# 0.00154f
C11689 _349_.A4 _340_.ZN 0.74814f
C11690 _242_.Z vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN 0.00833f
C11691 a_1916_21976# VPWR 0.297f
C11692 _355_.C a_23780_26344# 0.01337f
C11693 a_35616_24776# a_36544_24419# 1.16391f
C11694 _247_.ZN VPWR 0.30355f
C11695 a_46476_20937# _416_.ZN 0.00256f
C11696 a_23892_23588# VPWR 0.20621f
C11697 a_66652_8999# VPWR 0.29679f
C11698 a_16164_29480# a_16052_28292# 0.02666f
C11699 a_61612_13703# VPWR 0.31556f
C11700 a_1380_18884# a_1020_18840# 0.08717f
C11701 a_11772_2727# VPWR 0.36383f
C11702 a_25436_21543# a_25796_21640# 0.08663f
C11703 a_3172_18884# a_3620_18884# 0.01328f
C11704 _304_.B _261_.ZN 0.00123f
C11705 _304_.B a_52988_26680# 0.02173f
C11706 a_15132_29816# uio_oe[1] 0.00435f
C11707 _459_.CLK a_16700_29383# 0.01305f
C11708 a_5052_21976# a_4940_21543# 0.02634f
C11709 a_56708_11044# VPWR 0.21151f
C11710 a_52316_15704# a_52764_15704# 0.01288f
C11711 a_28672_31048# _340_.A2 0.00226f
C11712 _325_.A1 a_43668_19668# 0.08639f
C11713 a_18096_27165# VPWR 1.09608f
C11714 _474_.Q a_47259_20127# 0.00191f
C11715 a_63876_15748# a_63964_15704# 0.28563f
C11716 _462_.D a_35728_29480# 0.24395f
C11717 a_1468_27815# VPWR 0.29679f
C11718 a_35652_26344# a_35652_25156# 0.05841f
C11719 _304_.B _398_.C 0.15966f
C11720 _255_.I _242_.Z 0.02495f
C11721 _267_.ZN vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.02667f
C11722 a_29916_2727# a_30276_2824# 0.08717f
C11723 _265_.ZN VPWR 0.96172f
C11724 _459_.CLK _351_.A2 0.0323f
C11725 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I 0.0036f
C11726 _268_.A2 a_54000_30344# 0.00265f
C11727 a_4068_23588# a_4156_23544# 0.28563f
C11728 a_17472_28363# VPWR 1.11691f
C11729 a_3172_7908# a_3260_7864# 0.28563f
C11730 ui_in[4] ui_in[5] 0.01021f
C11731 a_4068_6340# a_4156_6296# 0.28563f
C11732 a_4964_4772# a_5052_4728# 0.28563f
C11733 a_19412_20452# a_19052_20408# 0.08717f
C11734 a_20756_20452# a_21204_20452# 0.01328f
C11735 a_7092_31048# a_7068_29383# 0.00134f
C11736 _390_.ZN vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.09001f
C11737 _474_.CLK _383_.ZN 0.41755f
C11738 vgaringosc.workerclkbuff_notouch_.I a_51457_29861# 0.24228f
C11739 a_55676_27815# a_56124_27815# 0.012f
C11740 a_2364_30951# a_2724_31048# 0.08717f
C11741 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN clk 0.00868f
C11742 a_24540_1592# a_24676_1256# 0.00168f
C11743 a_5500_1592# VPWR 0.3289f
C11744 a_55812_12612# a_55900_12568# 0.28563f
C11745 _459_.CLK a_16140_25112# 0.00189f
C11746 _459_.Q a_33164_24679# 0.01328f
C11747 a_59396_12612# a_59844_12612# 0.01328f
C11748 a_4964_12612# a_4940_12135# 0.00172f
C11749 _296_.ZN uo_out[3] 0.21465f
C11750 _284_.ZN uo_out[1] 2.02722f
C11751 a_23108_24776# a_23084_23544# 0.0016f
C11752 _371_.ZN _455_.Q 0.0457f
C11753 _355_.ZN a_27900_23111# 0.00118f
C11754 a_54332_1159# VPWR 0.30141f
C11755 a_61276_1159# a_61188_1256# 0.28563f
C11756 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I 0.01006f
C11757 a_33636_1636# a_33276_1592# 0.08707f
C11758 _359_.B a_41708_30644# 0.00158f
C11759 a_63068_18840# VPWR 0.29679f
C11760 _281_.A1 _422_.ZN 0.00151f
C11761 _451_.Q a_41440_23208# 0.00371f
C11762 a_51240_20452# _424_.B2 0.04056f
C11763 a_52024_20083# _424_.ZN 0.30582f
C11764 _399_.ZN _397_.Z 0.0628f
C11765 a_42684_27815# _330_.A1 0.00839f
C11766 a_43580_27815# a_43940_27912# 0.08674f
C11767 _452_.Q a_39796_22504# 0.03005f
C11768 a_21404_1159# a_21852_1159# 0.0131f
C11769 a_66316_10567# a_66676_10664# 0.08717f
C11770 _467_.D a_15604_27912# 0.0036f
C11771 a_52340_10664# a_52788_10664# 0.01328f
C11772 _311_.A2 a_38616_24328# 0.26811f
C11773 _244_.Z a_61412_26344# 0.00292f
C11774 a_5300_24776# a_5388_23111# 0.0027f
C11775 _304_.A1 a_41488_24072# 0.11248f
C11776 _474_.CLK _424_.B2 0.08103f
C11777 _408_.ZN a_52228_27912# 0.00974f
C11778 a_29716_31048# a_29788_30345# 0.00175f
C11779 a_24788_22020# VPWR 0.20595f
C11780 _355_.C a_22100_29480# 0.00664f
C11781 _363_.Z _335_.ZN 0.70144f
C11782 _416_.A1 a_43232_29480# 0.00638f
C11783 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN a_57132_23544# 0.0071f
C11784 a_34172_2727# VPWR 0.31816f
C11785 a_24004_21640# a_24452_21640# 0.01328f
C11786 a_51332_2824# a_51420_1159# 0.0027f
C11787 a_55476_13800# VPWR 0.20622f
C11788 a_32964_18884# a_32604_18840# 0.08717f
C11789 _459_.D a_30836_23588# 0.00152f
C11790 _261_.ZN VPWR 0.40868f
C11791 _352_.A2 a_25232_27165# 0.00112f
C11792 a_22188_30951# uio_out[6] 0.00161f
C11793 a_11012_29860# VPWR 0.21215f
C11794 a_52988_26680# VPWR 0.31648f
C11795 _409_.ZN a_50996_28292# 0.00363f
C11796 a_41160_29083# uo_out[3] 1.18363f
C11797 _327_.A2 a_43668_19668# 0.08427f
C11798 a_63292_11000# VPWR 0.31389f
C11799 a_2364_15271# a_2276_15368# 0.28563f
C11800 a_21068_21976# a_20956_21543# 0.02634f
C11801 a_21852_23111# VPWR 0.31389f
C11802 _459_.CLK a_26720_30301# 0.00114f
C11803 a_3708_15271# a_4156_15271# 0.0131f
C11804 _398_.C VPWR 1.96552f
C11805 _474_.Q _419_.Z 0.67868f
C11806 a_65756_17272# a_65668_15748# 0.0027f
C11807 a_62868_23208# a_63316_23208# 0.01328f
C11808 _467_.D a_16672_26841# 0.00159f
C11809 a_41340_2727# a_41252_2824# 0.28563f
C11810 a_61500_17272# a_62084_17316# 0.01675f
C11811 a_28000_29480# a_28928_29123# 1.16391f
C11812 _264_.B _260_.A2 0.43474f
C11813 a_4604_23544# a_4516_22020# 0.0027f
C11814 a_63180_16839# a_63540_16936# 0.08717f
C11815 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN 0.02096f
C11816 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN a_58252_18407# 0.01934f
C11817 _474_.Q _399_.A2 0.48339f
C11818 a_22212_1256# a_22660_1256# 0.01328f
C11819 a_64860_9432# a_65308_9432# 0.0131f
C11820 a_67012_9476# a_66652_9432# 0.08717f
C11821 a_21428_23588# a_21876_23588# 0.01328f
C11822 a_17844_23588# a_17932_23544# 0.28563f
C11823 _281_.ZN a_47636_23588# 0.00333f
C11824 a_66204_7864# a_66652_7864# 0.0131f
C11825 a_2724_25156# a_2812_25112# 0.28563f
C11826 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I 0.00967f
C11827 a_67100_6296# a_67548_6296# 0.0131f
C11828 a_1468_2727# a_1916_2727# 0.0131f
C11829 a_51532_13703# a_51980_13703# 0.01288f
C11830 a_65532_14136# a_65420_13703# 0.02634f
C11831 _459_.Q a_31348_25156# 0.00149f
C11832 a_40580_26344# a_41028_26344# 0.01328f
C11833 a_12892_29383# a_13340_29383# 0.0131f
C11834 a_17372_30951# a_17284_31048# 0.28563f
C11835 _495_.I a_41708_30644# 0.40236f
C11836 a_19300_1636# VPWR 0.23944f
C11837 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I 0.14912f
C11838 vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN a_67908_22020# 0.00591f
C11839 a_4156_30951# a_4828_30951# 0.00544f
C11840 a_49404_12568# a_49292_12135# 0.02634f
C11841 _250_.ZN _250_.B 0.11049f
C11842 a_16700_29816# _467_.D 0.00522f
C11843 _267_.A2 _267_.A1 0.34306f
C11844 a_46716_11000# a_47164_11000# 0.01288f
C11845 a_50660_11044# a_50748_11000# 0.28563f
C11846 a_62172_15271# a_62084_15368# 0.28563f
C11847 _371_.A3 a_29680_26724# 0.00899f
C11848 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I 0.04625f
C11849 a_31172_18504# VPWR 0.20348f
C11850 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN a_61300_16936# 0.00621f
C11851 a_40132_1636# a_40580_1636# 0.01328f
C11852 a_37780_16936# a_38228_16936# 0.01328f
C11853 a_51576_25896# a_51956_26183# 0.49319f
C11854 hold1.Z a_42796_23981# 0.00489f
C11855 a_54892_24679# a_55340_24679# 0.01222f
C11856 a_2276_26724# a_2724_26724# 0.01328f
C11857 _389_.ZN _424_.A2 0.00108f
C11858 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN VPWR 0.75852f
C11859 a_55208_22505# VPWR 0.18806f
C11860 _421_.A1 _402_.B 0.06981f
C11861 _424_.B1 _384_.A1 0.40147f
C11862 a_52228_27912# _412_.A1 0.00429f
C11863 _355_.C a_26148_28776# 0.00143f
C11864 _416_.A1 a_46156_25112# 0.00192f
C11865 _365_.ZN a_35874_27937# 0.03188f
C11866 a_5052_12568# VPWR 0.33516f
C11867 a_56572_2727# VPWR 0.31411f
C11868 a_48956_30951# a_49404_30951# 0.0131f
C11869 a_64412_18407# a_64324_18504# 0.28563f
C11870 a_2276_2824# a_2724_2824# 0.01328f
C11871 _474_.CLK a_44744_26355# 0.00105f
C11872 _459_.CLK a_27884_25641# 0.01996f
C11873 _330_.A1 _319_.ZN 0.60246f
C11874 a_57580_10567# VPWR 0.32122f
C11875 a_38428_15271# a_38788_15368# 0.08717f
C11876 a_62844_2727# a_62980_1636# 0.00154f
C11877 a_28012_21976# a_27900_21543# 0.02634f
C11878 _436_.B a_41099_26841# 0.04305f
C11879 a_19524_23208# VPWR 0.23492f
C11880 a_39884_27815# VPWR 0.32564f
C11881 a_1916_28248# a_2364_28248# 0.0131f
C11882 _330_.A1 a_36860_23111# 0.01038f
C11883 a_4516_28292# a_4156_28248# 0.08674f
C11884 _427_.ZN a_53660_21543# 0.0127f
C11885 a_4964_22020# a_5052_21976# 0.28563f
C11886 a_52316_2727# a_52676_2824# 0.08717f
C11887 a_39772_20408# _325_.A2 0.00346f
C11888 a_18380_23544# a_18292_22020# 0.0027f
C11889 a_27588_26344# VPWR 0.21165f
C11890 _393_.A3 VPWR 0.76708f
C11891 a_48420_18504# a_48868_18504# 0.01328f
C11892 a_16500_25156# a_16588_25112# 0.28563f
C11893 a_20084_25156# a_20532_25156# 0.01328f
C11894 a_30388_20452# a_30028_20408# 0.08717f
C11895 a_31732_20452# a_32180_20452# 0.01328f
C11896 a_48508_13703# a_48420_13800# 0.28563f
C11897 a_62396_14136# a_62420_13800# 0.00172f
C11898 a_37084_26247# _444_.D 0.00453f
C11899 a_21292_30951# a_21740_30951# 0.01255f
C11900 a_61188_20072# vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN 0.00504f
C11901 _317_.A2 a_35088_20893# 0.00807f
C11902 a_35628_16839# a_35540_16936# 0.28563f
C11903 a_62844_11000# a_62756_9476# 0.00151f
C11904 a_25436_1592# VPWR 0.33111f
C11905 a_4852_10664# a_4964_9476# 0.02666f
C11906 _304_.B a_53996_24679# 0.00189f
C11907 a_65980_12568# a_66428_12568# 0.01288f
C11908 a_23084_29383# _343_.A2 0.00857f
C11909 a_3172_1636# a_3620_1636# 0.01328f
C11910 a_47300_1636# a_46940_1592# 0.08663f
C11911 a_54020_11044# a_53660_11000# 0.08707f
C11912 _352_.ZN a_26580_23588# 0.00212f
C11913 a_56372_12232# a_56460_10567# 0.00151f
C11914 _459_.CLK a_32096_24419# 0.00286f
C11915 a_57580_23544# VPWR 0.3467f
C11916 a_17803_26841# a_16240_26795# 0.41622f
C11917 _474_.CLK a_55252_26724# 0.00305f
C11918 a_43804_1159# a_44252_1159# 0.0131f
C11919 a_55140_20452# vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I 0.00386f
C11920 _230_.I a_60276_29032# 0.0411f
C11921 a_2724_27912# a_2724_26724# 0.05841f
C11922 a_47636_18884# VPWR 0.18975f
C11923 a_54356_20072# a_54332_18840# 0.0016f
C11924 _346_.B a_20308_27912# 0.00951f
C11925 _455_.D a_20496_26344# 0.24751f
C11926 a_19860_20452# VPWR 0.21116f
C11927 a_37386_31048# VPWR 0.01407f
C11928 a_58500_12612# VPWR 0.21771f
C11929 a_56964_26724# a_57168_26724# 0.03324f
C11930 a_932_15748# a_1380_15748# 0.01328f
C11931 a_9532_2727# a_9668_1636# 0.00154f
C11932 a_47748_15368# a_48196_15368# 0.01328f
C11933 a_11324_29383# a_11236_29480# 0.28563f
C11934 a_15692_28248# a_15692_27815# 0.05841f
C11935 a_38584_28292# a_38772_28292# 0.00257f
C11936 a_64884_26724# a_64860_26247# 0.00172f
C11937 a_51444_10664# VPWR 0.20641f
C11938 a_49852_15271# a_49764_15368# 0.28563f
C11939 _258_.I _238_.ZN 0.47213f
C11940 a_1468_5863# a_1828_5960# 0.08717f
C11941 a_2364_4295# a_2724_4392# 0.08717f
C11942 _260_.A2 a_44786_24120# 0.02198f
C11943 _389_.ZN a_46804_28292# 0.00529f
C11944 _251_.A1 a_59652_25640# 0.8066f
C11945 a_51196_15271# a_51644_15271# 0.0131f
C11946 _334_.A1 a_35914_28776# 0.00327f
C11947 a_66876_15271# VPWR 0.32932f
C11948 _393_.ZN _393_.A1 0.7567f
C11949 _452_.CLK hold2.I 0.00387f
C11950 _475_.D a_46848_20893# 0.01952f
C11951 a_53996_25112# clk 0.00335f
C11952 a_63740_2727# a_63652_2824# 0.28563f
C11953 _416_.A1 _438_.A2 0.14493f
C11954 a_14796_21976# a_15244_21976# 0.01288f
C11955 a_18740_22020# a_18828_21976# 0.28563f
C11956 a_2812_15271# VPWR 0.30213f
C11957 a_32604_16839# a_33052_16839# 0.0131f
C11958 a_48060_30951# a_47972_31048# 0.28563f
C11959 a_29156_23208# a_29244_21543# 0.00151f
C11960 a_21316_1256# VPWR 0.20348f
C11961 a_28820_24072# a_29716_23588# 0.00591f
C11962 a_44612_1256# a_45060_1256# 0.01328f
C11963 a_67100_4728# VPWR 0.29679f
C11964 a_65308_7864# VPWR 0.30378f
C11965 a_22996_25156# a_23084_25112# 0.28563f
C11966 a_23868_2727# a_24316_2727# 0.0131f
C11967 a_11772_29383# VPWR 0.3802f
C11968 a_45284_13800# a_45732_13800# 0.01328f
C11969 a_56348_14136# a_56260_12612# 0.00151f
C11970 a_59372_13703# a_59732_13800# 0.08707f
C11971 a_3260_30951# VPWR 0.31951f
C11972 _384_.A1 _218_.ZN 0.07124f
C11973 a_46156_16839# a_46516_16936# 0.08707f
C11974 _474_.CLK a_49112_29885# 0.0325f
C11975 a_64412_29816# rst_n 0.02867f
C11976 a_49652_10664# a_49628_9432# 0.0016f
C11977 a_51444_10664# a_51332_9476# 0.02666f
C11978 a_53212_12568# a_53236_12232# 0.00172f
C11979 a_36884_16936# VPWR 0.2061f
C11980 a_63292_12568# a_63404_12135# 0.02634f
C11981 a_39100_1592# VPWR 0.29679f
C11982 a_5276_1159# a_5188_1256# 0.28563f
C11983 a_53996_24679# VPWR 0.29679f
C11984 _327_.Z VPWR 1.70918f
C11985 a_38472_30169# _437_.A1 0.00141f
C11986 a_4964_29860# a_5052_29816# 0.28563f
C11987 _383_.ZN _393_.A3 0.00888f
C11988 a_1020_29816# a_1468_29816# 0.01288f
C11989 _242_.Z vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.03512f
C11990 _397_.A2 _397_.Z 0.00638f
C11991 a_31172_17316# a_31620_17316# 0.01328f
C11992 _393_.A3 a_50068_27508# 0.00323f
C11993 a_48060_30951# VPWR 0.31143f
C11994 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN a_52756_29076# 0.00423f
C11995 a_60380_11000# a_60964_11044# 0.01675f
C11996 a_1380_2824# VPWR 0.20348f
C11997 a_50212_1636# a_50300_1592# 0.28563f
C11998 a_53796_1636# a_54244_1636# 0.01328f
C11999 a_47164_11000# a_47164_10567# 0.05841f
C12000 a_51108_11044# a_51084_10567# 0.00172f
C12001 _452_.CLK a_33076_20452# 0.00932f
C12002 a_61948_27815# a_62396_27815# 0.01222f
C12003 a_30724_20072# a_30724_18884# 0.05841f
C12004 a_2364_23111# a_2812_23111# 0.0131f
C12005 a_35204_31048# _294_.ZN 0.02587f
C12006 _459_.CLK a_17036_26247# 0.00781f
C12007 a_49404_18407# a_50324_18504# 0.00795f
C12008 a_43716_2824# a_43716_1636# 0.05841f
C12009 a_51668_18504# a_51756_16839# 0.00151f
C12010 a_41572_20072# _450_.D 0.0018f
C12011 a_47524_18504# VPWR 0.20897f
C12012 _432_.ZN a_41564_24679# 0.00512f
C12013 _452_.Q a_41476_24776# 0.00157f
C12014 a_19188_25156# VPWR 0.2297f
C12015 _352_.A2 a_25436_24679# 0.00129f
C12016 a_17036_27815# a_17396_27912# 0.08717f
C12017 a_30836_20452# VPWR 0.20595f
C12018 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN _324_.C 0.0275f
C12019 a_2724_27912# a_3172_27912# 0.01328f
C12020 _359_.B uo_out[0] 0.00216f
C12021 _343_.A2 a_22996_28292# 0.00236f
C12022 a_65084_12568# VPWR 0.32121f
C12023 a_34160_20523# a_34548_20937# 0.00393f
C12024 _243_.A1 _241_.Z 0.04536f
C12025 _358_.A2 a_30036_25940# 0.00893f
C12026 a_24676_2824# a_25124_2824# 0.01328f
C12027 _437_.A1 a_37556_23588# 0.02262f
C12028 _378_.I _378_.ZN 0.76311f
C12029 a_34052_22137# VPWR 0.00264f
C12030 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I a_65668_26344# 0.00132f
C12031 a_67348_16936# VPWR 0.2061f
C12032 _447_.Q _325_.A1 0.04651f
C12033 a_46852_15368# VPWR 0.20952f
C12034 a_33476_27912# uo_out[6] 0.01944f
C12035 _268_.A2 uio_in[0] 0.00104f
C12036 _304_.B _452_.CLK 0.21238f
C12037 a_50300_15271# VPWR 0.35986f
C12038 a_45732_14180# a_46180_14180# 0.01328f
C12039 a_31708_16839# VPWR 0.29679f
C12040 a_21740_30951# a_22100_31048# 0.0869f
C12041 a_43716_1256# VPWR 0.20348f
C12042 _268_.A1 _407_.ZN 0.00439f
C12043 vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN a_58836_14180# 0.00127f
C12044 _395_.A1 clkbuf_1_0__f_clk.I 0.05023f
C12045 a_2724_13800# a_2724_12612# 0.05841f
C12046 a_16052_23208# a_16052_22020# 0.05841f
C12047 a_5052_17272# VPWR 0.33516f
C12048 _417_.A2 _473_.Q 1.96661f
C12049 a_51644_12568# a_51556_11044# 0.00151f
C12050 a_16252_1159# a_16612_1256# 0.08717f
C12051 a_60268_12135# a_60716_12135# 0.01288f
C12052 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN 0.60388f
C12053 a_52900_1636# VPWR 0.2085f
C12054 _371_.A1 a_28112_27912# 0.01262f
C12055 a_46268_12135# a_46628_12232# 0.08717f
C12056 a_61052_27815# VPWR 0.31589f
C12057 a_9444_29480# a_9892_29480# 0.01328f
C12058 a_13252_1636# a_13340_1592# 0.28563f
C12059 a_9308_1592# a_9756_1592# 0.01288f
C12060 _304_.ZN _328_.A2 0.00992f
C12061 a_58687_31220# _270_.A2 0.04371f
C12062 a_58911_30644# a_59143_31198# 0.00209f
C12063 _230_.I _249_.A2 0.26937f
C12064 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I 0.05664f
C12065 a_31396_31048# _223_.I 0.01053f
C12066 a_54020_15368# a_54020_14180# 0.05841f
C12067 _350_.A2 _359_.B 0.23911f
C12068 a_23780_2824# VPWR 0.22423f
C12069 a_58052_11044# a_58028_10567# 0.00172f
C12070 a_54108_11000# a_54220_10567# 0.02634f
C12071 a_29468_1592# a_29468_1159# 0.05841f
C12072 a_67684_11044# a_67772_11000# 0.28563f
C12073 a_46628_31048# a_47076_31048# 0.01328f
C12074 _301_.A1 a_38784_22504# 0.00194f
C12075 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN 0.73131f
C12076 ui_in[6] ui_in[5] 0.01021f
C12077 _397_.Z a_48308_23588# 0.19087f
C12078 a_1468_23111# a_1380_23208# 0.28563f
C12079 _327_.A2 a_40668_19975# 0.00435f
C12080 a_5388_24679# a_5300_24776# 0.28563f
C12081 _448_.Q a_42784_22504# 0.0013f
C12082 a_22748_24679# a_23196_24679# 0.01288f
C12083 a_1380_9096# a_1828_9096# 0.01328f
C12084 a_66204_1159# a_66652_1159# 0.01255f
C12085 a_30812_19975# a_31260_19975# 0.0131f
C12086 a_36960_27912# _443_.D 0.31063f
C12087 _350_.A1 a_30388_28776# 0.02087f
C12088 a_2276_7528# a_2724_7528# 0.01328f
C12089 a_3172_5960# a_3620_5960# 0.01328f
C12090 a_5052_14136# VPWR 0.33516f
C12091 _424_.B1 clk 0.75172f
C12092 a_4068_4392# a_4852_4392# 0.00276f
C12093 a_1468_18407# a_1828_18504# 0.08717f
C12094 a_32156_18407# a_32604_18407# 0.0131f
C12095 a_27328_25227# a_28208_25641# 0.00306f
C12096 a_33376_23659# a_34304_24029# 1.16391f
C12097 a_53908_25156# a_54356_25156# 0.01328f
C12098 _260_.A1 a_44038_21236# 0.00758f
C12099 a_59372_12135# VPWR 0.31389f
C12100 a_8548_29480# VPWR 0.22423f
C12101 a_35292_15704# a_35740_15704# 0.01288f
C12102 a_45508_31048# VPWR 0.20364f
C12103 _365_.ZN _288_.ZN 0.06495f
C12104 _419_.Z a_51196_21543# 0.0028f
C12105 _474_.CLK a_53996_26680# 0.05962f
C12106 _431_.A3 a_39587_24372# 0.00455f
C12107 a_59620_27208# a_59828_26724# 0.02745f
C12108 a_21852_24679# VPWR 0.3142f
C12109 a_46492_15704# a_46492_15271# 0.05841f
C12110 a_50436_15748# a_50300_15271# 0.00168f
C12111 a_1380_7528# VPWR 0.20348f
C12112 a_3172_4392# VPWR 0.20993f
C12113 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_61076_23208# 0.02721f
C12114 _447_.Q _327_.A2 0.01723f
C12115 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I 0.63963f
C12116 a_45396_28292# a_45484_28248# 0.28563f
C12117 _417_.A2 _475_.D 0.03842f
C12118 a_34396_15704# VPWR 0.33659f
C12119 _452_.CLK VPWR 7.56333f
C12120 a_51240_19624# a_49896_18909# 0.00173f
C12121 _267_.A1 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.31028f
C12122 a_40464_27165# a_41099_26841# 0.02112f
C12123 a_51308_18407# a_51756_18407# 0.0131f
C12124 a_28460_21976# a_28908_21976# 0.01288f
C12125 _230_.I a_62564_29032# 0.49871f
C12126 _474_.CLK a_55788_24679# 0.02256f
C12127 _330_.A1 a_37360_19325# 0.01489f
C12128 a_54444_16839# a_54892_16839# 0.012f
C12129 a_50412_18407# VPWR 0.34813f
C12130 a_52452_14180# a_53124_14180# 0.00347f
C12131 a_65892_15368# a_65892_14180# 0.05841f
C12132 a_22996_28292# a_22636_28248# 0.08674f
C12133 _452_.CLK a_44364_17272# 0.00614f
C12134 a_47297_25596# _279_.Z 0.50602f
C12135 a_53548_16839# VPWR 0.31389f
C12136 _421_.A1 a_46352_22021# 0.12746f
C12137 a_66116_1256# VPWR 0.23483f
C12138 a_67012_1256# a_67460_1256# 0.01328f
C12139 a_46044_2727# a_46716_2727# 0.00544f
C12140 a_67124_13800# a_67572_13800# 0.01328f
C12141 a_50996_13800# a_51108_12612# 0.02666f
C12142 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN _408_.ZN 0.00158f
C12143 a_47164_18407# a_47300_17316# 0.00154f
C12144 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN VPWR 0.75536f
C12145 _260_.A1 a_41564_24679# 0.01362f
C12146 _304_.B a_41116_26247# 0.01784f
C12147 a_23108_23208# a_22996_22020# 0.02666f
C12148 _294_.A2 a_31920_29480# 0.04331f
C12149 a_59036_1592# VPWR 0.29679f
C12150 a_27676_1159# a_27588_1256# 0.28563f
C12151 a_57580_12135# a_57492_12232# 0.28563f
C12152 a_16028_1592# a_16700_1592# 0.00544f
C12153 a_40316_23233# VPWR 0.01199f
C12154 a_14684_29816# a_15132_29816# 0.01288f
C12155 a_14796_21543# VPWR 0.30073f
C12156 _448_.Q a_40244_21640# 0.00133f
C12157 _228_.ZN _324_.C 0.01906f
C12158 _474_.CLK a_57120_31048# 0.00898f
C12159 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I 0.78095f
C12160 a_47164_10567# a_47612_10567# 0.0131f
C12161 a_64996_11044# a_64972_10567# 0.00172f
C12162 a_59932_1592# a_60380_1592# 0.01288f
C12163 _260_.A1 _325_.A2 0.03365f
C12164 a_45956_2824# VPWR 0.20968f
C12165 _252_.ZN _244_.Z 0.53734f
C12166 _300_.ZN a_38764_20408# 0.00134f
C12167 a_21404_23111# a_21764_23208# 0.08707f
C12168 a_62308_26344# vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN 0.00149f
C12169 a_33276_23111# a_33724_23111# 0.012f
C12170 a_47948_23111# _324_.B 0.05473f
C12171 a_24988_24679# a_25348_24776# 0.08707f
C12172 _334_.A1 _402_.A1 0.00248f
C12173 a_49092_9476# VPWR 0.23086f
C12174 a_15692_21543# a_16140_21543# 0.0131f
C12175 a_62396_27815# a_62308_27912# 0.28563f
C12176 a_21204_31048# VPWR 0.19631f
C12177 a_59284_14180# VPWR 0.20697f
C12178 a_42596_15748# a_42236_15704# 0.08707f
C12179 _330_.A1 a_36996_21640# 0.00114f
C12180 a_1468_29816# a_1468_29383# 0.05841f
C12181 a_53236_12232# VPWR 0.20622f
C12182 a_5412_29860# a_5276_29383# 0.00168f
C12183 _411_.A2 _474_.Q 0.00205f
C12184 a_47076_2824# a_47524_2824# 0.01328f
C12185 a_58836_18884# a_58924_18840# 0.28563f
C12186 a_26756_24801# VPWR 0.01272f
C12187 a_25652_31048# _340_.A2 0.01225f
C12188 _250_.B a_63524_29098# 0.00164f
C12189 a_10876_29383# uio_oe[4] 0.00107f
C12190 a_7516_2727# a_7428_2824# 0.28563f
C12191 _447_.Q a_37084_21543# 0.01738f
C12192 a_48196_15748# VPWR 0.20595f
C12193 a_33948_19975# a_34644_20072# 0.01227f
C12194 a_31088_30301# VPWR 0.52849f
C12195 _397_.A1 clkbuf_1_0__f_clk.I 0.57202f
C12196 _378_.I uio_out[6] 0.049f
C12197 _237_.A1 a_60401_30300# 0.5712f
C12198 a_49988_9476# a_50436_9476# 0.01328f
C12199 a_22100_31048# a_22548_31048# 0.01328f
C12200 _452_.CLK a_36100_26344# 0.00782f
C12201 _248_.B1 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I 0.00281f
C12202 a_56260_14180# a_56348_14136# 0.28563f
C12203 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN a_64212_23588# 0.00102f
C12204 uo_out[5] uo_out[4] 0.08256f
C12205 ui_in[3] ui_in[1] 0.00561f
C12206 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN VPWR 0.80003f
C12207 a_10204_1592# a_10340_1256# 0.00168f
C12208 _400_.ZN _381_.A2 0.08688f
C12209 a_57940_13800# a_58052_12612# 0.02666f
C12210 a_54132_13800# a_54108_12568# 0.0016f
C12211 a_41099_26841# a_41564_26247# 0.02319f
C12212 _427_.A2 _424_.A1 0.47564f
C12213 VPWR uio_in[6] 0.00621f
C12214 a_41116_26247# VPWR 0.32721f
C12215 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN 0.01319f
C12216 a_1380_24776# a_1380_23588# 0.05841f
C12217 a_9084_1159# VPWR 0.3289f
C12218 a_38428_1159# a_39012_1256# 0.01675f
C12219 _436_.B a_41476_24776# 0.00762f
C12220 uio_oe[0] uio_out[7] 0.06851f
C12221 a_54132_12232# a_54580_12232# 0.01328f
C12222 a_932_4772# a_1380_4772# 0.01328f
C12223 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I 0.00171f
C12224 a_22972_1592# a_23420_1592# 0.01288f
C12225 a_51980_12135# a_52004_11044# 0.0016f
C12226 _305_.A2 _402_.B 0.00935f
C12227 _436_.ZN a_40468_25157# 0.00129f
C12228 a_58588_26247# VPWR 0.33759f
C12229 _244_.Z a_61500_26247# 0.00302f
C12230 a_2724_21640# VPWR 0.20782f
C12231 a_50436_17316# a_50076_17272# 0.08707f
C12232 a_61412_27912# VPWR 0.20862f
C12233 a_4940_10567# a_4852_10664# 0.28563f
C12234 _340_.A2 a_26720_30301# 0.02209f
C12235 a_932_1636# VPWR 0.22176f
C12236 _287_.A2 _352_.A2 0.04231f
C12237 a_43916_29816# _480_.Q 0.00497f
C12238 a_45012_29816# a_43232_29480# 0.00705f
C12239 _334_.A1 _359_.B 0.29093f
C12240 _459_.CLK a_24860_27209# 0.00157f
C12241 _402_.A1 a_49652_29480# 0.06521f
C12242 a_47524_31048# _474_.CLK 0.00156f
C12243 a_32380_23111# a_32292_23208# 0.28563f
C12244 a_61612_23111# VPWR 0.32897f
C12245 _311_.A2 a_38852_25156# 0.00491f
C12246 _452_.CLK a_36996_25156# 0.00224f
C12247 a_33152_22091# a_34080_22461# 1.16391f
C12248 a_59932_9432# VPWR 0.33981f
C12249 a_4964_23588# VPWR 0.21167f
C12250 _337_.A3 a_27588_26724# 0.01705f
C12251 a_54040_22366# a_54824_22045# 0.02307f
C12252 a_2364_3160# VPWR 0.30029f
C12253 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN 0.01057f
C12254 a_4964_6340# VPWR 0.21167f
C12255 a_52988_26680# a_53996_26680# 0.00323f
C12256 a_66876_14136# VPWR 0.31547f
C12257 _416_.A1 _402_.ZN 0.00342f
C12258 _474_.CLK a_54804_25156# 0.02341f
C12259 _397_.A2 _284_.B 0.31576f
C12260 a_2812_11000# VPWR 0.30213f
C12261 _474_.Q _399_.ZN 0.30289f
C12262 a_34448_25597# VPWR 0.75781f
C12263 a_49092_15748# a_49540_15748# 0.01328f
C12264 a_50748_20408# VPWR 0.34043f
C12265 _346_.A2 a_21600_26725# 0.11907f
C12266 _441_.ZN _301_.A1 0.00174f
C12267 a_65308_19975# a_65220_20072# 0.28563f
C12268 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN VPWR 0.7401f
C12269 _474_.CLK a_52204_18407# 0.00718f
C12270 _422_.ZN a_52997_20936# 0.00117f
C12271 a_30795_29977# a_31040_30345# 0.00232f
C12272 a_33412_18884# VPWR 0.20644f
C12273 a_52639_30644# VPWR 0.31337f
C12274 _359_.B a_35156_29860# 0.00139f
C12275 a_3260_26247# VPWR 0.30487f
C12276 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62732_26680# 0.01884f
C12277 a_18492_2727# a_18852_2824# 0.08717f
C12278 _304_.B a_41440_28363# 0.06826f
C12279 _260_.A2 a_44038_21236# 0.05147f
C12280 _334_.A1 a_36656_29123# 0.00393f
C12281 a_55588_9476# a_55676_9432# 0.28563f
C12282 _294_.ZN _335_.ZN 0.08684f
C12283 _362_.ZN _223_.ZN 0.01755f
C12284 a_26668_21976# a_26580_20452# 0.00151f
C12285 a_60964_14180# a_61052_14136# 0.28563f
C12286 a_50300_14136# a_50188_13703# 0.02634f
C12287 a_53212_17272# a_53124_15748# 0.00151f
C12288 a_4156_20408# a_4604_20408# 0.01222f
C12289 _428_.Z _427_.B1 0.0057f
C12290 _230_.I _250_.B 1.07586f
C12291 _455_.Q _346_.A2 1.72337f
C12292 a_48508_12568# a_48956_12568# 0.01288f
C12293 a_52452_12612# a_52540_12568# 0.28563f
C12294 a_64884_13800# a_64996_12612# 0.02666f
C12295 _460_.D a_33188_25940# 0.1116f
C12296 _411_.A2 _395_.A2 0.20813f
C12297 _424_.A1 a_54468_21640# 0.00275f
C12298 a_19076_24776# a_19188_23588# 0.02666f
C12299 a_31484_1159# VPWR 0.33352f
C12300 a_49852_1159# a_49764_1256# 0.28563f
C12301 _474_.CLK a_53660_21543# 0.00119f
C12302 _287_.A1 _293_.A2 0.3666f
C12303 _252_.ZN a_59605_25962# 0.00602f
C12304 a_30276_1636# a_29916_1592# 0.08707f
C12305 _330_.A1 a_36212_23588# 0.00134f
C12306 a_58924_12135# a_58948_11044# 0.0016f
C12307 _403_.ZN _470_.D 0.44912f
C12308 _304_.A1 _316_.A3 0.02998f
C12309 a_33636_21640# VPWR 0.21566f
C12310 a_34308_26344# a_35204_26344# 0.00455f
C12311 _281_.ZN a_51428_23340# 0.00151f
C12312 _438_.A2 _431_.A3 0.8676f
C12313 a_55116_10567# a_55476_10664# 0.08707f
C12314 a_1380_10664# a_1828_10664# 0.01328f
C12315 _424_.A1 a_52228_19368# 0.1637f
C12316 a_9980_1159# a_10428_1159# 0.0131f
C12317 a_43668_19668# VPWR 1.39729f
C12318 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN a_61188_20072# 0.07119f
C12319 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I 0.10027f
C12320 a_30948_23208# a_31396_23208# 0.01328f
C12321 _355_.C a_23332_26344# 0.01633f
C12322 _260_.A2 a_41564_24679# 0.04505f
C12323 a_1468_21976# VPWR 0.29679f
C12324 _402_.A1 a_41140_27912# 0.00546f
C12325 a_66204_8999# VPWR 0.31657f
C12326 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_56720_26344# 0.00172f
C12327 a_932_18884# a_1020_18840# 0.28563f
C12328 a_932_5960# VPWR 0.22176f
C12329 a_25436_21543# a_25348_21640# 0.28563f
C12330 a_23444_23588# VPWR 0.20665f
C12331 a_3620_21640# a_4068_21640# 0.01328f
C12332 a_61164_13703# VPWR 0.31556f
C12333 a_11324_2727# VPWR 0.32798f
C12334 a_39908_2824# a_39996_1159# 0.0027f
C12335 _355_.C a_17860_28777# 0.00103f
C12336 a_62308_27912# a_62756_27912# 0.01328f
C12337 _304_.B a_50176_26724# 0.00761f
C12338 a_56260_11044# VPWR 0.20595f
C12339 _459_.CLK a_16252_29383# 0.0041f
C12340 _325_.A1 a_43444_19668# 0.00312f
C12341 _282_.ZN _281_.ZN 0.38455f
C12342 a_17803_26841# VPWR 0.54588f
C12343 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I _256_.A2 0.08393f
C12344 a_1020_27815# VPWR 0.30073f
C12345 a_63876_15748# a_63516_15704# 0.08717f
C12346 a_66564_15748# a_67012_15748# 0.01328f
C12347 _265_.ZN a_41099_26841# 0.00521f
C12348 _323_.A3 a_38788_20072# 0.05218f
C12349 a_62508_23111# a_62956_23111# 0.0131f
C12350 a_29916_2727# a_29828_2824# 0.28563f
C12351 a_24228_26344# a_24080_25227# 0.00179f
C12352 a_41440_28363# VPWR 1.14095f
C12353 a_62420_22020# vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I 0.00293f
C12354 _375_.Z _346_.B 0.19669f
C12355 a_60964_9476# a_61412_9476# 0.01328f
C12356 a_4068_23588# a_3708_23544# 0.08717f
C12357 a_1468_23544# a_1916_23544# 0.0131f
C12358 a_10788_1256# a_11236_1256# 0.01328f
C12359 a_3172_7908# a_2812_7864# 0.08717f
C12360 a_2364_4728# a_2812_4728# 0.0131f
C12361 a_4964_4772# a_4604_4728# 0.08674f
C12362 a_4068_6340# a_3708_6296# 0.08717f
C12363 a_1468_6296# a_1916_6296# 0.0131f
C12364 a_3260_3160# a_3708_3160# 0.0131f
C12365 _390_.ZN a_50996_28292# 0.01526f
C12366 a_57692_14136# a_57580_13703# 0.02634f
C12367 a_18964_20452# a_19052_20408# 0.28563f
C12368 a_67884_16839# a_67908_15748# 0.0016f
C12369 a_2364_30951# a_2276_31048# 0.28563f
C12370 a_1468_29383# a_1916_29383# 0.0131f
C12371 a_57020_23111# clk 0.00133f
C12372 a_5052_1592# VPWR 0.3289f
C12373 _324_.C a_43736_25896# 0.04401f
C12374 _459_.Q a_32096_24419# 0.19507f
C12375 a_58388_13800# a_58476_12135# 0.00151f
C12376 a_2364_12568# a_2364_12135# 0.05841f
C12377 a_55812_12612# a_55452_12568# 0.08707f
C12378 _296_.ZN _388_.B 0.01265f
C12379 _395_.A2 _399_.ZN 0.11967f
C12380 _433_.ZN a_39796_22504# 0.00664f
C12381 _452_.Q _304_.ZN 0.26024f
C12382 _459_.CLK _358_.A3 0.1179f
C12383 _324_.B a_48529_22460# 0.04458f
C12384 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN 0.0847f
C12385 a_53660_1159# VPWR 0.35728f
C12386 a_60828_1159# a_61188_1256# 0.08717f
C12387 a_32592_25227# a_33472_25641# 0.00306f
C12388 a_35652_25156# a_36100_25156# 0.01328f
C12389 a_3708_11000# a_4156_11000# 0.0131f
C12390 _281_.A1 a_51108_21640# 0.00438f
C12391 a_65868_12135# a_65892_11044# 0.0016f
C12392 a_55924_12232# a_55812_11044# 0.02666f
C12393 a_62620_18840# VPWR 0.29679f
C12394 a_1380_16936# a_1828_16936# 0.01328f
C12395 a_33188_1636# a_33276_1592# 0.28563f
C12396 a_36772_1636# a_37220_1636# 0.01328f
C12397 _451_.Q a_41216_23208# 0.00909f
C12398 a_43580_27815# a_43492_27912# 0.28563f
C12399 a_42236_27815# _330_.A1 0.00692f
C12400 _399_.ZN a_46984_23588# 0.01244f
C12401 _451_.Q _325_.A1 0.11296f
C12402 _467_.D a_15156_27912# 0.00187f
C12403 _244_.Z a_60964_26344# 0.00843f
C12404 a_31620_18504# a_31620_17316# 0.05841f
C12405 a_66316_10567# a_66228_10664# 0.28563f
C12406 _251_.ZN VPWR 0.47766f
C12407 _336_.Z a_30724_26020# 0.16423f
C12408 a_24340_22020# VPWR 0.20595f
C12409 _355_.C a_21652_29480# 0.00657f
C12410 a_32516_18884# a_32604_18840# 0.28563f
C12411 a_55028_13800# VPWR 0.20622f
C12412 a_33724_2727# VPWR 0.31592f
C12413 a_4156_26247# a_4940_26247# 0.00443f
C12414 a_21740_30951# uio_out[6] 0.00321f
C12415 _327_.A2 a_43444_19668# 0.00185f
C12416 a_50176_26724# VPWR 0.01009f
C12417 a_54892_25112# a_55340_25112# 0.01255f
C12418 a_10564_29860# VPWR 0.21103f
C12419 a_62196_16936# a_62084_15748# 0.02666f
C12420 a_62844_11000# VPWR 0.31389f
C12421 a_1916_15271# a_2276_15368# 0.08717f
C12422 _287_.A2 _223_.ZN 0.08965f
C12423 _437_.ZN _301_.A1 0.01627f
C12424 a_21404_23111# VPWR 0.31389f
C12425 _459_.CLK a_25420_30345# 0.00163f
C12426 _261_.ZN a_39780_22805# 0.0228f
C12427 _384_.A3 _399_.A1 0.00232f
C12428 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN VPWR 0.93109f
C12429 _325_.ZN a_43916_16839# 0.00152f
C12430 _268_.A2 _274_.ZN 0.48722f
C12431 a_40892_2727# a_41252_2824# 0.08717f
C12432 a_63180_16839# a_63092_16936# 0.28563f
C12433 _281_.ZN a_47412_23588# 0.00839f
C12434 _474_.Q a_48516_24080# 0.00541f
C12435 a_66564_9476# a_66652_9432# 0.28563f
C12436 a_17844_23588# a_17484_23544# 0.08707f
C12437 a_16164_31048# uio_oe[1] 0.00802f
C12438 a_4516_25156# a_4964_25156# 0.01328f
C12439 a_2724_25156# a_2364_25112# 0.08717f
C12440 _435_.A3 _436_.ZN 0.13128f
C12441 a_54556_14136# a_54580_13800# 0.00172f
C12442 a_66004_20072# a_66116_18884# 0.02666f
C12443 a_24204_20408# a_24652_20408# 0.0131f
C12444 _459_.Q a_31124_25156# 0.00323f
C12445 a_16916_31048# a_17284_31048# 0.02601f
C12446 a_66652_17272# a_66540_16839# 0.02634f
C12447 a_57244_11000# a_57156_9476# 0.00151f
C12448 a_18852_1636# VPWR 0.21061f
C12449 a_62308_12612# a_62756_12612# 0.01328f
C12450 a_61297_30300# ui_in[2] 0.00638f
C12451 _324_.C _417_.A2 0.0258f
C12452 _452_.CLK _260_.ZN 0.11647f
C12453 _407_.ZN _398_.C 0.01389f
C12454 a_50660_11044# a_50300_11000# 0.08707f
C12455 a_61724_15271# a_62084_15368# 0.08717f
C12456 _371_.A3 a_28596_26725# 0.00102f
C12457 a_62868_12232# a_62756_11044# 0.02666f
C12458 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I a_58588_21543# 0.01035f
C12459 a_30724_18504# VPWR 0.22176f
C12460 _268_.A1 _274_.A2 0.55476f
C12461 _451_.Q _327_.A2 0.0415f
C12462 _284_.B a_48988_26369# 0.00117f
C12463 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN 0.08726f
C12464 a_32380_1159# a_32828_1159# 0.0131f
C12465 a_55312_22340# VPWR 0.39596f
C12466 a_62868_10664# a_63316_10664# 0.01328f
C12467 a_24900_24776# a_24988_23111# 0.00151f
C12468 a_25572_2824# a_25436_1592# 0.00154f
C12469 a_29380_2824# a_29380_1636# 0.05841f
C12470 a_66988_18407# a_67012_17316# 0.0016f
C12471 _384_.ZN _392_.A2 0.37564f
C12472 a_15244_26680# a_15244_26247# 0.05841f
C12473 _397_.A2 _474_.Q 0.11231f
C12474 a_37291_29535# a_37584_29123# 0.49241f
C12475 a_56124_2727# VPWR 0.31143f
C12476 a_62308_2824# a_62396_1159# 0.0027f
C12477 hold2.I _447_.Q 0.00769f
C12478 a_4604_12568# VPWR 0.33016f
C12479 a_63964_18407# a_64324_18504# 0.08717f
C12480 a_19612_26247# a_19524_26344# 0.28563f
C12481 a_36324_15368# a_36772_15368# 0.01328f
C12482 _416_.A1 a_46716_18407# 0.00136f
C12483 a_57132_10567# VPWR 0.32337f
C12484 _330_.A1 a_34160_20523# 0.06476f
C12485 _459_.CLK a_28256_25597# 0.01231f
C12486 a_38428_15271# a_38340_15368# 0.28563f
C12487 a_58252_16839# a_58700_16839# 0.01222f
C12488 a_19076_23208# VPWR 0.21778f
C12489 _436_.B a_41392_27165# 0.19704f
C12490 _373_.ZN _371_.A1 0.00108f
C12491 a_39772_15271# a_40220_15271# 0.0131f
C12492 _274_.A3 _267_.A2 0.4173f
C12493 a_38816_27555# VPWR 0.51085f
C12494 _261_.ZN a_39796_22504# 0.85252f
C12495 _260_.A1 _302_.Z 0.0246f
C12496 _460_.Q uo_out[4] 0.0607f
C12497 a_4068_28292# a_4156_28248# 0.28563f
C12498 a_52316_2727# a_52228_2824# 0.28563f
C12499 a_4964_22020# a_4604_21976# 0.08674f
C12500 a_2364_21976# a_2812_21976# 0.0131f
C12501 _237_.A1 a_60852_28292# 0.00142f
C12502 a_63964_17272# a_64412_17272# 0.0131f
C12503 a_27140_26344# VPWR 0.24076f
C12504 a_24340_23588# a_24788_23588# 0.01328f
C12505 a_67100_8999# a_67548_8999# 0.0131f
C12506 a_53212_29816# _274_.A3 0.00128f
C12507 a_33188_1256# a_33636_1256# 0.01328f
C12508 _441_.A2 _305_.A2 0.62753f
C12509 a_16500_25156# a_16140_25112# 0.08707f
C12510 a_2812_18840# a_2812_18407# 0.05841f
C12511 a_48060_13703# a_48420_13800# 0.08717f
C12512 a_62060_13703# a_62508_13703# 0.01288f
C12513 a_52540_14136# a_52452_12612# 0.00151f
C12514 a_12444_2727# a_12892_2727# 0.0131f
C12515 a_29940_20452# a_30028_20408# 0.28563f
C12516 a_36636_26247# _444_.D 0.00453f
C12517 _325_.A2 a_44276_20072# 0.10875f
C12518 a_35180_16839# a_35540_16936# 0.08707f
C12519 _268_.A1 a_56260_31048# 0.00322f
C12520 a_58063_30644# a_58911_30644# 0.00337f
C12521 a_24988_1592# VPWR 0.3289f
C12522 _330_.A1 a_38764_16839# 0.02422f
C12523 a_55900_12568# a_56012_12135# 0.02634f
C12524 a_16916_31048# a_17372_30951# 0.0065f
C12525 _304_.B a_53548_24679# 0.00379f
C12526 a_59844_12612# a_59820_12135# 0.00172f
C12527 a_1468_25112# a_1468_24679# 0.05841f
C12528 _304_.B a_40668_19975# 0.00283f
C12529 a_67117_30600# a_67741_30600# 0.10419f
C12530 _473_.Q a_45920_20523# 0.00103f
C12531 a_66900_18504# a_67348_18504# 0.01328f
C12532 _251_.A1 _250_.A2 0.084f
C12533 a_53572_11044# a_53660_11000# 0.28563f
C12534 a_57156_11044# a_57604_11044# 0.01328f
C12535 a_15132_1592# a_15132_1159# 0.05841f
C12536 a_42908_1592# a_43356_1592# 0.01288f
C12537 a_46852_1636# a_46940_1592# 0.28563f
C12538 _330_.A1 a_36996_17316# 0.0015f
C12539 a_48308_16936# a_48756_16936# 0.01328f
C12540 _395_.A3 _476_.Q 0.02465f
C12541 _371_.A1 a_28124_26680# 0.01448f
C12542 _337_.ZN _336_.Z 0.09991f
C12543 _459_.CLK a_31803_24831# 0.00131f
C12544 a_57132_23544# VPWR 0.32074f
C12545 _304_.A1 a_40656_23588# 0.00241f
C12546 a_19860_26724# a_20308_26724# 0.01328f
C12547 _474_.CLK a_54804_26724# 0.00591f
C12548 a_59172_23208# a_59172_22020# 0.05841f
C12549 a_58476_17272# a_58612_16936# 0.00168f
C12550 a_45820_18840# VPWR 0.33116f
C12551 _399_.ZN _427_.A2 0.24436f
C12552 _441_.A2 a_41440_23208# 0.00425f
C12553 _424_.A2 _384_.A1 0.09144f
C12554 a_20844_26680# a_20496_26344# 0.0074f
C12555 _346_.B a_19860_27912# 0.00169f
C12556 a_53616_29480# a_52756_29076# 0.00475f
C12557 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN a_56148_24776# 0.00459f
C12558 a_1916_27815# a_2364_27815# 0.0131f
C12559 _304_.B _447_.Q 0.0618f
C12560 a_19412_20452# VPWR 0.24625f
C12561 _275_.A2 a_50996_28292# 0.01776f
C12562 a_58052_12612# VPWR 0.2295f
C12563 a_56964_26724# a_56816_26724# 0.00128f
C12564 _359_.B _370_.ZN 0.22689f
C12565 _223_.I _294_.ZN 0.67965f
C12566 a_13252_2824# a_13700_2824# 0.01328f
C12567 _369_.ZN _371_.A1 1.15525f
C12568 _416_.A1 _384_.ZN 0.66913f
C12569 _395_.A1 _408_.ZN 0.00977f
C12570 a_10876_29383# a_11236_29480# 0.08717f
C12571 _474_.Q a_48308_23588# 0.06894f
C12572 a_36100_15748# a_35964_15271# 0.00168f
C12573 a_32156_15704# a_32156_15271# 0.05841f
C12574 a_50996_10664# VPWR 0.20977f
C12575 a_49180_15271# a_49764_15368# 0.01675f
C12576 a_57220_29861# _258_.ZN 0.00452f
C12577 a_1468_5863# a_1380_5960# 0.28563f
C12578 a_2364_4295# a_2276_4392# 0.28563f
C12579 a_932_21640# a_932_20452# 0.05841f
C12580 a_36188_26680# a_36636_26680# 0.01255f
C12581 _260_.A2 a_44162_24120# 0.06172f
C12582 _389_.ZN a_46580_28292# 0.01394f
C12583 _393_.ZN a_47525_29480# 0.00209f
C12584 _290_.ZN a_34292_28776# 0.00142f
C12585 _334_.A1 a_35710_28776# 0.00446f
C12586 _237_.A1 _238_.I 0.38236f
C12587 _404_.A1 _397_.A4 0.07707f
C12588 a_66428_15271# VPWR 0.3352f
C12589 _475_.D a_45920_20523# 0.27071f
C12590 a_18740_22020# a_18380_21976# 0.08707f
C12591 a_2364_15271# VPWR 0.30029f
C12592 a_63292_2727# a_63652_2824# 0.08717f
C12593 a_66788_15368# a_67236_15368# 0.01328f
C12594 a_47612_30951# a_47972_31048# 0.08717f
C12595 a_64860_7864# VPWR 0.30145f
C12596 a_20868_1256# VPWR 0.20348f
C12597 _325_.A2 a_37067_19001# 0.02582f
C12598 a_66652_4728# VPWR 0.29679f
C12599 a_22996_25156# a_22636_25112# 0.08674f
C12600 a_59372_13703# a_59284_13800# 0.28563f
C12601 _435_.A3 _439_.ZN 0.01511f
C12602 a_11324_29383# VPWR 0.34575f
C12603 a_2812_30951# VPWR 0.31677f
C12604 _474_.Q a_47860_21640# 0.00147f
C12605 a_46156_16839# a_46068_16936# 0.28563f
C12606 a_38652_1592# VPWR 0.32982f
C12607 a_4828_1159# a_5188_1256# 0.08717f
C12608 a_36436_16936# VPWR 0.2061f
C12609 a_49292_12135# a_49740_12135# 0.01288f
C12610 a_66788_12612# a_66764_12135# 0.00172f
C12611 a_53548_24679# VPWR 0.32888f
C12612 a_5948_1592# a_6396_1592# 0.01288f
C12613 a_17484_25112# a_17484_24679# 0.05841f
C12614 _242_.Z a_56404_27208# 0.00197f
C12615 a_40668_19975# VPWR 0.3094f
C12616 a_21428_25156# a_21404_24679# 0.00172f
C12617 _397_.A2 a_46984_23588# 0.5208f
C12618 a_4964_29860# a_4604_29816# 0.08707f
C12619 _304_.B vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.12792f
C12620 a_47612_30951# VPWR 0.31143f
C12621 a_67124_12232# a_67212_10567# 0.00151f
C12622 a_50212_1636# a_49852_1592# 0.08707f
C12623 _433_.ZN a_41476_24776# 0.00498f
C12624 _267_.A2 _324_.C 0.94364f
C12625 _452_.CLK a_32628_20452# 0.00245f
C12626 a_48284_15271# a_48420_14180# 0.00154f
C12627 a_2364_24679# a_2812_24679# 0.0131f
C12628 a_54780_1159# a_55228_1159# 0.0131f
C12629 _459_.CLK a_16588_26247# 0.00814f
C12630 a_67908_18884# a_67996_18840# 0.28563f
C12631 a_47076_18504# VPWR 0.20897f
C12632 a_63516_18840# a_63964_18840# 0.0131f
C12633 _362_.B _335_.ZN 2.42405f
C12634 _378_.I a_18096_27165# 0.00735f
C12635 a_18740_25156# VPWR 0.21333f
C12636 a_64212_23588# vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN 0.00126f
C12637 a_30388_20452# VPWR 0.20595f
C12638 a_17036_27815# a_16948_27912# 0.28563f
C12639 _447_.Q VPWR 2.78121f
C12640 _343_.A2 a_22548_28292# 0.00118f
C12641 _402_.A1 _234_.ZN 0.06557f
C12642 _245_.I1 clk 0.09342f
C12643 a_32068_15748# a_32516_15748# 0.01328f
C12644 a_64636_12568# VPWR 0.33393f
C12645 a_34160_20523# a_35723_20569# 0.41635f
C12646 _395_.A1 _412_.A1 0.40798f
C12647 a_45732_18504# a_45708_17272# 0.0016f
C12648 _243_.A1 a_57244_27815# 0.00235f
C12649 _402_.A1 a_49044_28292# 0.00148f
C12650 a_62564_29032# a_62944_29101# 0.00372f
C12651 _437_.A1 a_37108_23588# 0.00397f
C12652 _378_.I a_17472_28363# 0.02586f
C12653 a_37868_16839# a_37892_15748# 0.0016f
C12654 a_48104_30219# _397_.A2 0.25643f
C12655 a_66900_16936# VPWR 0.2061f
C12656 a_13364_31048# uio_oe[3] 0.00232f
C12657 _230_.I _252_.B 0.07976f
C12658 a_33028_27912# uo_out[6] 0.01624f
C12659 a_46404_15368# VPWR 0.20952f
C12660 a_25236_22020# a_25684_22020# 0.01328f
C12661 a_49852_15271# VPWR 0.34169f
C12662 _455_.D a_21600_26725# 0.09125f
C12663 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I _250_.C 0.12466f
C12664 a_43468_16839# a_43916_16839# 0.01288f
C12665 _417_.A2 _281_.A1 0.4483f
C12666 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I 0.04181f
C12667 a_31260_16839# VPWR 0.29679f
C12668 _404_.A1 a_44864_27165# 0.01911f
C12669 _313_.ZN a_36300_23544# 0.00123f
C12670 a_43268_1256# VPWR 0.20511f
C12671 a_21740_30951# a_21652_31048# 0.28563f
C12672 a_55588_1256# a_56036_1256# 0.01328f
C12673 a_34620_2727# a_35292_2727# 0.00544f
C12674 a_53460_24776# a_52852_24372# 0.13947f
C12675 a_55924_13800# a_56372_13800# 0.01328f
C12676 a_39236_17316# a_39212_16839# 0.00172f
C12677 _256_.A2 ui_in[1] 0.06064f
C12678 a_4604_17272# VPWR 0.33016f
C12679 _268_.A2 a_57220_29861# 0.15718f
C12680 vgaringosc.workerclkbuff_notouch_.I _393_.ZN 0.03015f
C12681 a_58388_10664# a_58500_9476# 0.02666f
C12682 a_52452_1636# VPWR 0.2085f
C12683 _355_.C a_30476_25112# 0.0237f
C12684 a_16252_1159# a_16164_1256# 0.28563f
C12685 _379_.Z a_18472_29076# 0.00757f
C12686 a_46268_12135# a_46180_12232# 0.28563f
C12687 a_13252_1636# a_12892_1592# 0.08707f
C12688 a_60604_27815# VPWR 0.31586f
C12689 a_66004_20072# a_66092_18407# 0.00151f
C12690 a_11460_29860# a_11908_29860# 0.01328f
C12691 a_53908_26724# a_54356_26724# 0.01328f
C12692 a_37892_17316# a_37980_17272# 0.28563f
C12693 a_33948_17272# a_34396_17272# 0.01288f
C12694 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN VPWR 0.48133f
C12695 a_47388_17272# a_47412_16936# 0.00172f
C12696 a_56708_1636# a_57156_1636# 0.01328f
C12697 a_67684_11044# a_67324_11000# 0.08707f
C12698 a_63740_11000# a_64188_11000# 0.01288f
C12699 a_23108_2824# VPWR 0.21435f
C12700 _455_.Q _455_.D 0.62709f
C12701 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I VPWR 0.70486f
C12702 a_40644_31048# uo_out[0] 0.01707f
C12703 a_1020_23111# a_1380_23208# 0.08717f
C12704 a_22300_23111# a_22748_23111# 0.01288f
C12705 a_4940_24679# a_5300_24776# 0.08674f
C12706 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I _245_.I1 0.08273f
C12707 _343_.A2 a_24100_29480# 0.02039f
C12708 a_6084_2824# a_6172_1159# 0.0027f
C12709 a_4604_14136# VPWR 0.33016f
C12710 a_1468_18407# a_1380_18504# 0.28563f
C12711 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I 0.64652f
C12712 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN a_59708_23111# 0.00121f
C12713 _474_.CLK _274_.A2 0.6735f
C12714 _402_.A1 _284_.A2 1.84393f
C12715 _448_.Q _330_.A2 0.01851f
C12716 a_27328_25227# a_27716_25641# 0.00393f
C12717 a_25643_25273# a_25928_25273# 0.00277f
C12718 _260_.A1 a_43814_21236# 0.03357f
C12719 a_61164_20408# vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN 0.00149f
C12720 a_58924_12135# VPWR 0.31389f
C12721 a_7876_29480# VPWR 0.20968f
C12722 a_35652_2824# a_36100_2824# 0.01328f
C12723 a_45060_31048# VPWR 0.20667f
C12724 a_63616_31128# ui_in[0] 0.43293f
C12725 vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN 0.73655f
C12726 a_35740_30951# _288_.ZN 0.00163f
C12727 a_21404_24679# VPWR 0.31394f
C12728 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_59620_23208# 0.00856f
C12729 _452_.Q _441_.B 0.00375f
C12730 _452_.CLK a_41099_26841# 0.02239f
C12731 a_2724_4392# VPWR 0.20782f
C12732 a_44812_16839# a_44836_15748# 0.0016f
C12733 _417_.A2 a_47271_21640# 0.003f
C12734 a_45396_28292# a_45036_28248# 0.08674f
C12735 a_35874_27937# VPWR 0.01105f
C12736 a_33948_15704# VPWR 0.30233f
C12737 a_2812_9432# a_3260_9432# 0.0131f
C12738 _474_.CLK a_55340_24679# 0.03545f
C12739 a_52452_14180# a_52540_14136# 0.28563f
C12740 _330_.A1 a_36060_19369# 0.0444f
C12741 a_62084_15368# a_61948_14136# 0.00154f
C12742 a_48508_14136# a_48956_14136# 0.01288f
C12743 a_22548_28292# a_22636_28248# 0.28563f
C12744 a_49404_18407# VPWR 0.33714f
C12745 a_53100_16839# VPWR 0.31389f
C12746 a_65668_1256# VPWR 0.23284f
C12747 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I a_65668_18884# 0.0022f
C12748 _325_.A2 a_41600_19376# 0.00318f
C12749 a_41432_17801# VPWR 0.19226f
C12750 a_58588_1592# VPWR 0.30503f
C12751 a_65780_10664# a_65668_9476# 0.02666f
C12752 a_27004_1159# a_27588_1256# 0.01675f
C12753 _358_.A3 a_31820_25112# 0.01535f
C12754 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN a_57604_14180# 0.0018f
C12755 a_54556_12568# a_54468_11044# 0.00151f
C12756 a_3172_12232# a_3620_12232# 0.01328f
C12757 a_57132_12135# a_57492_12232# 0.08707f
C12758 a_19748_1636# a_20196_1636# 0.01328f
C12759 a_40004_23233# VPWR 0.02193f
C12760 _452_.Q _328_.A2 0.00673f
C12761 a_5388_21543# VPWR 0.35526f
C12762 a_45620_17316# a_46404_17316# 0.00276f
C12763 a_4852_26344# a_4964_25156# 0.02666f
C12764 _474_.CLK a_56260_31048# 0.02517f
C12765 a_45508_2824# VPWR 0.20348f
C12766 a_61052_11000# a_61164_10567# 0.02634f
C12767 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN 0.02157f
C12768 a_21404_23111# a_21316_23208# 0.28563f
C12769 a_47948_23111# a_47860_23208# 0.28563f
C12770 a_16052_24776# a_16500_24776# 0.01328f
C12771 a_24988_24679# a_24900_24776# 0.28563f
C12772 _397_.A1 _412_.A1 0.75853f
C12773 a_48508_9432# VPWR 0.33981f
C12774 _424_.A2 clk 0.01063f
C12775 a_58836_14180# VPWR 0.19418f
C12776 a_61948_27815# a_62308_27912# 0.08674f
C12777 a_31620_18504# a_32068_18504# 0.01328f
C12778 _325_.A1 _325_.B 0.92049f
C12779 a_6084_31048# a_5948_29816# 0.00154f
C12780 a_42148_15748# a_42236_15704# 0.28563f
C12781 _330_.A1 a_36548_21640# 0.00357f
C12782 a_52788_12232# VPWR 0.20862f
C12783 _237_.A1 VPWR 0.80323f
C12784 a_58836_18884# a_58476_18840# 0.0869f
C12785 _402_.A1 a_39256_28292# 0.02652f
C12786 a_5052_20408# a_4940_19975# 0.02634f
C12787 a_59620_23208# vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I 0.0016f
C12788 a_25796_24776# VPWR 0.21584f
C12789 a_25100_30951# _340_.A2 0.01543f
C12790 a_51756_16839# a_51780_15748# 0.0016f
C12791 _447_.Q a_36636_21543# 0.02272f
C12792 a_31396_21640# a_31372_20408# 0.0016f
C12793 a_33188_21640# a_33076_20452# 0.02666f
C12794 a_7068_2727# a_7428_2824# 0.08717f
C12795 a_33948_19975# a_33860_20072# 0.28563f
C12796 a_47748_15748# VPWR 0.20595f
C12797 _452_.Q _300_.A2 0.00156f
C12798 _430_.ZN _301_.Z 0.00289f
C12799 _304_.B ui_in[7] 0.01645f
C12800 a_29788_30345# VPWR 0.39881f
C12801 _237_.A1 a_59332_29816# 0.05903f
C12802 _459_.CLK uo_out[1] 0.05356f
C12803 a_3260_14136# a_3260_13703# 0.05841f
C12804 a_56260_14180# a_55900_14136# 0.08717f
C12805 _459_.Q _358_.A3 0.72446f
C12806 _452_.CLK a_35652_26344# 0.01165f
C12807 _455_.Q _454_.D 0.06471f
C12808 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN a_63764_23588# 0.00471f
C12809 a_44571_26841# a_44856_26841# 0.00277f
C12810 a_62404_25156# vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN 0.00261f
C12811 a_45284_12612# a_45732_12612# 0.01328f
C12812 a_41099_26841# a_41116_26247# 0.00112f
C12813 a_67660_13703# a_67684_12612# 0.0016f
C12814 a_57020_2727# a_57468_2727# 0.0131f
C12815 _451_.Q hold2.I 0.02544f
C12816 _363_.Z a_35660_27508# 0.02593f
C12817 a_40668_26247# VPWR 0.29679f
C12818 _436_.B a_40973_24776# 0.03412f
C12819 a_38428_1159# a_38340_1256# 0.28563f
C12820 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN _258_.I 0.08097f
C12821 a_3172_9096# a_3172_7908# 0.05841f
C12822 a_932_20072# a_1380_20072# 0.01328f
C12823 a_68108_12135# a_68020_12232# 0.28563f
C12824 _294_.A2 uo_out[6] 0.18799f
C12825 a_4068_7528# a_4068_6340# 0.05841f
C12826 a_8636_1159# VPWR 0.33285f
C12827 a_8188_29816# uio_oe[6] 0.00453f
C12828 _436_.ZN a_40084_25156# 0.00589f
C12829 a_2276_21640# VPWR 0.20634f
C12830 _352_.A2 a_26580_23588# 0.02755f
C12831 _244_.Z a_61052_26247# 0.0064f
C12832 a_49988_17316# a_50076_17272# 0.28563f
C12833 a_60964_27912# VPWR 0.20815f
C12834 a_58028_10567# a_58476_10567# 0.01288f
C12835 a_47300_1636# a_47164_1159# 0.00168f
C12836 a_43356_1592# a_43356_1159# 0.05841f
C12837 a_65980_1592# a_66428_1592# 0.0131f
C12838 _340_.A2 a_25420_30345# 0.04221f
C12839 a_67908_2824# VPWR 0.21391f
C12840 a_4156_10567# a_4852_10664# 0.01227f
C12841 a_43916_29816# a_43232_29480# 0.00107f
C12842 _311_.A2 a_38628_25156# 0.02166f
C12843 a_31932_23111# a_32292_23208# 0.08707f
C12844 a_19972_23208# a_20420_23208# 0.01328f
C12845 a_61164_23111# VPWR 0.32628f
C12846 _452_.CLK a_36548_25156# 0.00398f
C12847 _337_.A3 a_27140_26724# 0.14927f
C12848 a_59484_9432# VPWR 0.31143f
C12849 a_4516_23588# VPWR 0.20862f
C12850 a_26556_21543# a_27004_21543# 0.01288f
C12851 a_66428_14136# VPWR 0.32136f
C12852 a_4516_6340# VPWR 0.20862f
C12853 a_5388_21543# a_5300_21640# 0.28563f
C12854 a_1916_3160# VPWR 0.297f
C12855 a_64548_2824# a_64548_1636# 0.05841f
C12856 a_2276_29480# a_2276_28292# 0.05841f
C12857 _327_.A2 _325_.B 0.09009f
C12858 _474_.CLK a_54356_25156# 0.06094f
C12859 a_33148_25641# VPWR 0.40163f
C12860 a_2364_11000# VPWR 0.30029f
C12861 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN 0.01312f
C12862 a_58052_2824# a_58500_2824# 0.01328f
C12863 a_50300_20408# VPWR 0.35348f
C12864 a_64860_19975# a_65220_20072# 0.08674f
C12865 _474_.CLK a_51756_18407# 0.00243f
C12866 a_67996_18840# a_67884_18407# 0.02634f
C12867 a_32964_18884# VPWR 0.20348f
C12868 a_52415_31220# VPWR 0.57393f
C12869 _359_.B a_34708_29860# 0.00169f
C12870 a_2812_26247# VPWR 0.30213f
C12871 a_18492_2727# a_18404_2824# 0.28563f
C12872 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62284_26680# 0.03107f
C12873 a_30724_26020# a_31932_26247# 0.00513f
C12874 _282_.ZN a_47636_25940# 0.20225f
C12875 _448_.Q _304_.A1 0.05643f
C12876 _355_.C a_20396_27815# 0.00641f
C12877 VPWR ui_in[7] 0.5946f
C12878 _251_.A1 vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN 0.00585f
C12879 _260_.A2 a_43814_21236# 0.00508f
C12880 _334_.A1 a_35728_29480# 0.01734f
C12881 a_53436_9432# a_53884_9432# 0.0131f
C12882 a_55588_9476# a_55228_9432# 0.08717f
C12883 a_63105_28293# vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN 0.00109f
C12884 _324_.C vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.13452f
C12885 a_64100_14180# a_64548_14180# 0.01328f
C12886 a_60268_14136# a_61052_14136# 0.00443f
C12887 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I 0.08504f
C12888 _230_.I a_63952_29480# 0.05f
C12889 _330_.A1 a_41188_18840# 0.06278f
C12890 _304_.B _451_.Q 0.48922f
C12891 a_24392_28248# _346_.A2 0.22177f
C12892 a_61076_13800# a_61052_12568# 0.0016f
C12893 _223_.I _362_.B 0.00104f
C12894 a_52452_12612# a_52092_12568# 0.08663f
C12895 _330_.A1 _444_.D 0.03109f
C12896 _424_.B1 _284_.A2 0.03353f
C12897 _424_.A1 a_54020_21640# 0.00622f
C12898 _411_.A2 a_47802_26724# 0.00931f
C12899 _362_.B _443_.D 0.00883f
C12900 a_21268_27912# a_21044_27508# 0.01342f
C12901 a_30812_1159# VPWR 0.32517f
C12902 _403_.ZN a_44961_27912# 0.07802f
C12903 a_49404_1159# a_49764_1256# 0.08717f
C12904 a_25884_1592# a_26332_1592# 0.01288f
C12905 a_29828_1636# a_29916_1592# 0.28563f
C12906 a_64884_12232# a_65332_12232# 0.01328f
C12907 _304_.A1 a_36764_22512# 0.00139f
C12908 a_37980_26247# _431_.A3 0.0038f
C12909 a_33188_21640# VPWR 0.20854f
C12910 _311_.A2 _302_.Z 0.00101f
C12911 a_31820_25112# a_31803_24831# 0.00112f
C12912 a_55116_10567# a_55028_10664# 0.28563f
C12913 a_15044_2824# a_15044_1636# 0.05841f
C12914 a_11236_2824# a_11100_1592# 0.00154f
C12915 a_1020_21976# VPWR 0.30073f
C12916 _402_.A1 a_40692_27912# 0.00267f
C12917 _230_.I vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN 0.17233f
C12918 _397_.A1 a_52304_26399# 0.00103f
C12919 a_45920_20523# _416_.ZN 0.00527f
C12920 a_55956_25940# a_56720_26344# 0.00399f
C12921 a_65756_8999# VPWR 0.31505f
C12922 a_22996_23588# VPWR 0.20595f
C12923 a_45088_29123# _393_.A1 0.00192f
C12924 a_15492_29480# a_15604_28292# 0.02666f
C12925 a_24988_21543# a_25348_21640# 0.08707f
C12926 a_10876_2727# VPWR 0.31831f
C12927 a_67548_5863# VPWR 0.32135f
C12928 a_2724_18884# a_3172_18884# 0.01328f
C12929 a_60716_13703# VPWR 0.33091f
C12930 _424_.A2 _416_.A3 0.0494f
C12931 _355_.C a_18028_28777# 0.01334f
C12932 _242_.Z VPWR 0.87331f
C12933 a_51868_15704# a_52316_15704# 0.01288f
C12934 a_55812_11044# VPWR 0.20595f
C12935 _256_.A2 _324_.C 3.18901f
C12936 _325_.A1 a_42811_19668# 0.00999f
C12937 _282_.ZN a_46156_25112# 0.00326f
C12938 a_26916_31048# _340_.A2 0.00798f
C12939 a_15244_26680# VPWR 0.30824f
C12940 a_63428_15748# a_63516_15704# 0.28563f
C12941 _265_.ZN a_41392_27165# 0.01734f
C12942 _323_.A3 a_38304_20072# 0.02435f
C12943 uo_out[1] uo_out[7] 0.00841f
C12944 a_63105_28293# VPWR 0.96468f
C12945 _336_.A1 _355_.B 0.67887f
C12946 _304_.B _384_.A3 0.03712f
C12947 _352_.ZN VPWR 1.10522f
C12948 a_29468_2727# a_29828_2824# 0.08717f
C12949 _284_.B _264_.B 0.03165f
C12950 a_48084_18884# a_48888_19243# 0.00302f
C12951 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I a_62060_20408# 0.00275f
C12952 a_21540_28292# VPWR 0.21433f
C12953 _260_.ZN _447_.Q 0.24508f
C12954 a_3620_23588# a_3708_23544# 0.28563f
C12955 a_3620_6340# a_3708_6296# 0.28563f
C12956 a_2724_7908# a_2812_7864# 0.28563f
C12957 _433_.ZN _304_.ZN 0.01019f
C12958 a_4516_4772# a_4604_4728# 0.28563f
C12959 a_18964_20452# a_18604_20408# 0.08717f
C12960 a_20308_20452# a_20756_20452# 0.01328f
C12961 _288_.ZN VPWR 0.90415f
C12962 _421_.B VPWR 0.50218f
C12963 a_55228_27815# a_55676_27815# 0.01222f
C12964 a_1916_30951# a_2276_31048# 0.08717f
C12965 a_37968_31048# _293_.A2 0.02497f
C12966 a_56572_23111# clk 0.00243f
C12967 a_4604_1592# VPWR 0.32824f
C12968 _451_.Q VPWR 3.03501f
C12969 a_55364_12612# a_55452_12568# 0.28563f
C12970 a_58948_12612# a_59396_12612# 0.01328f
C12971 _459_.Q a_31803_24831# 0.01431f
C12972 a_24652_30951# _459_.CLK 0.00154f
C12973 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I 0.0028f
C12974 _459_.CLK a_31484_26680# 0.00739f
C12975 _330_.A1 a_34715_22137# 0.00224f
C12976 a_25796_24776# a_25684_23588# 0.02666f
C12977 a_22660_24776# a_22636_23544# 0.0016f
C12978 a_60828_1159# a_60740_1256# 0.28563f
C12979 a_38759_24072# _441_.B 0.00293f
C12980 _243_.A1 a_58656_27912# 0.00652f
C12981 a_53212_1159# VPWR 0.3289f
C12982 a_32592_25227# a_32980_25641# 0.00393f
C12983 a_62172_18840# VPWR 0.30373f
C12984 _476_.Q _422_.ZN 0.43935f
C12985 a_33188_1636# a_32828_1592# 0.08707f
C12986 a_43132_27815# a_43492_27912# 0.0869f
C12987 _478_.D _384_.A1 0.51049f
C12988 a_41228_27815# _330_.A1 0.00839f
C12989 a_51892_10664# a_52340_10664# 0.01328f
C12990 a_65868_10567# a_66228_10664# 0.08717f
C12991 _244_.Z a_60516_26344# 0.04094f
C12992 a_20956_1159# a_21404_1159# 0.0131f
C12993 a_4852_24776# a_4940_23111# 0.00151f
C12994 a_23892_22020# VPWR 0.20595f
C12995 a_23556_21640# a_24004_21640# 0.01328f
C12996 a_32516_18884# a_32156_18840# 0.08717f
C12997 a_33276_2727# VPWR 0.31439f
C12998 _359_.B _296_.ZN 0.00259f
C12999 a_54580_13800# VPWR 0.20622f
C13000 a_50884_2824# a_50972_1159# 0.0027f
C13001 a_67324_15271# a_67772_15271# 0.012f
C13002 a_21292_30951# uio_out[6] 0.00722f
C13003 a_49952_26724# VPWR 0.00491f
C13004 a_10116_29860# VPWR 0.20944f
C13005 a_62396_11000# VPWR 0.31389f
C13006 a_1916_15271# a_1828_15368# 0.28563f
C13007 a_20620_21976# a_20508_21543# 0.02634f
C13008 a_20956_23111# VPWR 0.31389f
C13009 _437_.ZN a_37408_23208# 0.02692f
C13010 a_3260_15271# a_3708_15271# 0.0131f
C13011 _459_.CLK a_25792_30301# 0.0022f
C13012 _398_.C _279_.Z 1.36802f
C13013 _384_.A3 VPWR 3.15175f
C13014 _399_.ZN a_49405_22805# 0.00195f
C13015 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I _243_.A1 0.00679f
C13016 a_65308_17272# a_65220_15748# 0.00151f
C13017 vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I a_66676_20452# 0.00504f
C13018 a_62420_23208# a_62868_23208# 0.01328f
C13019 a_40892_2727# a_40804_2824# 0.28563f
C13020 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN 0.01519f
C13021 a_54780_18840# vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN 0.00335f
C13022 a_58388_18884# a_58252_18407# 0.00168f
C13023 a_62732_16839# a_63092_16936# 0.08717f
C13024 a_64412_9432# a_64860_9432# 0.0131f
C13025 a_66564_9476# a_66204_9432# 0.08717f
C13026 a_2276_25156# a_2364_25112# 0.28563f
C13027 a_14820_31048# uio_oe[1] 0.00726f
C13028 a_65756_7864# a_66204_7864# 0.0131f
C13029 a_67908_7908# a_67996_7864# 0.28563f
C13030 a_20980_23588# a_21428_23588# 0.01328f
C13031 a_17396_23588# a_17484_23544# 0.28563f
C13032 a_5052_7864# a_4940_7431# 0.02634f
C13033 a_21764_1256# a_22212_1256# 0.01328f
C13034 a_66652_6296# a_67100_6296# 0.0131f
C13035 a_67548_4728# a_67996_4728# 0.012f
C13036 a_65084_14136# a_64972_13703# 0.02634f
C13037 a_1020_2727# a_1468_2727# 0.0131f
C13038 a_51084_13703# a_51532_13703# 0.01288f
C13039 _359_.B a_41160_29083# 0.02598f
C13040 a_40132_26344# a_40580_26344# 0.01328f
C13041 a_12444_29383# a_12892_29383# 0.0131f
C13042 a_16252_30951# a_17284_31048# 0.0032f
C13043 a_16916_31048# a_16164_31048# 0.00639f
C13044 _416_.A2 a_48068_21236# 0.00997f
C13045 a_8627_30644# a_8636_29383# 0.00173f
C13046 a_18404_1636# VPWR 0.20839f
C13047 a_3708_30951# a_4156_30951# 0.0131f
C13048 a_67124_20452# a_66988_19975# 0.00168f
C13049 _250_.ZN a_61940_29076# 0.00195f
C13050 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I a_63316_20452# 0.00483f
C13051 a_53572_27912# a_52360_26355# 0.00103f
C13052 a_17508_29860# _467_.D 0.00153f
C13053 a_67796_18504# a_67884_16839# 0.00151f
C13054 a_61724_15271# a_61636_15368# 0.28563f
C13055 a_39548_1592# a_40132_1636# 0.01675f
C13056 a_5300_18504# VPWR 0.21406f
C13057 a_50212_11044# a_50300_11000# 0.28563f
C13058 a_46268_11000# a_46716_11000# 0.01288f
C13059 a_37332_16936# a_37780_16936# 0.01328f
C13060 a_34084_28776# a_37324_28776# 0.00576f
C13061 _437_.A1 _311_.A2 0.34962f
C13062 a_54444_24679# a_54892_24679# 0.01255f
C13063 _284_.B a_48560_26369# 0.01212f
C13064 a_1828_26724# a_2276_26724# 0.01328f
C13065 a_54824_22045# VPWR 1.10706f
C13066 _330_.ZN a_39324_17272# 0.00161f
C13067 _381_.Z _395_.A1 0.76764f
C13068 _371_.A3 a_31484_26680# 0.00668f
C13069 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN clk 0.00745f
C13070 _349_.A4 _373_.ZN 0.00573f
C13071 _416_.A1 a_41642_25156# 0.00192f
C13072 a_48508_30951# a_48956_30951# 0.0131f
C13073 hold2.I a_42161_24776# 0.52215f
C13074 a_4156_12568# VPWR 0.30552f
C13075 a_55676_2727# VPWR 0.31143f
C13076 a_63964_18407# a_63876_18504# 0.28563f
C13077 a_67796_16936# a_67772_15271# 0.00134f
C13078 a_4852_26344# a_5300_26344# 0.01328f
C13079 a_19164_26247# a_19524_26344# 0.08663f
C13080 a_1828_2824# a_2276_2824# 0.01328f
C13081 a_56460_10567# VPWR 0.34525f
C13082 a_37756_15271# a_38340_15368# 0.01675f
C13083 vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN 0.81938f
C13084 a_62396_2727# a_62532_1636# 0.00154f
C13085 a_27564_21976# a_27452_21543# 0.02634f
C13086 _436_.B a_40092_27209# 0.01472f
C13087 a_18628_23208# VPWR 0.23332f
C13088 _337_.A3 a_28891_25273# 0.0218f
C13089 _268_.A2 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.01067f
C13090 a_38523_27967# VPWR 0.36674f
C13091 _447_.Q _311_.Z 0.00461f
C13092 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I 0.94828f
C13093 a_1468_28248# a_1916_28248# 0.0131f
C13094 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN 0.00363f
C13095 a_4068_28292# a_3708_28248# 0.08717f
C13096 a_4516_22020# a_4604_21976# 0.28563f
C13097 _495_.I a_41160_29083# 0.46369f
C13098 a_38764_20408# _325_.A2 0.00347f
C13099 _301_.A1 _316_.A3 1.40951f
C13100 _345_.A2 VPWR 0.57877f
C13101 a_51868_2727# a_52228_2824# 0.08717f
C13102 a_67908_17316# a_67996_17272# 0.28563f
C13103 a_26746_26344# VPWR 0.01649f
C13104 a_47972_18504# a_48420_18504# 0.01328f
C13105 a_16052_25156# a_16140_25112# 0.28563f
C13106 a_19636_25156# a_20084_25156# 0.01328f
C13107 a_4964_18884# a_4940_18407# 0.00172f
C13108 a_61948_14136# a_61972_13800# 0.00172f
C13109 _276_.A2 _274_.A3 0.01067f
C13110 a_48060_13703# a_47972_13800# 0.28563f
C13111 a_31284_20452# a_31732_20452# 0.01328f
C13112 a_29356_20408# a_30028_20408# 0.00544f
C13113 a_16252_30951# uio_oe[1] 0.00493f
C13114 a_36188_26247# _444_.D 0.00453f
C13115 a_58063_30644# a_58687_31220# 0.10419f
C13116 a_35180_16839# a_35092_16936# 0.28563f
C13117 a_47524_22021# VPWR 0.60357f
C13118 a_62396_11000# a_62308_9476# 0.00151f
C13119 _373_.A2 _337_.A3 0.01184f
C13120 a_24540_1592# VPWR 0.33352f
C13121 a_65532_12568# a_65980_12568# 0.01288f
C13122 a_2724_1636# a_3172_1636# 0.01328f
C13123 a_22636_29383# a_23084_29383# 0.01255f
C13124 _304_.B a_40220_19975# 0.00193f
C13125 _430_.ZN _439_.ZN 0.02923f
C13126 _402_.A1 _419_.A4 0.05691f
C13127 _251_.A1 a_60940_28248# 0.00263f
C13128 a_55924_12232# a_56012_10567# 0.00151f
C13129 a_53572_11044# a_53212_11000# 0.08707f
C13130 a_46852_1636# a_46492_1592# 0.08707f
C13131 _330_.A1 a_36548_17316# 0.00457f
C13132 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I 0.00954f
C13133 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN 0.00998f
C13134 _371_.A1 a_27676_26680# 0.0018f
C13135 a_56684_23544# VPWR 0.31911f
C13136 _474_.CLK a_54356_26724# 0.02842f
C13137 _363_.Z _294_.ZN 0.29045f
C13138 a_48172_18840# a_48060_18407# 0.02634f
C13139 a_43356_1159# a_43804_1159# 0.0131f
C13140 a_54692_20452# a_55140_20452# 0.01328f
C13141 a_67684_21640# a_67884_19975# 0.00119f
C13142 a_2276_27912# a_2276_26724# 0.05841f
C13143 a_53412_29480# a_52756_29076# 0.02261f
C13144 _399_.ZN a_51332_24072# 0.10854f
C13145 _441_.A2 a_41216_23208# 0.00233f
C13146 _436_.ZN _441_.A3 0.06056f
C13147 a_18964_20452# VPWR 0.21483f
C13148 _459_.CLK _362_.ZN 0.02247f
C13149 a_56236_24679# a_56148_24776# 0.28563f
C13150 _441_.A2 _325_.A1 0.14039f
C13151 a_22100_31048# uio_out[6] 0.00112f
C13152 _304_.B a_42161_24776# 0.00127f
C13153 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I a_60212_25156# 0.6051f
C13154 _230_.I _243_.B2 0.52808f
C13155 a_57604_12612# VPWR 0.21273f
C13156 _359_.B a_29232_29931# 0.01392f
C13157 a_9084_2727# a_9220_1636# 0.00154f
C13158 a_10876_29383# a_10788_29480# 0.28563f
C13159 a_47300_15368# a_47748_15368# 0.01328f
C13160 vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN VPWR 0.73671f
C13161 a_15244_28248# a_15244_27815# 0.05841f
C13162 a_24864_29931# a_25252_30345# 0.00393f
C13163 a_50548_10664# VPWR 0.24134f
C13164 _304_.A1 a_42460_20452# 0.00316f
C13165 a_49180_15271# a_49092_15368# 0.28563f
C13166 a_1916_4295# a_2276_4392# 0.08717f
C13167 a_1020_5863# a_1380_5960# 0.08717f
C13168 _294_.A2 _460_.Q 0.36692f
C13169 _290_.ZN a_34084_28776# 0.02073f
C13170 _359_.B _335_.ZN 0.01955f
C13171 _260_.A2 a_43750_23544# 0.0116f
C13172 a_50748_15271# a_51196_15271# 0.0131f
C13173 a_65980_15271# VPWR 0.37796f
C13174 vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN 0.03163f
C13175 a_63292_2727# a_63204_2824# 0.28563f
C13176 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN 0.00292f
C13177 vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN 0.00147f
C13178 a_18292_22020# a_18380_21976# 0.28563f
C13179 a_1916_15271# VPWR 0.297f
C13180 a_32156_16839# a_32604_16839# 0.0131f
C13181 a_47612_30951# a_47524_31048# 0.28563f
C13182 _294_.ZN a_33812_29860# 0.00424f
C13183 a_28708_23208# a_28796_21543# 0.00151f
C13184 a_22548_25156# a_22636_25112# 0.28563f
C13185 a_64412_7864# VPWR 0.3038f
C13186 a_20420_1256# VPWR 0.20348f
C13187 a_28460_23544# a_28820_24072# 0.052f
C13188 a_44164_1256# a_44612_1256# 0.01328f
C13189 _325_.A2 a_37360_19325# 0.03402f
C13190 a_66204_4728# VPWR 0.31657f
C13191 _397_.A2 a_47802_26724# 0.00129f
C13192 a_58924_13703# a_59284_13800# 0.08707f
C13193 a_10876_29383# VPWR 0.33653f
C13194 a_55900_14136# a_55812_12612# 0.00151f
C13195 a_23196_2727# a_23868_2727# 0.00544f
C13196 _417_.Z a_49448_20072# 0.32258f
C13197 a_2364_30951# VPWR 0.31493f
C13198 _399_.A2 a_49013_22805# 0.00142f
C13199 a_45708_16839# a_46068_16936# 0.08707f
C13200 _330_.A1 a_44571_26841# 0.02405f
C13201 a_50996_10664# a_50884_9476# 0.02666f
C13202 a_49204_10664# a_49180_9432# 0.0016f
C13203 a_4828_1159# a_4740_1256# 0.28563f
C13204 a_35988_16936# VPWR 0.2061f
C13205 a_38204_1592# VPWR 0.3289f
C13206 a_40220_19975# VPWR 0.29679f
C13207 a_62844_12568# a_62956_12135# 0.02634f
C13208 _355_.C _349_.A4 0.23184f
C13209 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN 0.00287f
C13210 _230_.I a_59172_26724# 0.1049f
C13211 a_4516_29860# a_4604_29816# 0.28563f
C13212 _383_.A2 _395_.A1 0.00128f
C13213 _397_.A1 _381_.Z 0.08264f
C13214 a_30724_17316# a_31172_17316# 0.01328f
C13215 _304_.B a_50996_28292# 0.00413f
C13216 a_50660_11044# a_50636_10567# 0.00172f
C13217 a_46716_11000# a_46716_10567# 0.05841f
C13218 a_57044_17316# vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN 0.00172f
C13219 a_59932_11000# a_60380_11000# 0.012f
C13220 a_47164_30951# VPWR 0.31143f
C13221 _384_.A3 a_51240_23340# 0.55603f
C13222 a_49764_1636# a_49852_1592# 0.28563f
C13223 a_53348_1636# a_53796_1636# 0.01328f
C13224 _452_.CLK a_32180_20452# 0.00118f
C13225 _478_.D clk 0.05828f
C13226 a_61500_27815# a_61948_27815# 0.01222f
C13227 a_1916_23111# a_2364_23111# 0.0131f
C13228 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN a_52316_27815# 0.00403f
C13229 _459_.CLK a_16140_26247# 0.00816f
C13230 _270_.A2 _255_.ZN 0.01149f
C13231 a_49404_18407# a_49316_18504# 0.28563f
C13232 a_43268_2824# a_43268_1636# 0.05841f
C13233 a_51220_18504# a_51308_16839# 0.00151f
C13234 a_67212_20408# a_67012_18884# 0.00119f
C13235 a_46628_18504# VPWR 0.20897f
C13236 a_67908_18884# a_67548_18840# 0.08674f
C13237 a_18292_25156# VPWR 0.21366f
C13238 _474_.CLK vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN 0.01873f
C13239 a_2276_27912# a_2724_27912# 0.01328f
C13240 a_16588_27815# a_16948_27912# 0.08717f
C13241 _360_.ZN a_33148_25641# 0.00267f
C13242 a_42161_24776# VPWR 1.24496f
C13243 a_29940_20452# VPWR 0.22752f
C13244 _251_.A1 _246_.B2 0.94824f
C13245 a_64188_12568# VPWR 0.31479f
C13246 _402_.A1 a_40038_28720# 0.03943f
C13247 a_34160_20523# a_36016_20893# 0.02307f
C13248 _319_.ZN a_34716_20937# 0.2211f
C13249 a_24228_2824# a_24676_2824# 0.01328f
C13250 _229_.I _243_.A1 0.52187f
C13251 _355_.C _467_.D 0.69223f
C13252 _437_.A1 a_36660_23588# 0.00194f
C13253 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I VPWR 1.39532f
C13254 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_56388_25940# 0.00741f
C13255 _325_.B a_43284_18191# 0.00115f
C13256 a_66452_16936# VPWR 0.21187f
C13257 a_12916_31048# uio_oe[3] 0.01804f
C13258 a_32580_27912# uo_out[6] 0.01597f
C13259 a_45956_15368# VPWR 0.23027f
C13260 _300_.ZN _301_.Z 0.12141f
C13261 _436_.B _452_.Q 0.0014f
C13262 a_49180_15271# VPWR 0.32928f
C13263 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62148_29505# 0.0011f
C13264 a_45284_14180# a_45732_14180# 0.01328f
C13265 a_30812_16839# VPWR 0.30073f
C13266 a_21292_30951# a_21652_31048# 0.0869f
C13267 _397_.A4 _411_.A2 0.05089f
C13268 a_42820_1256# VPWR 0.25435f
C13269 a_1020_2727# a_932_2824# 0.28563f
C13270 a_2276_13800# a_2276_12612# 0.05841f
C13271 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I 0.0122f
C13272 a_53076_24776# a_52852_24372# 0.01342f
C13273 a_4156_17272# VPWR 0.30552f
C13274 _268_.A2 a_56596_29861# 0.15114f
C13275 a_15604_23208# a_15604_22020# 0.05841f
C13276 _355_.C a_30388_25156# 0.01959f
C13277 vgaringosc.workerclkbuff_notouch_.I a_45800_30345# 0.01984f
C13278 a_52004_1636# VPWR 0.2085f
C13279 a_15580_1159# a_16164_1256# 0.01675f
C13280 a_45820_12135# a_46180_12232# 0.08717f
C13281 a_8860_1592# a_9308_1592# 0.01288f
C13282 a_12804_1636# a_12892_1592# 0.28563f
C13283 a_8996_29480# a_9444_29480# 0.01328f
C13284 a_51196_12568# a_51108_11044# 0.00151f
C13285 a_59820_12135# a_60268_12135# 0.01288f
C13286 a_60156_27815# VPWR 0.31926f
C13287 _355_.ZN a_28012_24679# 0.05431f
C13288 _287_.A2 _459_.CLK 0.15759f
C13289 a_50996_28292# VPWR 0.13006f
C13290 a_37892_17316# a_37532_17272# 0.08663f
C13291 a_67236_11044# a_67324_11000# 0.28563f
C13292 a_45956_31048# a_46628_31048# 0.00347f
C13293 _362_.ZN uo_out[7] 0.0225f
C13294 a_53660_11000# a_53772_10567# 0.02634f
C13295 a_57604_11044# a_57580_10567# 0.00172f
C13296 a_53572_15368# a_53572_14180# 0.05841f
C13297 _459_.CLK a_16796_27209# 0.0554f
C13298 a_22660_2824# VPWR 0.20815f
C13299 a_29020_1592# a_29020_1159# 0.05841f
C13300 _455_.Q a_20844_26680# 0.01162f
C13301 a_62420_23208# a_62420_22020# 0.05841f
C13302 a_40196_31048# uo_out[0] 0.01747f
C13303 a_56148_24776# VPWR 0.20518f
C13304 _251_.A1 vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I 0.03005f
C13305 _448_.Q a_40004_22020# 0.00116f
C13306 a_1020_23111# a_932_23208# 0.28563f
C13307 a_4940_24679# a_4852_24776# 0.28563f
C13308 a_22300_24679# a_22748_24679# 0.01288f
C13309 a_65756_1159# a_66204_1159# 0.01255f
C13310 a_1828_7528# a_2276_7528# 0.01328f
C13311 _343_.A2 a_22996_29480# 0.00585f
C13312 _324_.C _395_.A1 1.28078f
C13313 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN a_59260_23111# 0.00655f
C13314 a_2724_5960# a_3172_5960# 0.01328f
C13315 a_3620_4392# a_4068_4392# 0.01328f
C13316 a_4156_14136# VPWR 0.30552f
C13317 hold2.Z hold1.Z 0.03847f
C13318 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I a_55228_28248# 0.00769f
C13319 _363_.Z a_33140_29860# 0.02317f
C13320 a_31708_18407# a_32156_18407# 0.0131f
C13321 a_35140_26680# a_35292_26247# 0.00161f
C13322 a_1020_18407# a_1380_18504# 0.08717f
C13323 _435_.ZN _434_.ZN 0.05451f
C13324 _441_.A3 _439_.ZN 0.06405f
C13325 _256_.A2 a_59796_29480# 0.00111f
C13326 _448_.Q a_38644_19368# 0.00274f
C13327 a_27328_25227# a_28891_25273# 0.41635f
C13328 a_7428_29480# VPWR 0.20348f
C13329 a_58476_12135# VPWR 0.32775f
C13330 a_34844_15704# a_35292_15704# 0.01288f
C13331 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I clk 0.00652f
C13332 _242_.Z a_57156_27912# 0.0022f
C13333 a_62532_30736# ui_in[0] 0.01344f
C13334 a_44612_31048# VPWR 0.20736f
C13335 a_20956_24679# VPWR 0.31389f
C13336 a_49988_15748# a_49852_15271# 0.00168f
C13337 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I VPWR 0.7389f
C13338 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_59172_23208# 0.00254f
C13339 _447_.Q a_39796_22504# 0.51589f
C13340 a_2276_4392# VPWR 0.20634f
C13341 _452_.CLK a_41392_27165# 0.02873f
C13342 a_44948_28292# a_45036_28248# 0.28563f
C13343 a_33500_15704# VPWR 0.30042f
C13344 _417_.A2 a_47047_21640# 0.00162f
C13345 _428_.Z _417_.A2 0.01151f
C13346 _316_.A3 a_37296_22020# 0.02791f
C13347 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I 0.02072f
C13348 a_34586_27912# VPWR 0.01579f
C13349 a_40464_27165# a_40092_27209# 0.10745f
C13350 a_4964_9476# a_5052_9432# 0.28563f
C13351 a_50860_18407# a_51308_18407# 0.0131f
C13352 a_28012_21976# a_28460_21976# 0.01288f
C13353 _330_.A1 a_36432_19325# 0.04831f
C13354 _474_.CLK a_54892_24679# 0.01323f
C13355 a_53996_16839# a_54444_16839# 0.01222f
C13356 a_48956_18407# VPWR 0.31587f
C13357 a_65444_15368# a_65444_14180# 0.05841f
C13358 a_52452_14180# a_52092_14136# 0.08663f
C13359 a_40040_17675# a_40804_15748# 0.00128f
C13360 a_21628_28248# a_22636_28248# 0.00323f
C13361 a_22548_28292# a_22996_28292# 0.01328f
C13362 a_52652_16839# VPWR 0.31389f
C13363 a_64996_1256# VPWR 0.21436f
C13364 _397_.A4 _399_.ZN 0.04045f
C13365 a_66564_1256# a_67012_1256# 0.01328f
C13366 _430_.ZN _303_.ZN 0.00276f
C13367 _383_.A2 _397_.A1 0.4727f
C13368 a_50548_13800# a_50660_12612# 0.02666f
C13369 a_66676_13800# a_67124_13800# 0.01328f
C13370 a_45596_2727# a_46044_2727# 0.0131f
C13371 a_46716_18407# a_46852_17316# 0.00154f
C13372 _475_.Q a_49828_22020# 0.00373f
C13373 a_48529_22460# a_48921_22020# 0.00762f
C13374 _325_.A2 a_42392_19243# 0.01495f
C13375 _319_.A2 VPWR 0.53838f
C13376 a_41536_17636# VPWR 0.40624f
C13377 a_22660_23208# a_22548_22020# 0.02666f
C13378 a_27004_1159# a_26916_1256# 0.28563f
C13379 a_63068_1592# a_63204_1256# 0.00168f
C13380 a_58140_1592# VPWR 0.33563f
C13381 a_57132_12135# a_57044_12232# 0.28563f
C13382 a_39178_23208# VPWR 0.01438f
C13383 a_14236_29816# a_14684_29816# 0.01288f
C13384 a_4940_21543# VPWR 0.31945f
C13385 _427_.B1 a_53300_23047# 0.00181f
C13386 _325_.B VPWR 0.52323f
C13387 a_45620_17316# a_45708_17272# 0.28563f
C13388 a_46716_10567# a_47164_10567# 0.0131f
C13389 a_45060_2824# VPWR 0.20348f
C13390 a_59484_1592# a_59932_1592# 0.01288f
C13391 _325_.A1 a_40580_20452# 0.00251f
C13392 a_32828_23111# a_33276_23111# 0.01288f
C13393 a_20956_23111# a_21316_23208# 0.08707f
C13394 a_24540_24679# a_24900_24776# 0.08707f
C13395 a_48060_9432# VPWR 0.31143f
C13396 a_15244_21543# a_15692_21543# 0.0131f
C13397 _287_.A2 _371_.A3 0.01166f
C13398 a_61948_27815# a_61860_27912# 0.28563f
C13399 _304_.B _402_.B 0.00342f
C13400 a_57604_14180# VPWR 0.21177f
C13401 _328_.A2 a_44484_19668# 0.00917f
C13402 a_52340_12232# VPWR 0.20595f
C13403 a_42148_15748# a_41788_15704# 0.08707f
C13404 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN 0.01248f
C13405 a_46628_2824# a_47076_2824# 0.01328f
C13406 a_4964_29860# a_4828_29383# 0.00168f
C13407 a_1020_29816# a_1020_29383# 0.05841f
C13408 _358_.A2 a_31348_25156# 0.00395f
C13409 a_58388_18884# a_58476_18840# 0.28563f
C13410 a_25348_24776# VPWR 0.20728f
C13411 clkbuf_1_0__f_clk.I clk 0.23599f
C13412 a_24652_30951# _340_.A2 0.0018f
C13413 _402_.A1 _381_.A2 0.81464f
C13414 a_43784_19369# _325_.ZN 0.02515f
C13415 a_7068_2727# a_6980_2824# 0.28563f
C13416 _447_.Q a_35816_21192# 0.40705f
C13417 a_47300_15748# VPWR 0.20595f
C13418 a_33500_19975# a_33860_20072# 0.08717f
C13419 a_34644_20072# a_34732_18407# 0.0027f
C13420 a_30160_30301# VPWR 0.18804f
C13421 _424_.ZN a_53100_18407# 0.00264f
C13422 _237_.A1 a_58116_30344# 0.01798f
C13423 _452_.CLK _304_.ZN 0.00199f
C13424 a_49540_9476# a_49988_9476# 0.01328f
C13425 a_21652_31048# a_22100_31048# 0.01328f
C13426 a_55812_14180# a_55900_14136# 0.28563f
C13427 a_59732_14180# a_60180_14180# 0.01328f
C13428 _452_.CLK a_35204_26344# 0.02076f
C13429 _459_.Q a_31484_26680# 0.00896f
C13430 a_21964_25112# a_21876_23588# 0.00151f
C13431 _455_.Q a_22064_27912# 0.01772f
C13432 _287_.A2 uo_out[7] 0.04286f
C13433 a_9756_1592# a_9892_1256# 0.00168f
C13434 a_57492_13800# a_57604_12612# 0.02666f
C13435 a_53684_13800# a_53660_12568# 0.0016f
C13436 _363_.Z a_35216_27533# 0.00175f
C13437 _245_.Z _244_.Z 0.12901f
C13438 a_932_24776# a_932_23588# 0.05841f
C13439 _441_.ZN _434_.ZN 0.01471f
C13440 _436_.ZN _300_.ZN 0.00612f
C13441 a_40220_26247# VPWR 0.31467f
C13442 _436_.B a_40357_24776# 0.10485f
C13443 a_7964_1159# VPWR 0.35728f
C13444 a_37980_1159# a_38340_1256# 0.08717f
C13445 a_51532_12135# a_51556_11044# 0.0016f
C13446 a_67660_12135# a_68020_12232# 0.08717f
C13447 a_53684_12232# a_54132_12232# 0.01328f
C13448 a_22524_1592# a_22972_1592# 0.01288f
C13449 _436_.ZN a_39860_25156# 0.01306f
C13450 a_59172_22020# vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I 0.00117f
C13451 a_4852_5960# a_4964_4772# 0.02666f
C13452 a_7740_29816# uio_oe[6] 0.00113f
C13453 _244_.Z a_60604_26247# 0.0239f
C13454 _352_.A2 a_26132_23588# 0.00313f
C13455 a_1828_21640# VPWR 0.20348f
C13456 _437_.A1 a_36860_23111# 0.00293f
C13457 a_60516_27912# VPWR 0.20789f
C13458 a_49988_17316# a_49628_17272# 0.08707f
C13459 _324_.C _397_.A1 0.25547f
C13460 _340_.A2 a_25792_30301# 0.06258f
C13461 _327_.A2 a_40580_20452# 0.00258f
C13462 a_4156_10567# a_4068_10664# 0.28563f
C13463 a_67460_2824# VPWR 0.20815f
C13464 _223_.I _359_.B 0.02993f
C13465 a_31932_23111# a_31844_23208# 0.28563f
C13466 _452_.CLK a_36100_25156# 0.00642f
C13467 _455_.Q a_27588_26724# 0.00136f
C13468 _337_.A3 a_25867_26841# 0.01295f
C13469 a_59036_9432# VPWR 0.31143f
C13470 a_4068_23588# VPWR 0.2157f
C13471 _402_.B VPWR 0.34348f
C13472 a_4940_21543# a_5300_21640# 0.08674f
C13473 a_4068_6340# VPWR 0.2157f
C13474 a_1468_3160# VPWR 0.29679f
C13475 a_65980_14136# VPWR 0.36289f
C13476 _474_.CLK a_53908_25156# 0.033f
C13477 a_14820_31048# a_14684_29816# 0.00154f
C13478 a_33520_25597# VPWR 0.19094f
C13479 a_48644_15748# a_49092_15748# 0.01328f
C13480 a_1916_11000# VPWR 0.297f
C13481 _334_.A1 _359_.ZN 0.01352f
C13482 a_11908_29860# a_11772_29383# 0.00168f
C13483 a_64860_19975# a_64772_20072# 0.28563f
C13484 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I a_65556_23588# 0.0159f
C13485 a_10004_31048# uio_oe[5] 0.00345f
C13486 _330_.A1 _439_.ZN 0.04097f
C13487 a_27884_25641# a_28228_25273# 0.00275f
C13488 a_41188_18840# _332_.Z 0.00129f
C13489 _252_.B _244_.Z 0.04222f
C13490 a_2364_26247# VPWR 0.30029f
C13491 a_52247_31220# VPWR 0.0043f
C13492 _427_.B2 a_52452_21236# 0.38122f
C13493 a_32516_18884# VPWR 0.20348f
C13494 _359_.B a_34260_29860# 0.00168f
C13495 a_18044_2727# a_18404_2824# 0.08717f
C13496 _355_.C a_19948_27815# 0.00623f
C13497 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_61836_26680# 0.00395f
C13498 _389_.ZN _381_.Z 0.08589f
C13499 _363_.Z _362_.B 0.12469f
C13500 a_55140_9476# a_55228_9432# 0.28563f
C13501 a_52764_17272# a_52676_15748# 0.00151f
C13502 a_26220_21976# a_26132_20452# 0.0027f
C13503 a_49852_14136# a_49740_13703# 0.02634f
C13504 _355_.ZN a_28372_23588# 0.00725f
C13505 a_3708_20408# a_4156_20408# 0.0131f
C13506 _474_.Q a_47776_20893# 0.00159f
C13507 _371_.A1 a_31964_28292# 0.00111f
C13508 _230_.I a_61940_29076# 0.03675f
C13509 a_57580_23544# vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN 0.00145f
C13510 _290_.ZN a_33776_29123# 0.06869f
C13511 _258_.ZN vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I 0.0376f
C13512 a_48060_12568# a_48508_12568# 0.01288f
C13513 a_52004_12612# a_52092_12568# 0.28563f
C13514 _424_.A1 a_53572_21640# 0.02961f
C13515 _248_.B1 a_63105_28293# 0.08067f
C13516 a_49404_1159# a_49316_1256# 0.28563f
C13517 a_18628_24776# a_18740_23588# 0.02666f
C13518 _454_.D a_22496_27967# 0.00159f
C13519 a_30364_1159# VPWR 0.29679f
C13520 a_58476_12135# a_58500_11044# 0.0016f
C13521 a_5300_9096# a_5388_7431# 0.0027f
C13522 a_48420_12232# a_48420_11044# 0.05841f
C13523 a_29828_1636# a_29468_1592# 0.08707f
C13524 a_32740_21640# VPWR 0.20692f
C13525 _474_.Q _395_.A3 0.53361f
C13526 _311_.A2 a_39172_22504# 0.00302f
C13527 _293_.A2 a_39884_27815# 0.00185f
C13528 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN a_66988_19975# 0.00149f
C13529 a_54668_10567# a_55028_10664# 0.08707f
C13530 a_9532_1159# a_9980_1159# 0.0131f
C13531 a_932_10664# a_1380_10664# 0.01328f
C13532 _325_.A2 a_43828_16936# 0.00466f
C13533 a_4964_22020# VPWR 0.21167f
C13534 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_63105_28293# 0.02613f
C13535 _330_.A1 _330_.ZN 0.69164f
C13536 a_30500_23208# a_30948_23208# 0.01328f
C13537 _402_.A1 a_39796_27912# 0.00546f
C13538 a_55956_25940# a_56368_26344# 0.00736f
C13539 a_22548_23588# VPWR 0.2267f
C13540 a_67100_5863# VPWR 0.29679f
C13541 a_65308_8999# VPWR 0.30378f
C13542 _223_.I a_32144_26724# 0.00142f
C13543 a_3172_21640# a_3620_21640# 0.01328f
C13544 a_60268_13703# VPWR 0.29679f
C13545 a_10428_2727# VPWR 0.31603f
C13546 a_24988_21543# a_24900_21640# 0.28563f
C13547 a_36548_21640# a_36016_20893# 0.03552f
C13548 _355_.C a_18400_28733# 0.0209f
C13549 a_61860_27912# a_62308_27912# 0.01328f
C13550 _392_.A2 _404_.A1 0.0055f
C13551 a_61388_15704# a_61276_15271# 0.02634f
C13552 a_4156_21976# a_4156_21543# 0.05841f
C13553 a_55364_11044# VPWR 0.20595f
C13554 a_14796_26680# VPWR 0.30073f
C13555 _421_.A1 _281_.ZN 0.14091f
C13556 a_26468_31048# _340_.A2 0.01661f
C13557 _282_.ZN a_46068_25156# 0.00521f
C13558 hold1.Z _448_.Q 0.05709f
C13559 a_63428_15748# a_63068_15704# 0.08717f
C13560 a_66116_15748# a_66564_15748# 0.01328f
C13561 _319_.ZN a_34732_19975# 0.07504f
C13562 a_62503_28293# VPWR 0.50384f
C13563 _388_.B uo_out[3] 0.06019f
C13564 clkbuf_1_0__f_clk.I _416_.A3 0.00327f
C13565 a_35204_26344# a_34448_25597# 0.0368f
C13566 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.00218f
C13567 a_24316_26247# VPWR 0.34058f
C13568 _373_.ZN a_25124_28776# 0.00331f
C13569 _304_.B a_52900_26724# 0.03724f
C13570 a_62060_23111# a_62508_23111# 0.0131f
C13571 a_29468_2727# a_29380_2824# 0.28563f
C13572 _439_.ZN _226_.ZN 0.26897f
C13573 _397_.A2 _397_.A4 0.09859f
C13574 _260_.ZN a_42161_24776# 0.08175f
C13575 a_19328_28733# VPWR 1.06626f
C13576 a_1020_23544# a_1468_23544# 0.0131f
C13577 a_3620_23588# a_3260_23544# 0.08717f
C13578 a_4516_7908# a_4964_7908# 0.01328f
C13579 a_2724_7908# a_2364_7864# 0.08717f
C13580 a_10340_1256# a_10788_1256# 0.01328f
C13581 a_60516_9476# a_60964_9476# 0.01328f
C13582 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN a_62196_23588# 0.00706f
C13583 a_1020_6296# a_1468_6296# 0.0131f
C13584 a_3620_6340# a_3260_6296# 0.08717f
C13585 a_67324_14136# a_67772_14136# 0.01288f
C13586 a_57244_14136# a_57132_13703# 0.02634f
C13587 a_1916_4728# a_2364_4728# 0.0131f
C13588 a_4516_4772# a_4156_4728# 0.08674f
C13589 a_2812_3160# a_3260_3160# 0.0131f
C13590 _474_.CLK _412_.ZN 0.13627f
C13591 a_67436_16839# a_67460_15748# 0.0016f
C13592 a_18516_20452# a_18604_20408# 0.28563f
C13593 a_6084_31048# a_6172_29383# 0.0027f
C13594 a_1020_29383# a_1468_29383# 0.0131f
C13595 a_1916_30951# a_1828_31048# 0.28563f
C13596 a_56124_23111# clk 0.00241f
C13597 a_4156_1592# VPWR 0.30551f
C13598 a_1916_12568# a_1916_12135# 0.05841f
C13599 _459_.Q a_30796_24463# 0.00534f
C13600 a_55364_12612# a_55004_12568# 0.08707f
C13601 a_57940_13800# a_58028_12135# 0.00151f
C13602 a_24196_31048# _459_.CLK 0.00494f
C13603 _424_.A2 _284_.A2 0.02633f
C13604 _330_.A1 a_35008_22461# 0.00722f
C13605 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_57020_23111# 0.00149f
C13606 _324_.B _475_.Q 0.5042f
C13607 a_55476_12232# a_55364_11044# 0.02666f
C13608 _476_.Q a_51108_21640# 0.00219f
C13609 _439_.ZN _300_.ZN 0.01819f
C13610 _437_.ZN _434_.ZN 0.03907f
C13611 a_52764_1159# VPWR 0.3289f
C13612 a_3260_11000# a_3708_11000# 0.0131f
C13613 a_38575_24072# _441_.B 0.00192f
C13614 a_60380_1159# a_60740_1256# 0.08717f
C13615 a_65420_12135# a_65444_11044# 0.0016f
C13616 a_52884_18884# VPWR 0.00419f
C13617 _459_.Q _362_.ZN 0.01296f
C13618 a_932_16936# a_1380_16936# 0.01328f
C13619 a_32740_1636# a_32828_1592# 0.28563f
C13620 a_36324_1636# a_36772_1636# 0.01328f
C13621 _346_.A2 a_23920_27555# 0.09002f
C13622 hold2.I _441_.A2 0.02681f
C13623 a_43132_27815# a_43044_27912# 0.28563f
C13624 a_56572_29383# vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.00273f
C13625 _424_.B1 _381_.A2 0.09901f
C13626 a_65868_10567# a_65780_10664# 0.28563f
C13627 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN 0.62315f
C13628 a_31172_18504# a_31172_17316# 0.05841f
C13629 a_63616_31128# _230_.I 0.00133f
C13630 a_23444_22020# VPWR 0.20595f
C13631 a_32068_18884# a_32156_18840# 0.28563f
C13632 a_32828_2727# VPWR 0.31143f
C13633 a_33860_18884# a_34308_18884# 0.01328f
C13634 a_54132_13800# VPWR 0.20622f
C13635 a_3708_26247# a_4156_26247# 0.0131f
C13636 _450_.D a_43400_18909# 0.00599f
C13637 a_20250_31048# uio_out[6] 0.00532f
C13638 a_54444_25112# a_54892_25112# 0.01255f
C13639 a_9668_29860# VPWR 0.20652f
C13640 a_61948_11000# VPWR 0.31389f
C13641 _417_.Z VPWR 0.67181f
C13642 a_1468_15271# a_1828_15368# 0.08717f
C13643 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN 0.73318f
C13644 a_20508_23111# VPWR 0.31389f
C13645 _444_.D a_38852_25156# 0.00199f
C13646 _383_.A2 _389_.ZN 0.0151f
C13647 _399_.ZN a_49013_22805# 0.00634f
C13648 a_52900_26724# VPWR 0.21724f
C13649 _416_.A1 _404_.A1 0.13437f
C13650 _362_.ZN _461_.D 0.09667f
C13651 _395_.A2 _395_.A3 0.20361f
C13652 vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I a_66228_20452# 0.02572f
C13653 a_40444_2727# a_40804_2824# 0.08717f
C13654 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN _267_.A1 0.68202f
C13655 vgaringosc.workerclkbuff_notouch_.I a_45088_29123# 0.00109f
C13656 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN a_57492_23588# 0.00769f
C13657 a_62732_16839# a_62644_16936# 0.28563f
C13658 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN 0.0209f
C13659 a_54780_18840# a_54892_18407# 0.02634f
C13660 a_17396_23588# a_17036_23544# 0.08707f
C13661 a_66116_9476# a_66204_9432# 0.28563f
C13662 a_67908_7908# a_67548_7864# 0.08663f
C13663 a_14372_31048# uio_oe[1] 0.00354f
C13664 a_4068_25156# a_4516_25156# 0.01328f
C13665 a_2276_25156# a_1916_25112# 0.08717f
C13666 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN VPWR 0.84762f
C13667 a_54108_14136# a_54132_13800# 0.00172f
C13668 a_23756_20408# a_24204_20408# 0.0131f
C13669 _452_.Q _433_.ZN 0.10828f
C13670 a_25460_20452# a_26132_20452# 0.00347f
C13671 _359_.B a_37584_29123# 0.017f
C13672 a_16252_30951# a_16164_31048# 0.28563f
C13673 a_66204_17272# a_66092_16839# 0.02634f
C13674 a_17956_1636# VPWR 0.2067f
C13675 a_56796_11000# a_56708_9476# 0.0027f
C13676 _362_.B a_35660_27508# 0.03878f
C13677 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I 0.00682f
C13678 a_61860_12612# a_62308_12612# 0.01328f
C13679 a_25884_27815# _351_.A2 0.00116f
C13680 a_63764_23208# vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I 0.00188f
C13681 a_48508_12568# a_48508_12135# 0.05841f
C13682 a_52452_12612# a_52428_12135# 0.00172f
C13683 a_17060_29860# _467_.D 0.00315f
C13684 _231_.ZN a_59172_23208# 0.00324f
C13685 a_5300_12232# a_5388_10567# 0.0027f
C13686 a_50212_11044# a_49852_11000# 0.08707f
C13687 a_61276_15271# a_61636_15368# 0.08717f
C13688 _304_.B _441_.A2 0.00522f
C13689 a_62420_12232# a_62308_11044# 0.02666f
C13690 _437_.A1 a_37532_25112# 0.0081f
C13691 a_4852_18504# VPWR 0.22733f
C13692 a_34084_28776# a_36828_28776# 0.00582f
C13693 _451_.Q a_39796_22504# 0.00241f
C13694 _284_.B a_48292_26369# 0.01859f
C13695 _327_.Z _328_.A2 0.42225f
C13696 _312_.ZN a_36084_23208# 0.01909f
C13697 a_62420_10664# a_62868_10664# 0.01328f
C13698 a_31932_1159# a_32380_1159# 0.0131f
C13699 a_24452_24776# a_24540_23111# 0.00151f
C13700 a_66540_18407# a_66564_17316# 0.0016f
C13701 a_28932_2824# a_28932_1636# 0.05841f
C13702 a_25124_2824# a_24988_1592# 0.00154f
C13703 _371_.A3 a_31031_27208# 0.00293f
C13704 _448_.Q _301_.A1 0.43934f
C13705 _330_.A1 _303_.ZN 0.01028f
C13706 a_14796_26680# a_14796_26247# 0.05841f
C13707 _276_.A2 a_51457_29861# 0.07616f
C13708 _395_.A3 a_50196_22805# 0.01448f
C13709 _448_.Q a_39236_20072# 0.00306f
C13710 _349_.A4 a_25962_29480# 0.00718f
C13711 _355_.C a_25124_28776# 0.05995f
C13712 _416_.A1 a_40468_25157# 0.01157f
C13713 a_7092_31048# uio_oe[7] 0.00345f
C13714 a_3708_12568# VPWR 0.33374f
C13715 a_55228_2727# VPWR 0.31143f
C13716 a_61860_2824# a_61948_1159# 0.0027f
C13717 _327_.A2 _331_.ZN 0.03959f
C13718 a_19164_26247# a_19076_26344# 0.28563f
C13719 a_63516_18407# a_63876_18504# 0.08717f
C13720 a_35876_15368# a_36324_15368# 0.01328f
C13721 a_56012_10567# VPWR 0.31547f
C13722 a_37756_15271# a_37668_15368# 0.28563f
C13723 a_33483_29535# a_33728_29167# 0.00232f
C13724 _436_.B a_40464_27165# 0.03628f
C13725 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I 0.018f
C13726 a_57468_16839# a_58252_16839# 0.00443f
C13727 a_17844_23208# VPWR 0.21215f
C13728 a_39324_15271# a_39772_15271# 0.0131f
C13729 a_37516_27599# VPWR 0.39937f
C13730 a_51240_19624# a_52024_20083# 0.02307f
C13731 a_3620_28292# a_3708_28248# 0.28563f
C13732 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.6546f
C13733 _301_.A1 a_36764_22512# 0.00271f
C13734 a_1916_21976# a_2364_21976# 0.0131f
C13735 a_4516_22020# a_4156_21976# 0.08674f
C13736 a_38316_20408# _325_.A2 0.0023f
C13737 a_51868_2727# a_51780_2824# 0.28563f
C13738 _284_.ZN hold2.I 0.62327f
C13739 a_52988_26680# _412_.ZN 0.00613f
C13740 a_67908_17316# a_67548_17272# 0.08674f
C13741 a_63516_17272# a_63964_17272# 0.0131f
C13742 _330_.A1 _397_.A4 0.08341f
C13743 a_23892_23588# a_24340_23588# 0.01328f
C13744 a_66652_8999# a_67100_8999# 0.0131f
C13745 vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN a_61636_18504# 0.00636f
C13746 a_16052_25156# a_15692_25112# 0.08707f
C13747 _459_.Q _287_.A2 1.91441f
C13748 a_32740_1256# a_33188_1256# 0.01328f
C13749 a_2364_18840# a_2364_18407# 0.05841f
C13750 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_60416_25156# 0.00612f
C13751 _402_.ZN _324_.B 0.02312f
C13752 a_47612_13703# a_47972_13800# 0.08717f
C13753 a_61612_13703# a_62060_13703# 0.01288f
C13754 _398_.C _412_.ZN 0.60364f
C13755 a_11772_2727# a_12444_2727# 0.00544f
C13756 a_52092_14136# a_52004_12612# 0.00151f
C13757 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN 0.08878f
C13758 a_15460_31048# uio_oe[1] 0.0965f
C13759 a_60604_27815# a_60740_26724# 0.00154f
C13760 a_58063_30644# a_58519_31220# 0.00165f
C13761 a_34732_16839# a_35092_16936# 0.08707f
C13762 _249_.A2 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN 0.0022f
C13763 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.02137f
C13764 a_46352_22021# VPWR 0.6939f
C13765 a_31620_1636# VPWR 0.2147f
C13766 a_4068_10664# a_4068_9476# 0.05841f
C13767 a_59396_12612# a_59372_12135# 0.00172f
C13768 a_55452_12568# a_55564_12135# 0.02634f
C13769 a_16252_30951# a_16916_31048# 0.00996f
C13770 a_1020_25112# a_1020_24679# 0.05841f
C13771 a_51791_30644# a_52639_30644# 0.00337f
C13772 a_66452_18504# a_66900_18504# 0.01328f
C13773 _441_.A2 VPWR 0.76286f
C13774 a_47860_16936# a_48308_16936# 0.01328f
C13775 a_14684_1592# a_14684_1159# 0.05841f
C13776 a_42460_1592# a_42908_1592# 0.01288f
C13777 a_46404_1636# a_46492_1592# 0.28563f
C13778 a_53124_11044# a_53212_11000# 0.28563f
C13779 a_56708_11044# a_57156_11044# 0.01328f
C13780 _362_.B a_36188_26680# 0.0165f
C13781 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62396_26247# 0.00316f
C13782 a_56236_23544# VPWR 0.31547f
C13783 _304_.A1 a_39760_23588# 0.00132f
C13784 a_18096_27165# a_19860_26724# 0.01233f
C13785 _474_.CLK a_53908_26724# 0.05115f
C13786 a_52964_29480# a_52756_29076# 0.01801f
C13787 a_58028_17272# a_58164_16936# 0.00168f
C13788 _424_.A2 a_52452_24072# 0.3802f
C13789 a_40416_18885# VPWR 0.59819f
C13790 a_12444_29816# uio_oe[3] 0.00188f
C13791 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN a_57044_23588# 0.00121f
C13792 a_1468_27815# a_1916_27815# 0.0131f
C13793 a_55788_24679# a_56148_24776# 0.08663f
C13794 a_18516_20452# VPWR 0.23295f
C13795 a_21652_31048# uio_out[6] 0.0022f
C13796 a_59652_25640# a_60212_25156# 0.3026f
C13797 a_57156_12612# VPWR 0.21061f
C13798 _268_.A2 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN 0.84072f
C13799 a_12804_2824# a_13252_2824# 0.01328f
C13800 _378_.ZN a_18096_27165# 0.00815f
C13801 a_10428_29383# a_10788_29480# 0.08717f
C13802 _226_.ZN _303_.ZN 0.02388f
C13803 _261_.ZN _452_.Q 0.11853f
C13804 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I 0.00204f
C13805 a_31708_15704# a_31708_15271# 0.05841f
C13806 a_35652_15748# a_35516_15271# 0.00168f
C13807 a_50100_10664# VPWR 0.21473f
C13808 a_48732_15271# a_49092_15368# 0.08717f
C13809 a_25772_21976# a_25796_21640# 0.00172f
C13810 a_56596_29861# a_56572_29383# 0.0013f
C13811 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN VPWR 0.95969f
C13812 _407_.A1 a_51048_26680# 0.00136f
C13813 a_1916_4295# a_1828_4392# 0.28563f
C13814 _260_.A2 a_43126_24119# 0.00277f
C13815 _284_.ZN _304_.B 1.65857f
C13816 a_65532_15271# VPWR 0.338f
C13817 a_17472_28363# _378_.ZN 0.28638f
C13818 a_62844_2727# a_63204_2824# 0.08717f
C13819 a_18292_22020# a_17932_21976# 0.08707f
C13820 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I 0.05733f
C13821 a_66340_15368# a_66788_15368# 0.01328f
C13822 a_1468_15271# VPWR 0.29679f
C13823 _436_.B a_41564_26247# 0.00349f
C13824 a_47164_30951# a_47524_31048# 0.08717f
C13825 clkbuf_1_0__f_clk.I _448_.Q 0.01019f
C13826 a_19972_1256# VPWR 0.2245f
C13827 _325_.A2 a_36060_19369# 0.01444f
C13828 _384_.ZN a_49828_22020# 0.0018f
C13829 a_65756_4728# VPWR 0.31505f
C13830 a_67908_7908# VPWR 0.2157f
C13831 a_22548_25156# a_22996_25156# 0.01328f
C13832 a_21964_25112# a_22636_25112# 0.00544f
C13833 _452_.CLK _328_.A2 0.00141f
C13834 _300_.ZN _303_.ZN 0.07999f
C13835 a_54804_16936# a_55004_15271# 0.00119f
C13836 a_10428_29383# VPWR 0.33392f
C13837 a_58924_13703# a_58836_13800# 0.28563f
C13838 a_44388_27912# a_44571_26841# 0.00123f
C13839 _330_.A1 a_44864_27165# 0.02426f
C13840 a_1916_30951# VPWR 0.31164f
C13841 a_45708_16839# a_45620_16936# 0.28563f
C13842 _427_.A2 _395_.A3 0.00233f
C13843 _474_.Q _427_.B1 0.00497f
C13844 _474_.CLK _427_.ZN 0.17452f
C13845 a_932_9476# a_1380_9476# 0.01328f
C13846 a_35540_16936# VPWR 0.2062f
C13847 a_37756_1592# VPWR 0.3289f
C13848 a_48508_12135# a_49292_12135# 0.00443f
C13849 a_66340_12612# a_66316_12135# 0.00172f
C13850 a_4156_1159# a_4740_1256# 0.01675f
C13851 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN VPWR 0.82124f
C13852 a_5500_1592# a_5948_1592# 0.01288f
C13853 a_39772_19975# VPWR 0.29679f
C13854 a_4516_29860# a_4156_29816# 0.08707f
C13855 _230_.I a_58052_26724# 0.00189f
C13856 a_17036_25112# a_17036_24679# 0.05841f
C13857 a_20980_25156# a_20956_24679# 0.00172f
C13858 a_46716_30951# VPWR 0.31605f
C13859 a_49764_1636# a_49404_1592# 0.08707f
C13860 a_66676_12232# a_66764_10567# 0.00151f
C13861 _433_.ZN a_40357_24776# 0.08615f
C13862 a_20672_30301# _346_.B 0.01517f
C13863 a_47836_15271# a_47972_14180# 0.00154f
C13864 _285_.Z uo_out[0] 0.0445f
C13865 a_1916_24679# a_2364_24679# 0.0131f
C13866 _416_.A1 a_46800_20937# 0.00142f
C13867 a_48956_18407# a_49316_18504# 0.08663f
C13868 a_54332_1159# a_54780_1159# 0.0131f
C13869 a_58276_25156# a_58364_25112# 0.28563f
C13870 a_63068_18840# a_63516_18840# 0.0131f
C13871 a_46180_18504# VPWR 0.20894f
C13872 a_67460_18884# a_67548_18840# 0.28563f
C13873 a_17844_25156# VPWR 0.20639f
C13874 a_29356_20408# VPWR 0.33981f
C13875 a_16588_27815# a_16500_27912# 0.28563f
C13876 _402_.A1 a_38584_28292# 0.35572f
C13877 a_63740_12568# VPWR 0.31389f
C13878 _319_.ZN a_35088_20893# 0.00766f
C13879 a_34160_20523# a_34716_20937# 0.8399f
C13880 a_31620_15748# a_32068_15748# 0.01328f
C13881 _251_.A1 a_57220_29861# 0.06703f
C13882 _371_.ZN _350_.A1 0.06344f
C13883 a_16240_26795# uio_out[7] 0.00151f
C13884 _355_.C a_17060_29480# 0.00403f
C13885 a_59652_25640# VPWR 0.5652f
C13886 _436_.B _433_.ZN 0.16305f
C13887 _316_.ZN _319_.A3 0.01319f
C13888 a_37420_16839# a_37444_15748# 0.0016f
C13889 _378_.I a_21540_28292# 0.00163f
C13890 _352_.A2 VPWR 2.81236f
C13891 a_45416_29885# _397_.A2 0.00131f
C13892 a_66004_16936# VPWR 0.26985f
C13893 a_32132_27912# uo_out[6] 0.00223f
C13894 a_45284_15368# VPWR 0.20968f
C13895 a_11460_31048# uio_oe[3] 0.00176f
C13896 _284_.ZN VPWR 4.53823f
C13897 _256_.A2 _249_.A2 0.06072f
C13898 a_24788_22020# a_25236_22020# 0.01328f
C13899 a_43020_16839# a_43468_16839# 0.01288f
C13900 a_48732_15271# VPWR 0.2987f
C13901 _436_.ZN _264_.B 0.00379f
C13902 _417_.A2 _476_.Q 0.20012f
C13903 a_5388_16839# VPWR 0.35526f
C13904 a_64100_27912# vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN 0.00147f
C13905 a_55140_1256# a_55588_1256# 0.01328f
C13906 a_21292_30951# a_21204_31048# 0.28563f
C13907 a_42148_1256# VPWR 0.21708f
C13908 a_34172_2727# a_34620_2727# 0.0131f
C13909 a_55476_13800# a_55924_13800# 0.01328f
C13910 _304_.B a_40580_20452# 0.00753f
C13911 a_3708_17272# VPWR 0.33374f
C13912 a_57940_10664# a_58052_9476# 0.02666f
C13913 a_15580_1159# a_15492_1256# 0.28563f
C13914 a_51556_1636# VPWR 0.2085f
C13915 a_45820_12135# a_45732_12232# 0.28563f
C13916 vgaringosc.workerclkbuff_notouch_.I a_48104_30219# 0.03249f
C13917 _379_.Z a_18264_29480# 0.31604f
C13918 a_12804_1636# a_12444_1592# 0.08707f
C13919 _249_.A2 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I 0.00385f
C13920 a_58911_30644# a_59955_30600# 0.01189f
C13921 a_27328_25227# a_28012_24679# 0.00107f
C13922 _355_.ZN a_27172_24328# 0.05441f
C13923 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN VPWR 0.70746f
C13924 a_52988_26680# a_53908_26724# 0.00795f
C13925 a_11012_29860# a_11460_29860# 0.01328f
C13926 a_62404_25156# clk 0.00205f
C13927 _416_.A1 _435_.A3 0.70971f
C13928 a_33500_17272# a_33948_17272# 0.01288f
C13929 a_37444_17316# a_37532_17272# 0.28563f
C13930 a_46940_17272# a_46964_16936# 0.00172f
C13931 a_22212_2824# VPWR 0.20815f
C13932 a_56260_1636# a_56708_1636# 0.01328f
C13933 a_63292_11000# a_63740_11000# 0.01288f
C13934 a_67236_11044# a_66876_11000# 0.08707f
C13935 _459_.CLK a_17168_27165# 0.05286f
C13936 _442_.ZN a_39968_26841# 0.00242f
C13937 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN 0.00635f
C13938 a_55700_24776# VPWR 0.20348f
C13939 vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I VPWR 0.73158f
C13940 _311_.A2 _312_.ZN 0.70047f
C13941 a_39748_31048# uo_out[0] 0.01953f
C13942 a_21852_23111# a_22300_23111# 0.01288f
C13943 a_4156_24679# a_4852_24776# 0.01227f
C13944 a_3708_14136# VPWR 0.33374f
C13945 a_23084_29383# a_22996_29480# 0.28563f
C13946 _343_.A2 a_22548_29480# 0.00208f
C13947 a_5636_2824# a_5724_1159# 0.0027f
C13948 _363_.Z a_32916_29860# 0.0031f
C13949 _451_.Q a_41476_24776# 0.00252f
C13950 a_1020_18407# a_932_18504# 0.28563f
C13951 _352_.A2 a_28903_24776# 0.07196f
C13952 _229_.I _250_.C 0.18629f
C13953 _448_.Q a_39268_18840# 0.00166f
C13954 a_27328_25227# a_29184_25597# 0.02307f
C13955 _355_.ZN a_27884_25641# 0.21547f
C13956 _447_.Q _304_.ZN 0.12902f
C13957 _274_.A2 ui_in[7] 0.00628f
C13958 _272_.A2 ui_in[4] 0.0683f
C13959 a_6980_29480# VPWR 0.20348f
C13960 a_58028_12135# VPWR 0.33765f
C13961 _346_.B a_21044_27508# 0.43165f
C13962 a_35204_2824# a_35652_2824# 0.01328f
C13963 _265_.ZN _436_.B 0.05952f
C13964 _223_.ZN a_31396_26724# 0.00367f
C13965 a_44164_31048# VPWR 0.20789f
C13966 a_61860_30736# ui_in[0] 0.00219f
C13967 a_30795_29977# _337_.ZN 0.00127f
C13968 a_20508_24679# VPWR 0.31389f
C13969 _327_.A2 a_45732_18504# 0.12066f
C13970 _255_.I _246_.B2 0.16482f
C13971 _452_.CLK a_40092_27209# 0.02359f
C13972 a_1828_4392# VPWR 0.20348f
C13973 a_44364_16839# a_44388_15748# 0.0016f
C13974 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN 0.01092f
C13975 a_25348_21640# a_25460_20452# 0.02666f
C13976 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN a_64188_27815# 0.00209f
C13977 a_33052_15704# VPWR 0.29736f
C13978 a_2364_9432# a_2812_9432# 0.0131f
C13979 a_4964_9476# a_4604_9432# 0.08674f
C13980 a_14004_31048# uio_oe[3] 0.00142f
C13981 _474_.CLK a_54444_24679# 0.00911f
C13982 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _411_.A2 0.01938f
C13983 _330_.A1 a_35504_18955# 0.05942f
C13984 _261_.ZN a_40357_24776# 0.02849f
C13985 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN 0.00338f
C13986 a_48060_14136# a_48508_14136# 0.01288f
C13987 a_48508_18407# VPWR 0.32807f
C13988 a_52004_14180# a_52092_14136# 0.28563f
C13989 a_61636_15368# a_61500_14136# 0.00154f
C13990 a_52204_16839# VPWR 0.31389f
C13991 a_64548_1256# VPWR 0.20655f
C13992 _384_.A1 a_54088_22895# 0.01307f
C13993 a_60268_13703# a_60292_12612# 0.0016f
C13994 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I _241_.I0 0.62032f
C13995 a_40580_20452# VPWR 0.21241f
C13996 _475_.Q a_49604_22020# 0.00577f
C13997 _325_.A2 a_41188_18840# 0.52489f
C13998 a_41048_17341# VPWR 1.14252f
C13999 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN a_67684_24776# 0.03377f
C14000 a_65332_10664# a_65220_9476# 0.02666f
C14001 a_57692_1592# VPWR 0.33799f
C14002 a_26556_1159# a_26916_1256# 0.08717f
C14003 _284_.A2 hold1.Z 0.00345f
C14004 a_56460_12135# a_57044_12232# 0.01675f
C14005 a_19300_1636# a_19748_1636# 0.01328f
C14006 a_54108_12568# a_54020_11044# 0.00151f
C14007 a_2724_12232# a_3172_12232# 0.01328f
C14008 a_4156_21543# VPWR 0.3269f
C14009 _452_.Q _327_.Z 0.42044f
C14010 a_45620_17316# a_45260_17272# 0.0869f
C14011 _412_.A1 clk 0.03298f
C14012 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.00392f
C14013 _474_.CLK _268_.A1 0.83055f
C14014 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN _250_.A2 0.00134f
C14015 a_62980_1636# a_63652_1636# 0.00347f
C14016 _436_.B _261_.ZN 0.00975f
C14017 _237_.A1 a_58340_29860# 0.00132f
C14018 a_44612_2824# VPWR 0.20348f
C14019 _294_.ZN _362_.B 0.00895f
C14020 a_20956_23111# a_20868_23208# 0.28563f
C14021 a_24540_24679# a_24452_24776# 0.28563f
C14022 a_15604_24776# a_16052_24776# 0.01328f
C14023 _319_.A3 a_37384_19624# 0.52345f
C14024 a_47612_9432# VPWR 0.31143f
C14025 a_61500_27815# a_61860_27912# 0.08674f
C14026 a_57156_14180# VPWR 0.21376f
C14027 a_31172_18504# a_31620_18504# 0.01328f
C14028 _284_.A2 a_45396_25156# 0.01347f
C14029 a_5636_31048# a_5500_29816# 0.00154f
C14030 _328_.A2 a_43668_19668# 0.04196f
C14031 a_51892_12232# VPWR 0.20595f
C14032 a_41700_15748# a_41788_15704# 0.28563f
C14033 a_45284_15748# a_45732_15748# 0.01328f
C14034 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I VPWR 0.83408f
C14035 _358_.A2 a_31124_25156# 0.01232f
C14036 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN a_65108_23588# 0.00107f
C14037 _459_.Q a_35008_27533# 0.02852f
C14038 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I 0.00745f
C14039 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN 0.09042f
C14040 a_49492_18840# a_49840_19001# 0.00277f
C14041 a_58388_18884# a_58028_18840# 0.0869f
C14042 a_24900_24776# VPWR 0.20622f
C14043 _304_.A1 a_33724_23111# 0.0172f
C14044 a_24196_31048# _340_.A2 0.00101f
C14045 a_55208_22505# _427_.ZN 0.01434f
C14046 a_32740_21640# a_32628_20452# 0.02666f
C14047 a_30948_21640# a_30924_20408# 0.0016f
C14048 a_51308_16839# a_51332_15748# 0.0016f
C14049 a_43888_19204# _325_.ZN 0.2926f
C14050 a_6620_2727# a_6980_2824# 0.08717f
C14051 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN 0.0091f
C14052 _294_.ZN a_32628_26725# 0.04654f
C14053 a_46852_15748# VPWR 0.20595f
C14054 a_33500_19975# a_33412_20072# 0.28563f
C14055 _424_.A2 _419_.A4 0.07589f
C14056 a_22996_29480# a_22996_28292# 0.05841f
C14057 _251_.A1 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.03997f
C14058 vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN 0.03727f
C14059 _241_.I0 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.68736f
C14060 _459_.Q a_31031_27208# 0.00754f
C14061 _424_.ZN VPWR 0.23295f
C14062 _274_.A1 a_52756_29076# 0.51431f
C14063 a_2812_14136# a_2812_13703# 0.05841f
C14064 a_55812_14180# a_55452_14136# 0.08717f
C14065 a_29716_31048# uo_out[7] 0.01025f
C14066 a_24304_26795# a_25867_26841# 0.41635f
C14067 a_56572_2727# a_57020_2727# 0.0131f
C14068 _384_.A1 _473_.Q 0.18121f
C14069 a_67212_13703# a_67236_12612# 0.0016f
C14070 _384_.ZN _324_.B 0.00467f
C14071 _223_.ZN VPWR 0.97374f
C14072 a_37556_23588# _437_.ZN 0.02403f
C14073 a_39772_26247# VPWR 0.32117f
C14074 a_7516_1159# VPWR 0.3289f
C14075 a_37980_1159# a_37892_1256# 0.28563f
C14076 a_2724_9096# a_2724_7908# 0.05841f
C14077 a_67660_12135# a_67572_12232# 0.28563f
C14078 a_3620_7528# a_3620_6340# 0.05841f
C14079 _334_.A1 _285_.Z 0.0939f
C14080 _363_.Z _359_.B 0.08982f
C14081 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I clk 0.04737f
C14082 _352_.A2 a_25684_23588# 0.00291f
C14083 a_1380_21640# VPWR 0.20348f
C14084 a_49540_17316# a_49628_17272# 0.28563f
C14085 a_53124_17316# a_53572_17316# 0.01328f
C14086 a_60068_27912# VPWR 0.15903f
C14087 a_3708_10567# a_4068_10664# 0.08717f
C14088 a_57580_10567# a_58028_10567# 0.01288f
C14089 _365_.ZN _459_.CLK 0.02999f
C14090 a_67012_2824# VPWR 0.20815f
C14091 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_56124_28248# 0.00166f
C14092 a_65532_1592# a_65980_1592# 0.0131f
C14093 a_42908_1592# a_42908_1159# 0.05841f
C14094 a_46852_1636# a_46716_1159# 0.00168f
C14095 _350_.A2 _371_.A1 2.16162f
C14096 a_19524_23208# a_19972_23208# 0.01328f
C14097 a_31484_23111# a_31844_23208# 0.08707f
C14098 _452_.CLK a_35652_25156# 0.02106f
C14099 a_3620_23588# VPWR 0.22347f
C14100 _337_.A3 a_26160_27165# 0.20796f
C14101 a_58588_9432# VPWR 0.31968f
C14102 a_64100_2824# a_64100_1636# 0.05841f
C14103 a_46356_24072# VPWR 0.81231f
C14104 a_25884_21543# a_26556_21543# 0.00544f
C14105 a_3620_6340# VPWR 0.22347f
C14106 a_4940_21543# a_4852_21640# 0.28563f
C14107 a_1020_3160# VPWR 0.30073f
C14108 a_59708_23111# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.00111f
C14109 a_1828_29480# a_1828_28292# 0.05841f
C14110 a_65532_14136# VPWR 0.32412f
C14111 a_39884_27815# _436_.B 0.06595f
C14112 _452_.CLK a_34308_18884# 0.00702f
C14113 a_1468_11000# VPWR 0.29679f
C14114 _260_.ZN _441_.A2 0.18006f
C14115 a_32592_25227# VPWR 1.11545f
C14116 a_8996_31048# uio_oe[5] 0.00409f
C14117 a_57380_2824# a_58052_2824# 0.00347f
C14118 vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN VPWR 0.75297f
C14119 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I a_65108_23588# 0.00347f
C14120 a_64412_19975# a_64772_20072# 0.08674f
C14121 _355_.B a_28796_23111# 0.00164f
C14122 a_67548_18840# a_67436_18407# 0.02634f
C14123 a_32068_18884# VPWR 0.20348f
C14124 _359_.B a_33812_29860# 0.0017f
C14125 a_1916_26247# VPWR 0.297f
C14126 a_18044_2727# a_17956_2824# 0.28563f
C14127 a_35723_20569# a_35504_18955# 0.00113f
C14128 _355_.C a_19500_27815# 0.00306f
C14129 _421_.A1 a_47636_25940# 0.00452f
C14130 _402_.A1 _400_.ZN 0.45357f
C14131 a_52988_9432# a_53436_9432# 0.0131f
C14132 a_55140_9476# a_54780_9432# 0.08717f
C14133 _427_.B1 _427_.A2 0.23479f
C14134 a_62503_28293# a_62844_27815# 0.0013f
C14135 _452_.CLK _452_.Q 0.08967f
C14136 a_63652_14180# a_64100_14180# 0.01328f
C14137 _371_.A1 a_31516_28292# 0.00309f
C14138 _355_.ZN a_27924_23588# 0.00441f
C14139 _230_.I a_59572_29076# 0.01025f
C14140 _228_.ZN ui_in[4] 0.04772f
C14141 _290_.ZN a_33483_29535# 0.01214f
C14142 _452_.CLK a_35044_21640# 0.00116f
C14143 a_64212_13800# a_64100_12612# 0.02666f
C14144 a_52004_12612# a_51644_12568# 0.08707f
C14145 _438_.ZN a_40244_21640# 0.214f
C14146 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I 0.00179f
C14147 _424_.A1 a_53108_21640# 0.00128f
C14148 _281_.ZN a_51620_19911# 0.00192f
C14149 _370_.B _352_.A2 0.16012f
C14150 a_29916_1159# VPWR 0.29679f
C14151 a_48956_1159# a_49316_1256# 0.08717f
C14152 a_64212_12232# a_64884_12232# 0.00347f
C14153 a_25436_1592# a_25884_1592# 0.01288f
C14154 a_29380_1636# a_29468_1592# 0.28563f
C14155 _304_.B vgaringosc.ro_inv4.inv_array_notouch_\[3\].I 0.78282f
C14156 _304_.A1 a_38576_22504# 0.0025f
C14157 a_32292_21640# VPWR 0.20692f
C14158 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I a_64412_19975# 0.02465f
C14159 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN 0.00157f
C14160 a_37980_26247# a_37892_26344# 0.28563f
C14161 _452_.Q a_40316_23233# 0.00171f
C14162 _311_.A2 a_38968_22504# 0.00414f
C14163 a_54668_10567# a_54580_10664# 0.28563f
C14164 a_5188_29480# a_5388_27815# 0.00119f
C14165 a_53796_1636# a_53660_1159# 0.00168f
C14166 a_49852_1592# a_49852_1159# 0.05841f
C14167 a_35816_21192# _319_.A2 0.00237f
C14168 a_10788_2824# a_10652_1592# 0.00154f
C14169 a_14596_2824# a_14596_1636# 0.05841f
C14170 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I 0.00998f
C14171 a_47544_20127# VPWR 0.00204f
C14172 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_62503_28293# 0.02723f
C14173 _330_.A1 a_37408_18504# 0.07293f
C14174 a_4516_22020# VPWR 0.20862f
C14175 a_34308_24776# a_34756_24776# 0.01328f
C14176 a_64860_8999# VPWR 0.30145f
C14177 a_15044_29480# a_15156_28292# 0.02666f
C14178 a_66652_5863# VPWR 0.29679f
C14179 a_24540_21543# a_24900_21640# 0.08707f
C14180 _334_.A1 a_37444_26724# 0.00171f
C14181 _351_.A2 _351_.ZN 0.17399f
C14182 a_21964_23544# VPWR 0.34385f
C14183 _416_.A1 _416_.A2 0.14555f
C14184 a_2276_18884# a_2724_18884# 0.01328f
C14185 a_9980_2727# VPWR 0.31446f
C14186 a_59820_13703# VPWR 0.29679f
C14187 _459_.CLK a_29856_29123# 0.02964f
C14188 a_51420_15704# a_51868_15704# 0.01288f
C14189 a_54916_11044# VPWR 0.20595f
C14190 a_18044_29816# _379_.Z 0.00639f
C14191 a_57580_23544# _231_.I 0.03525f
C14192 a_26020_31048# _340_.A2 0.02217f
C14193 a_15156_26724# VPWR 0.20551f
C14194 a_62279_28293# VPWR 0.00688f
C14195 a_62980_15748# a_63068_15704# 0.28563f
C14196 _230_.I _257_.B 0.04524f
C14197 _319_.ZN a_33948_19975# 0.00507f
C14198 a_23868_26247# VPWR 0.32237f
C14199 _336_.A2 _355_.B 0.40381f
C14200 a_29020_2727# a_29380_2824# 0.08717f
C14201 a_47636_18884# a_48084_18884# 0.01328f
C14202 _337_.A3 _351_.A2 0.01338f
C14203 a_3172_23588# a_3260_23544# 0.28563f
C14204 a_2276_7908# a_2364_7864# 0.28563f
C14205 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN a_61748_23588# 0.04674f
C14206 a_19035_28409# VPWR 0.55721f
C14207 a_4068_4772# a_4156_4728# 0.28563f
C14208 a_3172_6340# a_3260_6296# 0.28563f
C14209 _279_.Z _421_.B 0.01042f
C14210 a_49764_26724# _395_.A2 0.23131f
C14211 a_4964_3204# a_5052_3160# 0.28563f
C14212 a_17932_20408# a_18604_20408# 0.00544f
C14213 a_19860_20452# a_20308_20452# 0.01328f
C14214 _369_.ZN _336_.A1 0.00333f
C14215 a_1468_30951# a_1828_31048# 0.08717f
C14216 _258_.I vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I 0.01965f
C14217 a_18760_29032# a_18028_28777# 0.00619f
C14218 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN _256_.A2 0.0822f
C14219 a_66787_30600# vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I 0.0026f
C14220 a_3708_1592# VPWR 0.33374f
C14221 a_54916_12612# a_55004_12568# 0.28563f
C14222 a_58500_12612# a_58948_12612# 0.01328f
C14223 _459_.Q a_31168_24419# 0.0075f
C14224 _365_.ZN uo_out[7] 0.02996f
C14225 _359_.B uo_out[3] 0.05647f
C14226 a_23084_30951# _459_.CLK 0.00613f
C14227 a_46198_27060# _284_.A2 0.0071f
C14228 a_25348_24776# a_25236_23588# 0.02666f
C14229 a_47860_23208# _475_.Q 0.02453f
C14230 a_52316_1159# VPWR 0.3289f
C14231 _284_.ZN _260_.ZN 0.00139f
C14232 a_60380_1159# a_60292_1256# 0.28563f
C14233 _317_.A2 _316_.A3 0.4788f
C14234 a_32740_1636# a_32380_1592# 0.08707f
C14235 a_34448_25597# a_35652_25156# 0.00712f
C14236 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I VPWR 1.1897f
C14237 a_52436_18884# VPWR 0.00636f
C14238 _346_.A2 a_23627_27967# 0.0284f
C14239 _478_.D a_52452_24072# 0.01597f
C14240 a_42684_27815# a_43044_27912# 0.0869f
C14241 _331_.ZN VPWR 0.50189f
C14242 a_65420_10567# a_65780_10664# 0.08717f
C14243 a_51444_10664# a_51892_10664# 0.01328f
C14244 a_36524_18407# a_36548_17316# 0.0016f
C14245 a_20508_1159# a_20956_1159# 0.0131f
C14246 _284_.A2 clkbuf_1_0__f_clk.I 0.00558f
C14247 a_22996_22020# VPWR 0.20595f
C14248 _424_.B1 _427_.B2 0.12711f
C14249 a_62532_30736# _230_.I 0.17687f
C14250 _260_.A1 a_42796_23981# 0.00135f
C14251 _334_.A1 _371_.A1 0.69256f
C14252 a_23108_21640# a_23556_21640# 0.01328f
C14253 a_32068_18884# a_31708_18840# 0.08717f
C14254 a_50436_2824# a_50524_1159# 0.0027f
C14255 a_53684_13800# VPWR 0.20622f
C14256 a_32380_2727# VPWR 0.31143f
C14257 a_66876_15271# a_67324_15271# 0.01222f
C14258 VPWR uio_in[4] 0.00217f
C14259 a_9220_29860# VPWR 0.2085f
C14260 a_7964_29383# uio_oe[6] 0.00107f
C14261 a_61500_11000# VPWR 0.31389f
C14262 _431_.A3 _435_.A3 0.07827f
C14263 a_20172_21976# a_20060_21543# 0.02634f
C14264 a_1468_15271# a_1380_15368# 0.28563f
C14265 _359_.B _371_.A2 0.02931f
C14266 _444_.D a_38628_25156# 0.00694f
C14267 a_20060_23111# VPWR 0.31389f
C14268 a_2812_15271# a_3260_15271# 0.0131f
C14269 _384_.A3 _279_.Z 0.00152f
C14270 a_26720_30301# _337_.A3 0.00137f
C14271 a_42392_19243# a_42896_18504# 0.00388f
C14272 a_64860_17272# a_64772_15748# 0.00151f
C14273 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _397_.A2 0.00547f
C14274 a_61972_23208# a_62420_23208# 0.01328f
C14275 _435_.ZN _432_.ZN 0.02401f
C14276 a_60852_15748# vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I 0.07161f
C14277 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN a_60940_15704# 0.0019f
C14278 a_40444_2727# a_40356_2824# 0.28563f
C14279 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN a_57044_23588# 0.00678f
C14280 _355_.C _336_.A1 0.11942f
C14281 a_62284_16839# a_62644_16936# 0.08717f
C14282 a_21316_1256# a_21764_1256# 0.01328f
C14283 a_66116_9476# a_65756_9432# 0.08717f
C14284 a_16948_23588# a_17036_23544# 0.28563f
C14285 a_20532_23588# a_20980_23588# 0.01328f
C14286 a_67460_7908# a_67548_7864# 0.28563f
C14287 a_65308_7864# a_65756_7864# 0.0131f
C14288 _265_.ZN a_41564_26247# 0.01602f
C14289 VPWR uio_out[7] 1.29888f
C14290 a_1828_25156# a_1916_25112# 0.28563f
C14291 _495_.I uo_out[3] 0.01183f
C14292 a_66204_6296# a_66652_6296# 0.0131f
C14293 a_67100_4728# a_67548_4728# 0.0131f
C14294 a_58924_18840# VPWR 0.33768f
C14295 a_50636_13703# a_51084_13703# 0.01288f
C14296 _359_.B a_37291_29535# 0.01867f
C14297 a_25460_20452# a_25548_20408# 0.28563f
C14298 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN clk 0.40687f
C14299 a_15460_31048# a_16164_31048# 0.00391f
C14300 a_11772_29383# a_12444_29383# 0.00544f
C14301 _427_.A2 _422_.ZN 0.06126f
C14302 a_39684_26344# a_40132_26344# 0.01328f
C14303 _294_.A2 uo_out[2] 0.13082f
C14304 a_17508_1636# VPWR 0.20402f
C14305 a_66676_20452# a_66540_19975# 0.00168f
C14306 a_63316_23208# vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I 0.00214f
C14307 a_3260_30951# a_3708_30951# 0.0131f
C14308 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I 0.02298f
C14309 _470_.D hold2.I 0.00169f
C14310 a_16612_29860# _467_.D 0.00196f
C14311 _251_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.00765f
C14312 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I 0.61715f
C14313 a_45820_11000# a_46268_11000# 0.01288f
C14314 a_49764_11044# a_49852_11000# 0.28563f
C14315 a_61276_15271# a_61188_15368# 0.28563f
C14316 a_67348_18504# a_67436_16839# 0.00151f
C14317 a_4068_18504# VPWR 0.22146f
C14318 a_36884_16936# a_37332_16936# 0.01328f
C14319 a_39100_1592# a_39548_1592# 0.012f
C14320 _437_.A1 a_37084_25112# 0.00332f
C14321 _336_.A2 a_25643_25273# 0.00377f
C14322 a_34084_28776# a_36420_28776# 0.00589f
C14323 a_58063_30644# _255_.ZN 0.00284f
C14324 a_53996_24679# a_54444_24679# 0.01255f
C14325 a_40668_19975# _328_.A2 0.00308f
C14326 a_1380_26724# a_1828_26724# 0.01328f
C14327 a_29856_29123# uo_out[7] 0.0234f
C14328 _330_.ZN a_39236_17316# 0.00142f
C14329 _424_.A2 _381_.A2 0.01311f
C14330 _470_.Q _395_.A1 0.01064f
C14331 _274_.A3 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.00431f
C14332 _371_.A3 a_30847_27208# 0.00292f
C14333 _427_.ZN vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN 0.00872f
C14334 a_6084_31048# uio_oe[7] 0.00409f
C14335 _448_.Q a_38788_20072# 0.04882f
C14336 _370_.B _223_.ZN 0.43953f
C14337 a_35728_29480# a_37584_29123# 0.02307f
C14338 a_36656_29123# a_37291_29535# 0.02112f
C14339 a_48060_30951# a_48508_30951# 0.0131f
C14340 a_54780_2727# VPWR 0.31143f
C14341 _330_.A1 _452_.D 0.50748f
C14342 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I 0.62415f
C14343 a_3260_12568# VPWR 0.30487f
C14344 a_1380_2824# a_1828_2824# 0.01328f
C14345 a_63516_18407# a_63428_18504# 0.28563f
C14346 a_18716_26247# a_19076_26344# 0.08674f
C14347 a_67348_16936# a_67324_15271# 0.00134f
C14348 a_4068_26344# a_4852_26344# 0.00276f
C14349 _452_.CLK _436_.B 0.60048f
C14350 a_55564_10567# VPWR 0.31547f
C14351 a_56964_26724# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.01221f
C14352 a_27116_21976# a_27004_21543# 0.02634f
C14353 a_37308_15271# a_37668_15368# 0.08717f
C14354 a_17396_23208# VPWR 0.20348f
C14355 a_61948_2727# a_62084_1636# 0.00154f
C14356 _337_.A3 a_27884_25641# 0.00218f
C14357 _230_.I vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I 0.06188f
C14358 _268_.A2 a_53616_29480# 0.00355f
C14359 a_37888_27555# VPWR 0.18835f
C14360 _340_.A2 a_29716_31048# 0.00974f
C14361 vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I a_67908_22020# 0.07069f
C14362 a_3620_28292# a_3260_28248# 0.08717f
C14363 a_1020_28248# a_1468_28248# 0.0131f
C14364 a_51420_2727# a_51780_2824# 0.08717f
C14365 a_4068_22020# a_4156_21976# 0.28563f
C14366 _424_.B2 a_52436_18884# 0.002f
C14367 a_67460_17316# a_67548_17272# 0.28563f
C14368 a_37964_18191# a_37892_17316# 0.00175f
C14369 a_53704_23219# a_55116_22895# 0.00393f
C14370 a_47524_18504# a_47972_18504# 0.01328f
C14371 a_29804_30951# _287_.A2 0.00119f
C14372 _459_.Q a_29716_31048# 0.0018f
C14373 a_15604_25156# a_15692_25112# 0.28563f
C14374 a_19188_25156# a_19636_25156# 0.01328f
C14375 a_47612_13703# a_47524_13800# 0.28563f
C14376 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_60064_25156# 0.00199f
C14377 a_61500_14136# a_61524_13800# 0.00172f
C14378 a_30836_20452# a_31284_20452# 0.01328f
C14379 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I a_55228_20408# 0.00608f
C14380 a_14908_30951# uio_oe[1] 0.04244f
C14381 a_34732_16839# a_34644_16936# 0.28563f
C14382 _279_.Z a_47524_22021# 0.00443f
C14383 a_26108_30951# a_24864_29931# 0.00102f
C14384 _218_.ZN _427_.B2 0.00985f
C14385 a_61948_11000# a_61860_9476# 0.00151f
C14386 a_31172_1636# VPWR 0.20847f
C14387 a_65084_12568# a_65532_12568# 0.01288f
C14388 a_2276_1636# a_2724_1636# 0.01328f
C14389 a_22188_29383# a_22636_29383# 0.01255f
C14390 a_51791_30644# a_52415_31220# 0.10419f
C14391 _284_.B a_43600_25640# 0.00154f
C14392 _237_.A1 ui_in[2] 0.05982f
C14393 _304_.B _470_.D 0.03289f
C14394 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN 0.8201f
C14395 a_67772_24679# VPWR 0.33084f
C14396 _447_.Q _300_.A2 0.6984f
C14397 a_52540_11000# a_53212_11000# 0.00544f
C14398 a_51791_30644# ui_in[7] 0.00629f
C14399 a_4852_15368# a_4964_14180# 0.02666f
C14400 a_55476_12232# a_55564_10567# 0.00151f
C14401 a_46404_1636# a_46044_1592# 0.08707f
C14402 _362_.B a_32628_26725# 0.01027f
C14403 _459_.CLK a_30240_24776# 0.00972f
C14404 a_55788_23544# VPWR 0.32256f
C14405 _304_.A1 a_39536_23588# 0.00241f
C14406 a_47724_18840# a_47612_18407# 0.02634f
C14407 a_48888_19243# a_49404_18407# 0.00138f
C14408 _474_.CLK a_52988_26680# 0.00427f
C14409 a_42908_1159# a_43356_1159# 0.0131f
C14410 a_54244_20452# a_54692_20452# 0.01328f
C14411 a_1828_27912# a_1828_26724# 0.05841f
C14412 a_55228_15704# a_55364_15368# 0.00168f
C14413 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN a_61188_15368# 0.0037f
C14414 _441_.A2 a_39780_22805# 0.01717f
C14415 _275_.A2 uio_in[0] 0.02921f
C14416 _436_.ZN a_41564_24679# 0.00342f
C14417 _261_.ZN _433_.ZN 0.02641f
C14418 _424_.A2 a_51988_24072# 0.00233f
C14419 a_55788_24679# a_55700_24776# 0.28563f
C14420 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN a_56596_23588# 0.00135f
C14421 vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN 0.14823f
C14422 a_17932_20408# VPWR 0.34338f
C14423 a_21204_31048# uio_out[6] 0.00589f
C14424 _255_.ZN vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I 0.03541f
C14425 _474_.CLK _398_.C 0.0888f
C14426 _358_.A3 _358_.A2 0.5273f
C14427 a_56708_12612# VPWR 0.21151f
C14428 a_67348_16936# a_67796_16936# 0.01328f
C14429 a_8636_2727# a_8772_1636# 0.00154f
C14430 a_10428_29383# a_10340_29480# 0.28563f
C14431 _378_.ZN a_17803_26841# 0.00295f
C14432 a_46852_15368# a_47300_15368# 0.01328f
C14433 a_24864_29931# a_26427_29977# 0.41635f
C14434 a_58612_16936# vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN 0.00174f
C14435 a_14796_28248# a_14796_27815# 0.05841f
C14436 a_49652_10664# VPWR 0.21204f
C14437 a_48732_15271# a_48644_15368# 0.28563f
C14438 a_57492_23588# VPWR 0.21685f
C14439 a_1468_4295# a_1828_4392# 0.08717f
C14440 a_37444_26724# a_37532_26680# 0.28563f
C14441 _260_.A1 a_43380_20452# 0.00167f
C14442 _249_.A2 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN 0.0014f
C14443 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I 0.04607f
C14444 _260_.A2 a_42796_23981# 0.00667f
C14445 a_35616_24776# _304_.A1 0.00162f
C14446 a_50300_15271# a_50748_15271# 0.0131f
C14447 _252_.ZN _231_.ZN 0.26012f
C14448 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_58364_25112# 0.00144f
C14449 a_65084_15271# VPWR 0.33974f
C14450 a_21428_22020# a_21876_22020# 0.01328f
C14451 a_17844_22020# a_17932_21976# 0.28563f
C14452 _229_.I _258_.I 0.0044f
C14453 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN 0.0024f
C14454 a_1020_15271# VPWR 0.30073f
C14455 _421_.A1 _475_.Q 0.20321f
C14456 a_62844_2727# a_62756_2824# 0.28563f
C14457 a_47164_30951# a_47076_31048# 0.28563f
C14458 a_57132_17272# vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I 0.001f
C14459 a_31708_16839# a_32156_16839# 0.0131f
C14460 _436_.B a_41116_26247# 0.02793f
C14461 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I 0.00136f
C14462 a_40244_21640# a_40692_21640# 0.01328f
C14463 _384_.ZN a_49172_27508# 0.00115f
C14464 a_43716_1256# a_44164_1256# 0.01328f
C14465 a_67460_7908# VPWR 0.20348f
C14466 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN _324_.C 1.75827f
C14467 a_28012_23544# a_28460_23544# 0.01222f
C14468 a_19300_1256# VPWR 0.24258f
C14469 a_28260_23208# a_28348_21543# 0.00151f
C14470 _384_.ZN a_49604_22020# 0.00621f
C14471 a_65308_4728# VPWR 0.30378f
C14472 _325_.A2 a_36432_19325# 0.01357f
C14473 a_22748_2727# a_23196_2727# 0.0131f
C14474 a_4940_13703# a_4964_12612# 0.0016f
C14475 a_58476_13703# a_58836_13800# 0.08707f
C14476 a_9980_29383# VPWR 0.33235f
C14477 a_55452_14136# a_55364_12612# 0.00151f
C14478 a_4852_13800# a_5300_13800# 0.01328f
C14479 a_36060_19369# a_36076_18407# 0.0019f
C14480 _381_.Z clk 0.01791f
C14481 a_1468_30951# VPWR 0.31143f
C14482 _330_.A1 a_43564_27209# 0.00635f
C14483 a_45260_16839# a_45620_16936# 0.08707f
C14484 _417_.A2 a_53300_23047# 0.00107f
C14485 _324_.C _384_.A1 0.01273f
C14486 a_37308_1592# VPWR 0.3289f
C14487 a_4156_1159# a_4068_1256# 0.28563f
C14488 a_35092_16936# VPWR 0.23246f
C14489 a_50548_10664# a_50436_9476# 0.02666f
C14490 _474_.CLK a_55208_22505# 0.03933f
C14491 a_62396_12568# a_62508_12135# 0.02634f
C14492 _416_.A3 _473_.Q 0.2174f
C14493 _250_.A2 VPWR 0.20136f
C14494 a_39324_19975# VPWR 0.31495f
C14495 _470_.D VPWR 0.25796f
C14496 _397_.A1 _470_.Q 0.06628f
C14497 a_7652_29860# a_8100_29860# 0.01328f
C14498 a_4068_29860# a_4156_29816# 0.28563f
C14499 a_59484_11000# a_59932_11000# 0.01288f
C14500 a_50212_11044# a_50188_10567# 0.00172f
C14501 a_46268_11000# a_46268_10567# 0.05841f
C14502 a_46044_30951# VPWR 0.33981f
C14503 a_52900_1636# a_53348_1636# 0.01328f
C14504 a_49316_1636# a_49404_1592# 0.28563f
C14505 ui_in[4] ui_in[3] 0.03336f
C14506 _371_.ZN a_28112_27912# 0.00918f
C14507 a_61052_27815# a_61500_27815# 0.01255f
C14508 _416_.A1 a_46308_20937# 0.00103f
C14509 a_1468_23111# a_1916_23111# 0.0131f
C14510 a_48956_18407# a_48868_18504# 0.28563f
C14511 vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN 0.63963f
C14512 a_50772_18504# a_50860_16839# 0.00151f
C14513 a_42820_2824# a_42820_1636# 0.05841f
C14514 a_66764_20408# a_66564_18884# 0.00119f
C14515 a_67460_18884# a_67100_18840# 0.08674f
C14516 a_45732_18504# VPWR 0.1322f
C14517 a_58276_25156# a_57916_25112# 0.08674f
C14518 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I ui_in[1] 0.00416f
C14519 a_17396_25156# VPWR 0.20348f
C14520 a_28908_20408# VPWR 0.31143f
C14521 a_16140_27815# a_16500_27912# 0.08717f
C14522 a_1828_27912# a_2276_27912# 0.01328f
C14523 _360_.ZN a_32592_25227# 0.0066f
C14524 _437_.A1 _444_.D 0.17041f
C14525 a_63292_12568# VPWR 0.31389f
C14526 a_23780_2824# a_24228_2824# 0.01328f
C14527 a_34160_20523# a_35088_20893# 1.16391f
C14528 _251_.A1 a_56596_29861# 0.00417f
C14529 _474_.CLK _393_.A3 0.02807f
C14530 _378_.I a_19328_28733# 0.03747f
C14531 _447_.Q a_38325_22804# 0.00708f
C14532 a_17844_21640# a_17844_20452# 0.05841f
C14533 a_65332_16936# VPWR 0.21901f
C14534 a_45416_29885# a_46828_30345# 0.00393f
C14535 a_44836_15368# VPWR 0.20895f
C14536 _416_.A3 _475_.D 0.12373f
C14537 a_48284_15271# VPWR 0.29679f
C14538 _349_.A4 a_26468_27912# 0.0017f
C14539 _412_.B2 VPWR 0.53489f
C14540 a_4940_16839# VPWR 0.31945f
C14541 _359_.B a_34756_24776# 0.0011f
C14542 a_41700_1256# VPWR 0.20828f
C14543 a_67996_3160# a_67996_2727# 0.05841f
C14544 a_1828_13800# a_1828_12612# 0.05841f
C14545 _304_.B a_40132_20452# 0.00605f
C14546 _441_.ZN _260_.A1 0.00162f
C14547 a_3260_17272# VPWR 0.30487f
C14548 _416_.A1 a_46252_19759# 0.03717f
C14549 a_15156_23208# a_15156_22020# 0.05841f
C14550 a_15132_1159# a_15492_1256# 0.08717f
C14551 vgaringosc.workerclkbuff_notouch_.I a_45904_30180# 0.02463f
C14552 a_51108_1636# VPWR 0.20855f
C14553 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I VPWR 0.71567f
C14554 a_59372_12135# a_59820_12135# 0.01288f
C14555 a_45372_12135# a_45732_12232# 0.08717f
C14556 _379_.Z a_17786_29480# 0.00898f
C14557 a_50748_12568# a_50660_11044# 0.00151f
C14558 a_8548_29480# a_8996_29480# 0.01328f
C14559 a_12356_1636# a_12444_1592# 0.28563f
C14560 a_58252_18407# VPWR 0.3947f
C14561 a_37444_17316# a_37084_17272# 0.08707f
C14562 a_45508_31048# a_45956_31048# 0.01328f
C14563 a_57156_11044# a_57132_10567# 0.00172f
C14564 a_53212_11000# a_53324_10567# 0.02634f
C14565 a_28572_1592# a_28572_1159# 0.05841f
C14566 _459_.CLK a_16240_26795# 0.09976f
C14567 a_66788_11044# a_66876_11000# 0.28563f
C14568 a_21764_2824# VPWR 0.20815f
C14569 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I 0.00104f
C14570 _424_.A1 a_52408_19759# 0.03693f
C14571 _285_.Z _234_.ZN 0.00355f
C14572 a_55252_24776# VPWR 0.20348f
C14573 a_39300_31048# uo_out[0] 0.00408f
C14574 _448_.Q a_42168_22504# 0.06311f
C14575 a_21852_24679# a_22300_24679# 0.01288f
C14576 a_4156_24679# a_4068_24776# 0.28563f
C14577 _412_.ZN a_53548_24679# 0.00219f
C14578 _386_.A4 _400_.ZN 0.00326f
C14579 a_65084_1159# a_65756_1159# 0.00544f
C14580 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN a_56684_17272# 0.006f
C14581 a_1380_7528# a_1828_7528# 0.01328f
C14582 a_4940_19975# a_5388_19975# 0.01222f
C14583 a_3172_4392# a_3620_4392# 0.01328f
C14584 a_3260_14136# VPWR 0.30487f
C14585 a_49764_2824# a_49764_1636# 0.05841f
C14586 a_22636_29383# a_22996_29480# 0.0869f
C14587 a_2276_5960# a_2724_5960# 0.01328f
C14588 a_31260_18407# a_31708_18407# 0.0131f
C14589 _352_.A2 a_28679_24776# 0.00241f
C14590 _229_.I a_62148_29505# 0.00106f
C14591 _355_.ZN a_28256_25597# 0.0069f
C14592 a_27328_25227# a_27884_25641# 0.8399f
C14593 a_24636_25641# a_24980_25273# 0.00275f
C14594 a_57580_12135# VPWR 0.32122f
C14595 a_6532_29480# VPWR 0.20348f
C14596 a_34396_15704# a_34844_15704# 0.01288f
C14597 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I 0.62316f
C14598 _370_.ZN _371_.A1 0.00693f
C14599 a_43716_31048# VPWR 0.20654f
C14600 _287_.A1 _288_.ZN 2.10174f
C14601 vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN VPWR 0.71884f
C14602 _359_.B _294_.ZN 0.0375f
C14603 a_20060_24679# VPWR 0.31431f
C14604 _393_.ZN a_46837_29076# 0.00104f
C14605 a_60401_30300# _246_.B2 0.55152f
C14606 _274_.ZN _267_.ZN 0.00202f
C14607 _421_.A1 _402_.ZN 0.25645f
C14608 _397_.A2 _392_.A2 0.05149f
C14609 a_1380_4392# VPWR 0.20348f
C14610 _452_.CLK a_40464_27165# 0.01823f
C14611 _260_.A2 _435_.ZN 0.33478f
C14612 _301_.Z _302_.Z 0.00244f
C14613 a_32604_15704# VPWR 0.29679f
C14614 a_50412_18407# a_50860_18407# 0.0131f
C14615 a_4516_9476# a_4604_9432# 0.28563f
C14616 _359_.B a_29351_28293# 0.00557f
C14617 a_13452_30951# uio_oe[3] 0.00377f
C14618 a_27564_21976# a_28012_21976# 0.01288f
C14619 a_43736_25896# _284_.B 0.02613f
C14620 _474_.CLK a_53996_24679# 0.00698f
C14621 a_52004_14180# a_51644_14136# 0.08707f
C14622 a_64996_15368# a_64996_14180# 0.05841f
C14623 a_53548_16839# a_53996_16839# 0.01222f
C14624 a_48060_18407# VPWR 0.31435f
C14625 a_21628_28248# a_22548_28292# 0.00795f
C14626 a_49652_16936# a_49628_15704# 0.0016f
C14627 a_53460_16936# a_53572_15748# 0.02666f
C14628 a_51756_16839# VPWR 0.31389f
C14629 a_66116_1256# a_66564_1256# 0.01328f
C14630 a_64100_1256# VPWR 0.20363f
C14631 _384_.A1 a_54192_22851# 0.00205f
C14632 _248_.B1 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.71727f
C14633 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I clk 0.07422f
C14634 _416_.A3 a_47252_18884# 0.02258f
C14635 a_45148_2727# a_45596_2727# 0.0131f
C14636 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I a_56124_28248# 0.00311f
C14637 a_50100_13800# a_50212_12612# 0.02666f
C14638 a_66228_13800# a_66676_13800# 0.01328f
C14639 a_46268_18407# a_46404_17316# 0.00154f
C14640 a_56036_28292# _241_.I0 0.00424f
C14641 a_40132_20452# VPWR 0.20664f
C14642 a_57244_1592# VPWR 0.33431f
C14643 a_26556_1159# a_26468_1256# 0.28563f
C14644 a_62620_1592# a_62756_1256# 0.00168f
C14645 a_56460_12135# a_56372_12232# 0.28563f
C14646 a_47948_23111# VPWR 0.31517f
C14647 _397_.A1 a_52744_26031# 0.00272f
C14648 _474_.Q a_51108_21640# 0.03603f
C14649 a_13788_29816# a_14236_29816# 0.01288f
C14650 a_3708_21543# VPWR 0.33374f
C14651 a_45172_17316# a_45260_17272# 0.28563f
C14652 a_4068_26344# a_4068_25156# 0.05841f
C14653 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN 0.07317f
C14654 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.00999f
C14655 a_52639_30644# _268_.A1 0.00181f
C14656 a_44164_2824# VPWR 0.20348f
C14657 a_46268_10567# a_46716_10567# 0.0131f
C14658 a_62980_1636# a_63068_1592# 0.28563f
C14659 a_59036_1592# a_59484_1592# 0.01288f
C14660 _229_.I _255_.ZN 0.00155f
C14661 _237_.A1 a_61297_30300# 0.01432f
C14662 a_20508_23111# a_20868_23208# 0.08707f
C14663 a_32380_23111# a_32828_23111# 0.01288f
C14664 a_24092_24679# a_24452_24776# 0.08707f
C14665 _319_.A3 a_36836_20072# 0.00219f
C14666 a_47164_9432# VPWR 0.31143f
C14667 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I a_65756_27815# 0.00769f
C14668 a_61500_27815# a_61412_27912# 0.28563f
C14669 a_56708_14180# VPWR 0.20637f
C14670 a_14796_21543# a_15244_21543# 0.0131f
C14671 _293_.A2 _288_.ZN 0.02652f
C14672 a_48708_29816# a_49104_30345# 0.00232f
C14673 _284_.A2 a_44948_25156# 0.00653f
C14674 a_41700_15748# a_41340_15704# 0.08707f
C14675 _452_.Q _447_.Q 0.51002f
C14676 a_51444_12232# VPWR 0.20595f
C14677 a_45956_2824# a_46628_2824# 0.00347f
C14678 a_57940_18884# a_58028_18840# 0.28563f
C14679 a_57828_25156# clk 0.00546f
C14680 a_4156_20408# a_4156_19975# 0.05841f
C14681 a_24452_24776# VPWR 0.20622f
C14682 a_55312_22340# _427_.ZN 0.22847f
C14683 _294_.A2 _358_.A3 0.02322f
C14684 a_43400_18909# _325_.ZN 0.2968f
C14685 a_43888_19204# a_43784_19369# 0.10745f
C14686 _294_.ZN a_32144_26724# 0.02375f
C14687 a_6620_2727# a_6532_2824# 0.28563f
C14688 a_33052_19975# a_33412_20072# 0.08717f
C14689 a_46404_15748# VPWR 0.2267f
C14690 _384_.A1 _281_.A1 0.10307f
C14691 a_49092_9476# a_49540_9476# 0.01328f
C14692 _397_.A2 _416_.A1 0.11313f
C14693 _384_.A3 a_52036_22504# 0.00167f
C14694 a_56124_28248# vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.00564f
C14695 _241_.I0 a_56036_27912# 0.00828f
C14696 a_21204_31048# a_21652_31048# 0.01328f
C14697 a_4964_14180# a_4940_13703# 0.00172f
C14698 a_55364_14180# a_55452_14136# 0.28563f
C14699 a_59284_14180# a_59732_14180# 0.01328f
C14700 a_67884_19975# VPWR 0.34862f
C14701 _459_.Q a_30847_27208# 0.00832f
C14702 a_21516_25112# a_21428_23588# 0.00151f
C14703 _442_.ZN _311_.A2 0.00214f
C14704 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I a_61836_23544# 0.00303f
C14705 _351_.ZN a_24860_27209# 0.21984f
C14706 a_24304_26795# a_26160_27165# 0.02307f
C14707 a_43564_27209# a_43908_26841# 0.00275f
C14708 a_9308_1592# a_9444_1256# 0.00168f
C14709 a_53236_13800# a_53212_12568# 0.0016f
C14710 a_57044_13800# a_57156_12612# 0.02666f
C14711 a_37108_23588# _437_.ZN 0.0027f
C14712 _419_.A4 clkbuf_1_0__f_clk.I 0.04914f
C14713 _230_.I vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN 0.45015f
C14714 a_39324_26247# VPWR 0.32254f
C14715 _324_.C clk 0.02142f
C14716 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN VPWR 0.80029f
C14717 a_18096_27165# a_19188_25156# 0.0011f
C14718 a_37532_1159# a_37892_1256# 0.08717f
C14719 a_51084_12135# a_51108_11044# 0.0016f
C14720 a_53236_12232# a_53684_12232# 0.01328f
C14721 a_7068_1159# VPWR 0.3289f
C14722 a_67212_12135# a_67572_12232# 0.08717f
C14723 a_22076_1592# a_22524_1592# 0.01288f
C14724 a_932_3204# a_1380_3204# 0.01328f
C14725 a_932_21640# VPWR 0.22176f
C14726 a_49540_17316# a_49180_17272# 0.08707f
C14727 a_59172_27912# VPWR 0.63526f
C14728 _475_.Q a_49034_21640# 0.00137f
C14729 a_66564_2824# VPWR 0.21098f
C14730 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_55676_28248# 0.00665f
C14731 _304_.ZN _325_.B 0.00182f
C14732 a_67684_1636# a_67772_1592# 0.28563f
C14733 a_3708_10567# a_3620_10664# 0.28563f
C14734 _231_.ZN vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN 0.0103f
C14735 _350_.A2 a_30388_28776# 1.98589f
C14736 _443_.D a_37392_27967# 0.00159f
C14737 _441_.ZN _260_.A2 0.11611f
C14738 a_31484_23111# a_31396_23208# 0.28563f
C14739 _452_.CLK a_34155_25273# 0.00853f
C14740 _337_.A3 a_24860_27209# 0.00742f
C14741 a_59260_23111# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.00123f
C14742 _285_.Z a_39256_28292# 0.31509f
C14743 a_3172_23588# VPWR 0.20993f
C14744 a_58140_9432# VPWR 0.35372f
C14745 a_65084_14136# VPWR 0.32121f
C14746 a_3172_6340# VPWR 0.20993f
C14747 a_4156_21543# a_4852_21640# 0.01227f
C14748 a_4964_3204# VPWR 0.21167f
C14749 a_38816_27555# _436_.B 0.0029f
C14750 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN clk 0.09051f
C14751 a_14372_31048# a_14236_29816# 0.00154f
C14752 _452_.CLK a_33860_18884# 0.00362f
C14753 a_11460_29860# a_11324_29383# 0.00168f
C14754 a_48196_15748# a_48644_15748# 0.01328f
C14755 a_1020_11000# VPWR 0.30073f
C14756 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I a_64660_23588# 0.0017f
C14757 a_64412_19975# a_64324_20072# 0.28563f
C14758 _392_.A2 _330_.A1 0.00117f
C14759 _452_.CLK _433_.ZN 0.001f
C14760 a_31088_30301# a_30795_29977# 0.49319f
C14761 a_31620_18884# VPWR 0.20348f
C14762 a_1468_26247# VPWR 0.29679f
C14763 a_17596_2727# a_17956_2824# 0.08717f
C14764 _451_.Q _300_.A2 0.19119f
C14765 _432_.ZN a_41488_24072# 0.01198f
C14766 _474_.CLK vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN 0.04678f
C14767 a_54692_9476# a_54780_9432# 0.28563f
C14768 _389_.ZN _470_.Q 0.08844f
C14769 _417_.A2 _474_.D 0.01422f
C14770 a_62503_28293# a_62396_27815# 0.00101f
C14771 _398_.C a_53996_24679# 0.00176f
C14772 _408_.ZN _284_.A2 0.00165f
C14773 a_49404_14136# a_49292_13703# 0.02634f
C14774 _371_.A1 a_31068_28292# 0.00553f
C14775 a_3260_20408# a_3708_20408# 0.0131f
C14776 a_52316_17272# a_52228_15748# 0.00151f
C14777 _230_.I a_59348_29076# 0.00171f
C14778 _324_.C vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I 0.0341f
C14779 _452_.CLK a_34308_21640# 0.01364f
C14780 a_67548_2727# a_67996_2727# 0.01222f
C14781 a_47612_12568# a_48060_12568# 0.01288f
C14782 a_51556_12612# a_51644_12568# 0.28563f
C14783 _256_.A2 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN 0.02941f
C14784 a_22064_27912# a_23920_27555# 0.02307f
C14785 a_29468_1159# VPWR 0.29679f
C14786 a_58028_12135# a_58052_11044# 0.0016f
C14787 a_48956_1159# a_48868_1256# 0.28563f
C14788 a_47972_12232# a_47972_11044# 0.05841f
C14789 a_4852_9096# a_4940_7431# 0.00151f
C14790 a_67772_12568# a_67684_11044# 0.00151f
C14791 a_29380_1636# a_29020_1592# 0.08707f
C14792 _452_.Q a_41432_17801# 0.00254f
C14793 a_37532_26247# a_37892_26344# 0.08663f
C14794 a_31844_21640# VPWR 0.20692f
C14795 a_41116_26247# a_41564_26247# 0.01222f
C14796 _452_.Q a_40004_23233# 0.00291f
C14797 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_58948_26344# 0.00167f
C14798 _319_.A3 a_38228_20452# 0.00171f
C14799 a_31820_25112# a_30240_24776# 0.00516f
C14800 a_54220_10567# a_54580_10664# 0.08707f
C14801 a_60852_28292# a_60940_28248# 0.28563f
C14802 a_9084_1159# a_9532_1159# 0.0131f
C14803 a_46596_20127# VPWR 0.00246f
C14804 _330_.A1 a_36436_18504# 0.01037f
C14805 a_30052_23208# a_30500_23208# 0.01328f
C14806 _229_.I a_61836_26680# 0.00109f
C14807 _275_.A2 _274_.ZN 0.00152f
C14808 a_4068_22020# VPWR 0.2157f
C14809 a_58588_26247# a_59036_26247# 0.01222f
C14810 _351_.A2 a_24304_26795# 0.07718f
C14811 a_21516_23544# VPWR 0.31547f
C14812 a_64412_8999# VPWR 0.30566f
C14813 _334_.A1 a_36996_26724# 0.00167f
C14814 _303_.ZN _325_.A2 0.00136f
C14815 a_2724_21640# a_3172_21640# 0.01328f
C14816 a_59372_13703# VPWR 0.29679f
C14817 a_24540_21543# a_24452_21640# 0.28563f
C14818 a_9532_2727# VPWR 0.31143f
C14819 a_66204_5863# VPWR 0.31657f
C14820 a_51084_28248# _397_.A4 0.01737f
C14821 _459_.CLK a_29563_29535# 0.02066f
C14822 a_61412_27912# a_61860_27912# 0.01328f
C14823 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I a_56836_27208# 0.00117f
C14824 _324_.C _241_.Z 0.00239f
C14825 a_54468_11044# VPWR 0.20595f
C14826 _265_.ZN _452_.CLK 0.06289f
C14827 a_3708_21976# a_3708_21543# 0.05841f
C14828 a_25012_31048# _340_.A2 0.01259f
C14829 a_14708_26724# VPWR 0.22176f
C14830 _319_.ZN a_33500_19975# 0.00235f
C14831 a_65668_15748# a_66116_15748# 0.01328f
C14832 a_62980_15748# a_62620_15704# 0.08717f
C14833 vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN VPWR 0.72773f
C14834 _448_.Q _317_.A2 0.02153f
C14835 a_28036_26724# _355_.B 0.00355f
C14836 _319_.ZN a_35180_18407# 0.00144f
C14837 a_61612_23111# a_62060_23111# 0.0131f
C14838 a_23420_26247# VPWR 0.31863f
C14839 a_29020_2727# a_28932_2824# 0.28563f
C14840 _431_.A3 _430_.ZN 0.14382f
C14841 _416_.A1 _330_.A1 0.2255f
C14842 a_3172_23588# a_2812_23544# 0.08717f
C14843 _337_.A3 a_24900_27912# 0.01027f
C14844 a_16588_28248# VPWR 0.30535f
C14845 a_59932_9432# a_60516_9476# 0.01675f
C14846 a_14372_31048# a_14820_31048# 0.01328f
C14847 a_9892_1256# a_10340_1256# 0.01328f
C14848 a_3172_6340# a_2812_6296# 0.08717f
C14849 a_2276_7908# a_1916_7864# 0.08717f
C14850 a_4068_7908# a_4516_7908# 0.01328f
C14851 _251_.A1 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I 0.1539f
C14852 a_1468_4728# a_1916_4728# 0.0131f
C14853 a_4068_4772# a_3708_4728# 0.08717f
C14854 a_2364_3160# a_2812_3160# 0.0131f
C14855 a_4964_3204# a_4604_3160# 0.08674f
C14856 _412_.A1 _284_.A2 0.00928f
C14857 a_5636_31048# a_5724_29383# 0.0027f
C14858 a_66988_16839# a_67012_15748# 0.0016f
C14859 a_48529_22460# VPWR 0.48035f
C14860 a_66876_14136# a_67324_14136# 0.01288f
C14861 _311_.A2 _435_.ZN 0.00304f
C14862 _258_.I a_56484_29480# 0.0148f
C14863 _337_.A3 a_28596_26725# 0.002f
C14864 a_1468_30951# a_1380_31048# 0.28563f
C14865 a_3260_1592# VPWR 0.30486f
C14866 a_57492_13800# a_57580_12135# 0.00151f
C14867 a_54916_12612# a_54556_12568# 0.08707f
C14868 _324_.C hold2.Z 0.31381f
C14869 _395_.A1 a_50084_24328# 0.05733f
C14870 a_1468_12568# a_1468_12135# 0.05841f
C14871 _459_.Q a_30240_24776# 0.01153f
C14872 _459_.CLK a_21428_25156# 0.00649f
C14873 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I 0.0245f
C14874 _359_.B _388_.B 0.66268f
C14875 a_22636_30951# _459_.CLK 0.00253f
C14876 _459_.CLK a_31396_26724# 0.00176f
C14877 a_59932_1159# a_60292_1256# 0.08717f
C14878 a_36148_21976# _316_.A3 0.02813f
C14879 a_51868_1159# VPWR 0.3289f
C14880 a_64972_12135# a_64996_11044# 0.0016f
C14881 a_55028_12232# a_54916_11044# 0.02666f
C14882 a_34448_25597# a_34155_25273# 0.49241f
C14883 a_2812_11000# a_3260_11000# 0.0131f
C14884 a_35876_1636# a_36324_1636# 0.01328f
C14885 a_32292_1636# a_32380_1592# 0.28563f
C14886 _238_.I a_60940_28248# 0.00108f
C14887 a_50748_20408# a_51240_20452# 0.05364f
C14888 _346_.A2 a_22620_27599# 0.00784f
C14889 a_42684_27815# a_42596_27912# 0.28563f
C14890 _393_.ZN _397_.A1 0.1153f
C14891 a_37352_19001# VPWR 0.00204f
C14892 _285_.Z _296_.ZN 0.60753f
C14893 _452_.CLK _261_.ZN 0.00162f
C14894 a_65420_10567# a_65332_10664# 0.28563f
C14895 a_30724_18504# a_30724_17316# 0.05841f
C14896 a_61860_30736# _230_.I 0.30047f
C14897 _416_.A3 _416_.ZN 0.06519f
C14898 a_22548_22020# VPWR 0.2267f
C14899 _260_.A1 a_41488_24072# 0.31301f
C14900 _334_.A1 a_30388_28776# 0.01525f
C14901 a_31620_18884# a_31708_18840# 0.28563f
C14902 a_31932_2727# VPWR 0.31143f
C14903 _352_.ZN a_26548_24372# 0.38404f
C14904 a_52639_30644# _474_.CLK 0.01137f
C14905 a_53236_13800# VPWR 0.20622f
C14906 a_33412_18884# a_33860_18884# 0.01328f
C14907 a_3260_26247# a_3708_26247# 0.0131f
C14908 _349_.A4 _454_.Q 1.4108f
C14909 a_8772_29860# VPWR 0.2293f
C14910 a_53996_25112# a_54444_25112# 0.01255f
C14911 _304_.B _459_.CLK 0.22918f
C14912 a_61052_11000# VPWR 0.3185f
C14913 a_1020_15271# a_1380_15368# 0.08717f
C14914 a_19612_23111# VPWR 0.32678f
C14915 _304_.A1 _438_.ZN 0.00154f
C14916 _346_.ZN VPWR 0.24171f
C14917 _432_.ZN a_40880_23588# 0.00633f
C14918 _261_.ZN a_40316_23233# 0.00157f
C14919 _251_.A1 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.06133f
C14920 a_39996_2727# a_40356_2824# 0.08717f
C14921 vgaringosc.workerclkbuff_notouch_.I a_43788_29167# 0.00235f
C14922 a_54332_18840# a_54444_18407# 0.02634f
C14923 _371_.ZN _373_.ZN 0.13654f
C14924 a_62284_16839# a_62196_16936# 0.28563f
C14925 a_65668_9476# a_65756_9432# 0.28563f
C14926 _474_.Q _417_.A2 1.14825f
C14927 a_1828_25156# a_1468_25112# 0.08717f
C14928 a_67460_7908# a_67100_7864# 0.08717f
C14929 a_16948_23588# a_16588_23544# 0.08707f
C14930 a_4156_7864# a_4156_7431# 0.05841f
C14931 a_3620_25156# a_4068_25156# 0.01328f
C14932 _448_.Q _434_.ZN 0.0248f
C14933 a_40644_31048# uo_out[3] 0.00336f
C14934 a_58476_18840# VPWR 0.34238f
C14935 _388_.B _495_.I 0.86031f
C14936 a_65220_20072# a_65220_18884# 0.05841f
C14937 a_64188_14136# a_64300_13703# 0.02634f
C14938 a_53660_14136# a_53684_13800# 0.00172f
C14939 _359_.B a_36284_29167# 0.03912f
C14940 a_25460_20452# a_25100_20408# 0.08717f
C14941 a_23308_20408# a_23756_20408# 0.0131f
C14942 a_15460_31048# a_14820_31048# 0.00782f
C14943 a_14908_30951# a_16164_31048# 0.00231f
C14944 a_51196_21543# a_51108_21640# 0.28563f
C14945 a_52004_12612# a_51980_12135# 0.00172f
C14946 a_48060_12568# a_48060_12135# 0.05841f
C14947 a_61412_12612# a_61860_12612# 0.01328f
C14948 a_17060_1636# VPWR 0.20348f
C14949 a_22064_27912# a_22944_27599# 0.00306f
C14950 _332_.Z _452_.D 0.05228f
C14951 _386_.A4 a_47924_28292# 0.01988f
C14952 a_52228_27912# a_52360_26355# 0.00128f
C14953 _359_.B _362_.B 1.03674f
C14954 a_932_7908# VPWR 0.22176f
C14955 a_61972_12232# a_61860_11044# 0.02666f
C14956 a_49764_11044# a_49404_11000# 0.08707f
C14957 a_4852_12232# a_4940_10567# 0.00151f
C14958 a_3620_18504# VPWR 0.22347f
C14959 _437_.A1 a_36636_25112# 0.00119f
C14960 _336_.A2 a_25936_25597# 0.18009f
C14961 a_29563_29535# uo_out[7] 0.01133f
C14962 a_61972_10664# a_62420_10664# 0.01328f
C14963 a_67684_1636# a_67548_1159# 0.00168f
C14964 a_31484_1159# a_31932_1159# 0.0131f
C14965 _330_.ZN a_37980_17272# 0.01564f
C14966 _371_.A3 a_31396_26724# 0.19293f
C14967 _448_.Q a_36772_23208# 0.00184f
C14968 a_24004_24776# a_24092_23111# 0.00151f
C14969 a_66092_18407# a_66116_17316# 0.0016f
C14970 a_28484_2824# a_28484_1636# 0.05841f
C14971 a_24676_2824# a_24540_1592# 0.00154f
C14972 _383_.A2 a_49652_29480# 0.00309f
C14973 _424_.A2 _427_.B2 0.05631f
C14974 _448_.Q a_38304_20072# 0.00964f
C14975 _416_.A1 a_39860_25156# 0.01444f
C14976 _330_.A1 a_41776_18504# 0.01968f
C14977 a_33636_21640# a_34308_21640# 0.00347f
C14978 a_36656_29123# a_36284_29167# 0.10745f
C14979 a_35728_29480# a_37291_29535# 0.41635f
C14980 a_54332_2727# VPWR 0.31605f
C14981 a_58588_21543# vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I 0.00124f
C14982 a_2812_12568# VPWR 0.30213f
C14983 a_63068_18407# a_63428_18504# 0.08717f
C14984 a_18716_26247# a_18628_26344# 0.28563f
C14985 _381_.A2 clkbuf_1_0__f_clk.I 0.01156f
C14986 a_35428_15368# a_35876_15368# 0.01328f
C14987 _340_.A2 uio_out[2] 0.14967f
C14988 _246_.B2 _238_.I 0.49399f
C14989 a_59036_26247# _251_.ZN 0.03945f
C14990 _311_.A2 _441_.ZN 0.00185f
C14991 _459_.CLK VPWR 8.13118f
C14992 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I a_58028_20408# 0.00581f
C14993 a_55116_10567# VPWR 0.31547f
C14994 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I _231_.I 0.0015f
C14995 a_37308_15271# a_37220_15368# 0.28563f
C14996 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I 0.04837f
C14997 a_16948_23208# VPWR 0.20348f
C14998 _362_.B a_36656_29123# 0.00732f
C14999 _337_.A3 a_28256_25597# 0.00202f
C15000 _268_.A2 a_53412_29480# 0.00564f
C15001 _230_.I a_64324_29860# 0.00253f
C15002 a_51240_19624# a_51620_19911# 0.49319f
C15003 a_38876_15271# a_39324_15271# 0.0131f
C15004 a_3172_28292# a_3260_28248# 0.28563f
C15005 a_58364_25112# vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN 0.00448f
C15006 a_4068_22020# a_3708_21976# 0.08717f
C15007 a_1468_21976# a_1916_21976# 0.0131f
C15008 a_51420_2727# a_51332_2824# 0.28563f
C15009 _301_.A1 a_38576_22504# 0.05041f
C15010 a_63068_17272# a_63516_17272# 0.0131f
C15011 a_67460_17316# a_67100_17272# 0.08674f
C15012 a_66204_8999# a_66652_8999# 0.0131f
C15013 a_32292_1256# a_32740_1256# 0.01328f
C15014 a_15604_25156# a_15244_25112# 0.08707f
C15015 a_67100_7431# a_67548_7431# 0.0131f
C15016 a_23444_23588# a_23892_23588# 0.01328f
C15017 a_29804_30951# a_29716_31048# 0.28563f
C15018 a_1916_18840# a_1916_18407# 0.05841f
C15019 _324_.C a_45036_28248# 0.00912f
C15020 a_61164_13703# a_61612_13703# 0.01288f
C15021 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_59226_25156# 0.011f
C15022 a_51644_14136# a_51556_12612# 0.00151f
C15023 a_11324_2727# a_11772_2727# 0.0131f
C15024 a_47164_13703# a_47524_13800# 0.08717f
C15025 _384_.A3 _412_.ZN 0.02367f
C15026 a_55140_20452# a_55228_20408# 0.28563f
C15027 a_14460_30951# uio_oe[1] 0.00531f
C15028 _460_.D a_33024_25273# 0.00208f
C15029 a_25100_30951# _342_.ZN 0.00313f
C15030 a_24564_31048# _459_.CLK 0.00629f
C15031 a_33948_16839# a_34644_16936# 0.01227f
C15032 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN 0.00277f
C15033 a_65072_29860# vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.0025f
C15034 a_3620_10664# a_3620_9476# 0.05841f
C15035 a_30724_1636# VPWR 0.20348f
C15036 a_58948_12612# a_58924_12135# 0.00172f
C15037 a_55004_12568# a_55116_12135# 0.02634f
C15038 _424_.B1 a_52452_21236# 0.03131f
C15039 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN a_64772_26344# 0.07013f
C15040 _284_.B a_43192_25640# 0.00345f
C15041 a_15460_31048# a_16252_30951# 0.00279f
C15042 _431_.A3 _441_.A3 0.09003f
C15043 _451_.Q _452_.Q 2.57666f
C15044 a_51791_30644# a_52247_31220# 0.00165f
C15045 a_63092_26724# vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN 0.00561f
C15046 _388_.B _386_.ZN 0.00744f
C15047 a_66004_18504# a_66452_18504# 0.01328f
C15048 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I 0.76464f
C15049 a_56260_11044# a_56708_11044# 0.01328f
C15050 a_45956_1636# a_46044_1592# 0.28563f
C15051 a_42012_1592# a_42460_1592# 0.01288f
C15052 a_14236_1592# a_14236_1159# 0.05841f
C15053 a_47412_16936# a_47860_16936# 0.01328f
C15054 _250_.A2 a_62844_27815# 0.03007f
C15055 _352_.A2 _336_.Z 0.89523f
C15056 _459_.CLK a_28903_24776# 0.00191f
C15057 a_58164_18504# a_58252_16839# 0.0027f
C15058 a_55340_23544# VPWR 0.32732f
C15059 a_17803_26841# a_18096_27165# 0.58767f
C15060 a_48888_19243# a_48956_18407# 0.03137f
C15061 _260_.A1 a_40880_23588# 0.01447f
C15062 _395_.A2 _417_.A2 0.005f
C15063 _399_.ZN a_47636_23588# 0.00128f
C15064 a_17484_20408# VPWR 0.31184f
C15065 a_55340_24679# a_55700_24776# 0.08674f
C15066 a_1020_27815# a_1468_27815# 0.0131f
C15067 _400_.ZN _424_.A2 0.03511f
C15068 _248_.B1 _250_.A2 0.47752f
C15069 a_56260_12612# VPWR 0.20595f
C15070 a_12356_2824# a_12804_2824# 0.01328f
C15071 _355_.C _371_.ZN 0.13373f
C15072 a_9980_29383# a_10340_29480# 0.08717f
C15073 _342_.ZN a_25420_30345# 0.21523f
C15074 a_41440_28363# _265_.ZN 0.29556f
C15075 a_24864_29931# a_26720_30301# 0.02307f
C15076 a_35204_15748# a_35068_15271# 0.00168f
C15077 a_31260_15704# a_31260_15271# 0.05841f
C15078 a_49204_10664# VPWR 0.23151f
C15079 a_48284_15271# a_48644_15368# 0.08717f
C15080 a_25324_21976# a_25348_21640# 0.00172f
C15081 _324_.C a_49652_29480# 0.01669f
C15082 a_37444_26724# a_37084_26680# 0.0869f
C15083 a_1468_4295# a_1380_4392# 0.28563f
C15084 a_57044_23588# VPWR 0.21283f
C15085 _260_.A1 a_43156_20452# 0.00143f
C15086 _260_.A2 a_41488_24072# 0.01358f
C15087 _334_.A1 a_34292_28776# 0.00123f
C15088 a_37179_24831# a_37556_23588# 0.0306f
C15089 a_64412_15271# VPWR 0.32824f
C15090 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_57916_25112# 0.0165f
C15091 _252_.ZN a_58948_26344# 0.00432f
C15092 _247_.ZN _251_.ZN 0.0034f
C15093 _441_.B a_39178_23208# 0.007f
C15094 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN _250_.A2 0.23746f
C15095 a_62396_2727# a_62756_2824# 0.08717f
C15096 a_17844_22020# a_17484_21976# 0.08707f
C15097 _371_.A3 VPWR 1.2317f
C15098 a_67996_15704# VPWR 0.35098f
C15099 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I 0.09629f
C15100 vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN 0.02105f
C15101 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN a_65668_26344# 0.00755f
C15102 a_56684_17272# vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I 0.01189f
C15103 _436_.B a_40668_26247# 0.02981f
C15104 a_46716_30951# a_47076_31048# 0.08717f
C15105 a_65892_15368# a_66340_15368# 0.01328f
C15106 a_58836_17316# a_58700_16839# 0.00168f
C15107 _384_.ZN a_48988_27508# 0.00109f
C15108 a_21964_25112# a_22548_25156# 0.01675f
C15109 a_67012_7908# VPWR 0.20348f
C15110 _452_.CLK _327_.Z 0.0366f
C15111 a_18852_1256# VPWR 0.21061f
C15112 _325_.A2 a_35504_18955# 0.01652f
C15113 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN 0.01485f
C15114 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN 0.01997f
C15115 a_64860_4728# VPWR 0.30145f
C15116 a_58476_13703# a_58388_13800# 0.28563f
C15117 a_9532_29383# VPWR 0.32962f
C15118 a_54356_16936# a_54556_15271# 0.00119f
C15119 _460_.Q a_33188_25940# 0.33856f
C15120 a_1020_30951# VPWR 0.31538f
C15121 _330_.A1 a_43936_27165# 0.00795f
C15122 _275_.ZN _407_.A1 0.00128f
C15123 a_45260_16839# a_45172_16936# 0.28563f
C15124 _379_.A2 _379_.Z 0.31137f
C15125 a_3708_1159# a_4068_1256# 0.08717f
C15126 a_34644_16936# VPWR 0.24112f
C15127 _474_.CLK a_55312_22340# 0.08809f
C15128 _437_.A1 _439_.ZN 0.31128f
C15129 a_36860_1592# VPWR 0.3289f
C15130 a_44961_27912# VPWR 1.01094f
C15131 a_60940_28248# VPWR 0.33584f
C15132 a_5052_1592# a_5500_1592# 0.01288f
C15133 a_38876_19975# VPWR 0.31592f
C15134 a_65892_12612# a_65868_12135# 0.00172f
C15135 a_48060_12135# a_48508_12135# 0.0131f
C15136 a_20532_25156# a_20508_24679# 0.00172f
C15137 a_16588_25112# a_16588_24679# 0.05841f
C15138 _474_.D a_50644_21640# 0.01252f
C15139 a_4068_29860# a_3708_29816# 0.08707f
C15140 a_45596_30951# VPWR 0.31143f
C15141 _441_.A2 _304_.ZN 0.00168f
C15142 a_66228_12232# a_66316_10567# 0.00151f
C15143 a_49316_1636# a_48956_1592# 0.08707f
C15144 _238_.ZN _252_.B 0.11541f
C15145 a_47388_15271# a_47524_14180# 0.00154f
C15146 _371_.ZN a_27908_27912# 0.0018f
C15147 _346_.B _455_.Q 0.05809f
C15148 a_1468_24679# a_1916_24679# 0.0131f
C15149 a_53660_1159# a_54332_1159# 0.00544f
C15150 a_48508_18407# a_48868_18504# 0.08717f
C15151 a_40132_20072# a_40580_20072# 0.01328f
C15152 _328_.A2 _325_.B 0.05801f
C15153 VPWR uo_out[7] 0.78146f
C15154 a_57828_25156# a_57916_25112# 0.28563f
C15155 _416_.A1 a_38616_24328# 0.00465f
C15156 a_16948_25156# VPWR 0.20348f
C15157 a_67012_18884# a_67100_18840# 0.28563f
C15158 a_34980_22895# a_35188_22895# 0.00334f
C15159 a_44744_18559# VPWR 0.00204f
C15160 a_62620_18840# a_63068_18840# 0.0131f
C15161 a_16140_27815# a_16052_27912# 0.28563f
C15162 _294_.A2 uo_out[1] 0.02637f
C15163 a_28460_20408# VPWR 0.31143f
C15164 a_59226_25156# vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN 0.00206f
C15165 a_62844_12568# VPWR 0.31389f
C15166 a_31172_15748# a_31620_15748# 0.01328f
C15167 _311_.A2 _437_.ZN 0.24771f
C15168 _447_.Q a_38131_22804# 0.00786f
C15169 a_36972_16839# a_36996_15748# 0.0016f
C15170 _393_.A1 _392_.A2 0.0364f
C15171 _378_.I a_19035_28409# 0.07068f
C15172 _480_.Q VPWR 0.44345f
C15173 _304_.B _281_.ZN 0.0065f
C15174 a_45416_29885# a_46336_30345# 0.00306f
C15175 a_64884_16936# VPWR 0.21058f
C15176 a_44388_15368# VPWR 0.20348f
C15177 a_64188_27815# vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN 0.00354f
C15178 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN a_64884_26724# 0.07105f
C15179 _416_.A3 a_47271_21640# 0.03185f
C15180 a_58164_16936# vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN 0.0356f
C15181 a_24340_22020# a_24788_22020# 0.01328f
C15182 a_47836_15271# VPWR 0.29679f
C15183 a_42572_16839# a_43020_16839# 0.01288f
C15184 a_4156_16839# VPWR 0.3269f
C15185 a_50792_26344# VPWR 0.61021f
C15186 _303_.ZN _302_.Z 0.08462f
C15187 a_64660_23208# vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN 0.00429f
C15188 a_41252_1256# VPWR 0.20663f
C15189 a_54692_1256# a_55140_1256# 0.01328f
C15190 _393_.ZN _389_.ZN 0.1447f
C15191 a_55028_13800# a_55476_13800# 0.01328f
C15192 a_33724_2727# a_34172_2727# 0.0131f
C15193 vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN clk 0.08707f
C15194 _304_.B a_39684_20452# 0.0073f
C15195 a_37980_17272# a_37868_16839# 0.02634f
C15196 _474_.CLK a_57132_23544# 0.00166f
C15197 a_57492_10664# a_57604_9476# 0.02666f
C15198 a_2812_17272# VPWR 0.30213f
C15199 _416_.A1 a_46624_19715# 0.02629f
C15200 a_60212_25156# vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I 0.0021f
C15201 vgaringosc.workerclkbuff_notouch_.I a_45416_29885# 0.06361f
C15202 a_50660_1636# VPWR 0.23171f
C15203 a_58612_16936# VPWR 0.21827f
C15204 a_15132_1159# a_15044_1256# 0.28563f
C15205 a_45372_12135# a_45284_12232# 0.28563f
C15206 a_12356_1636# a_11996_1592# 0.08707f
C15207 VPWR uio_in[0] 0.33416f
C15208 a_58687_31220# a_58911_30644# 0.53809f
C15209 a_57580_18407# VPWR 0.33273f
C15210 a_10564_29860# a_11012_29860# 0.01328f
C15211 a_36996_17316# a_37084_17272# 0.28563f
C15212 a_33052_17272# a_33500_17272# 0.01288f
C15213 a_66788_11044# a_66428_11000# 0.08707f
C15214 a_62844_11000# a_63292_11000# 0.01288f
C15215 a_46492_17272# a_46516_16936# 0.00172f
C15216 _330_.A1 _431_.A3 0.2728f
C15217 _424_.A1 a_52512_19715# 0.0326f
C15218 a_21316_2824# VPWR 0.20815f
C15219 a_55812_1636# a_56260_1636# 0.01328f
C15220 _285_.Z a_40038_28720# 0.00467f
C15221 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN 0.06365f
C15222 a_54804_24776# VPWR 0.20348f
C15223 a_21404_23111# a_21852_23111# 0.01288f
C15224 a_3708_24679# a_4068_24776# 0.08717f
C15225 a_5188_2824# a_5276_1159# 0.0027f
C15226 a_22636_29383# a_22548_29480# 0.28563f
C15227 a_2812_14136# VPWR 0.30213f
C15228 _246_.B2 VPWR 1.53725f
C15229 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I a_58836_18884# 0.02618f
C15230 a_27328_25227# a_28256_25597# 1.16391f
C15231 a_37892_15748# a_38564_15748# 0.00347f
C15232 a_37360_19325# a_37964_18191# 0.00131f
C15233 a_6084_29480# VPWR 0.20348f
C15234 a_57132_12135# VPWR 0.32337f
C15235 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN clk 0.05152f
C15236 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I VPWR 0.79491f
C15237 a_34532_2824# a_35204_2824# 0.00347f
C15238 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I a_62508_21976# 0.00452f
C15239 a_29232_29931# _371_.A1 0.00132f
C15240 a_62420_22020# vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I 0.0042f
C15241 _370_.ZN a_30388_28776# 0.00113f
C15242 a_43268_31048# VPWR 0.20482f
C15243 a_64884_26724# VPWR 0.15276f
C15244 _334_.A1 a_38472_30169# 0.01844f
C15245 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN VPWR 0.76404f
C15246 a_59332_29816# _246_.B2 0.00166f
C15247 _388_.B _386_.A4 0.02486f
C15248 a_19612_24679# VPWR 0.32678f
C15249 a_45128_26031# _402_.ZN 0.00472f
C15250 _417_.A2 _427_.A2 0.41183f
C15251 a_24900_21640# a_25012_20452# 0.02666f
C15252 a_43916_16839# a_43940_15748# 0.0016f
C15253 _378_.I uio_out[7] 0.1629f
C15254 _281_.ZN VPWR 2.16339f
C15255 a_32156_15704# VPWR 0.29679f
C15256 _417_.A2 a_51196_21543# 0.01341f
C15257 _301_.Z a_39172_22504# 0.00246f
C15258 _436_.B _451_.Q 0.10034f
C15259 a_1916_9432# a_2364_9432# 0.0131f
C15260 a_4516_9476# a_4156_9432# 0.08674f
C15261 _371_.A1 _335_.ZN 0.14889f
C15262 _381_.Z a_49044_28292# 0.00525f
C15263 a_13004_30951# uio_oe[3] 0.01121f
C15264 _474_.CLK a_53548_24679# 0.00599f
C15265 _416_.A1 _393_.A1 0.38919f
C15266 a_61188_15368# a_61052_14136# 0.00154f
C15267 _363_.Z a_33060_31048# 0.00107f
C15268 a_51556_14180# a_51644_14136# 0.28563f
C15269 a_47612_18407# VPWR 0.31399f
C15270 a_47612_14136# a_48060_14136# 0.01288f
C15271 a_51308_16839# VPWR 0.31389f
C15272 a_63652_1256# VPWR 0.20348f
C15273 _384_.A1 a_53704_23219# 0.03509f
C15274 _370_.B _459_.CLK 0.29054f
C15275 a_59820_13703# a_59844_12612# 0.0016f
C15276 _416_.A3 a_47028_18884# 0.00882f
C15277 a_56036_28292# a_56124_28248# 0.28563f
C15278 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I clk 0.00114f
C15279 a_39684_20452# VPWR 0.19456f
C15280 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.74483f
C15281 a_45620_17316# VPWR 0.21241f
C15282 a_64884_10664# a_64772_9476# 0.02666f
C15283 a_26108_1159# a_26468_1256# 0.08717f
C15284 a_56796_1592# VPWR 0.33245f
C15285 a_2276_12232# a_2724_12232# 0.01328f
C15286 _397_.A1 a_52848_25987# 0.00195f
C15287 a_53660_12568# a_53572_11044# 0.00151f
C15288 a_18852_1636# a_19300_1636# 0.01328f
C15289 a_56012_12135# a_56372_12232# 0.08663f
C15290 _474_.Q a_50644_21640# 0.00196f
C15291 _448_.Q a_40332_21543# 0.03335f
C15292 a_3260_21543# VPWR 0.30487f
C15293 _452_.Q a_40220_19975# 0.03465f
C15294 vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I VPWR 0.71372f
C15295 a_45172_17316# a_44812_17272# 0.0869f
C15296 a_52415_31220# _268_.A1 0.02222f
C15297 a_43716_2824# VPWR 0.20348f
C15298 _230_.I a_59620_27208# 0.00251f
C15299 a_62980_1636# a_62620_1592# 0.08663f
C15300 a_20508_23111# a_20420_23208# 0.28563f
C15301 a_24092_24679# a_24004_24776# 0.28563f
C15302 a_15156_24776# a_15604_24776# 0.01328f
C15303 _319_.A3 a_36612_20072# 0.00658f
C15304 _433_.ZN _447_.Q 0.0095f
C15305 a_46716_9432# VPWR 0.31143f
C15306 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I 0.00406f
C15307 a_61052_27815# a_61412_27912# 0.0869f
C15308 a_56260_14180# VPWR 0.20348f
C15309 _325_.A2 a_37408_18504# 0.00147f
C15310 a_30724_18504# a_31172_18504# 0.01328f
C15311 _284_.A2 a_44500_25156# 0.01051f
C15312 a_5188_31048# a_5052_29816# 0.00154f
C15313 a_44836_15748# a_45284_15748# 0.01328f
C15314 vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I VPWR 0.96123f
C15315 a_50996_12232# VPWR 0.2093f
C15316 a_41252_15748# a_41340_15704# 0.28563f
C15317 a_57940_18884# a_57580_18840# 0.0869f
C15318 _362_.ZN a_33028_27912# 0.00651f
C15319 _412_.A1 _419_.A4 0.61949f
C15320 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I a_56796_15271# 0.00257f
C15321 a_24004_24776# VPWR 0.20622f
C15322 a_55312_22340# a_55208_22505# 0.10745f
C15323 a_54824_22045# _427_.ZN 0.26624f
C15324 _381_.Z _284_.A2 0.03529f
C15325 a_43400_18909# a_43784_19369# 1.16391f
C15326 _294_.A2 a_31484_26680# 0.04073f
C15327 a_50860_16839# a_50884_15748# 0.0016f
C15328 a_6172_2727# a_6532_2824# 0.08717f
C15329 a_32292_21640# a_32180_20452# 0.02666f
C15330 a_30500_21640# a_30476_20408# 0.0016f
C15331 a_45820_15704# VPWR 0.35662f
C15332 a_33052_19975# a_32964_20072# 0.28563f
C15333 a_22548_29480# a_22548_28292# 0.05841f
C15334 _251_.A1 a_57168_26724# 0.00634f
C15335 _384_.A3 a_51618_22504# 0.00737f
C15336 a_67436_19975# VPWR 0.32937f
C15337 _431_.A3 a_39860_25156# 0.00106f
C15338 _229_.I vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.00176f
C15339 a_2364_14136# a_2364_13703# 0.05841f
C15340 _459_.Q a_31396_26724# 0.00636f
C15341 a_55364_14180# a_55004_14136# 0.08717f
C15342 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I 0.75616f
C15343 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN ena 0.04703f
C15344 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I _274_.A2 0.02717f
C15345 _474_.CLK vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.01013f
C15346 _351_.ZN a_25232_27165# 0.00506f
C15347 a_24304_26795# a_24860_27209# 0.8399f
C15348 vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN a_58476_13703# 0.0011f
C15349 a_56124_2727# a_56572_2727# 0.0131f
C15350 a_4604_12568# a_5052_12568# 0.01222f
C15351 a_66764_13703# a_66788_12612# 0.0016f
C15352 a_36660_23588# _437_.ZN 0.00103f
C15353 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN 0.0194f
C15354 a_53660_17272# VPWR 0.34784f
C15355 a_18096_27165# a_18740_25156# 0.00111f
C15356 a_2276_9096# a_2276_7908# 0.05841f
C15357 a_6620_1159# VPWR 0.3289f
C15358 a_37532_1159# a_37444_1256# 0.28563f
C15359 a_67212_12135# a_67124_12232# 0.28563f
C15360 a_3172_7528# a_3172_6340# 0.05841f
C15361 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN a_57132_18407# 0.00115f
C15362 a_4068_5960# a_4068_4772# 0.05841f
C15363 a_34396_21543# VPWR 0.31319f
C15364 _438_.ZN a_40004_22020# 0.00146f
C15365 a_22059_26399# a_21876_25156# 0.00123f
C15366 a_49092_17316# a_49180_17272# 0.28563f
C15367 _370_.B _371_.A3 0.0109f
C15368 a_52676_17316# a_53124_17316# 0.01328f
C15369 a_65084_1592# a_65532_1592# 0.0131f
C15370 a_67684_1636# a_67324_1592# 0.08674f
C15371 a_27676_26680# a_27676_26247# 0.05841f
C15372 a_3260_10567# a_3620_10664# 0.08717f
C15373 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_55228_28248# 0.031f
C15374 a_57132_10567# a_57580_10567# 0.01288f
C15375 a_66116_2824# VPWR 0.2417f
C15376 a_40264_30320# uo_out[3] 0.0034f
C15377 a_19076_23208# a_19524_23208# 0.01328f
C15378 a_31036_23111# a_31396_23208# 0.08707f
C15379 _452_.CLK a_34448_25597# 0.04094f
C15380 _455_.Q a_26160_27165# 0.00429f
C15381 _337_.A3 a_25232_27165# 0.00457f
C15382 a_25436_21543# a_25884_21543# 0.012f
C15383 a_57692_9432# VPWR 0.31961f
C15384 a_2724_23588# VPWR 0.20782f
C15385 a_4156_21543# a_4068_21640# 0.28563f
C15386 a_2724_6340# VPWR 0.20782f
C15387 a_4516_3204# VPWR 0.20862f
C15388 a_1380_29480# a_1380_28292# 0.05841f
C15389 a_63652_2824# a_63652_1636# 0.05841f
C15390 a_64636_14136# VPWR 0.33393f
C15391 _231_.ZN a_59226_25156# 0.00229f
C15392 a_38816_27555# a_39884_27815# 0.00506f
C15393 a_31820_25112# VPWR 0.33057f
C15394 a_4964_11044# VPWR 0.21167f
C15395 _252_.ZN _247_.B 0.05353f
C15396 a_63964_19975# a_64324_20072# 0.08717f
C15397 a_50660_20452# VPWR 0.21651f
C15398 a_56932_2824# a_57380_2824# 0.01328f
C15399 _386_.ZN a_47700_28292# 0.0118f
C15400 a_67100_18840# a_66988_18407# 0.02634f
C15401 _428_.Z _384_.A1 0.08832f
C15402 _427_.B2 a_49988_21236# 0.00216f
C15403 a_1020_26247# VPWR 0.30073f
C15404 a_31172_18884# VPWR 0.20348f
C15405 a_17596_2727# a_17508_2824# 0.28563f
C15406 a_62732_26680# a_63180_26680# 0.01255f
C15407 _359_.B a_32916_29860# 0.01497f
C15408 a_27140_26344# a_27588_26344# 0.01328f
C15409 _370_.B uo_out[7] 0.35004f
C15410 _454_.Q a_25124_28776# 0.2252f
C15411 a_54692_9476# a_54332_9432# 0.08717f
C15412 _417_.A2 a_50196_21640# 0.00193f
C15413 _398_.C a_53548_24679# 0.00301f
C15414 a_63204_14180# a_63652_14180# 0.01328f
C15415 _408_.ZN a_51048_26680# 0.00165f
C15416 _261_.ZN _447_.Q 0.41464f
C15417 _452_.CLK a_33636_21640# 0.06495f
C15418 a_51556_12612# a_51196_12568# 0.08707f
C15419 a_63764_13800# a_63652_12612# 0.02666f
C15420 a_29020_1159# VPWR 0.29679f
C15421 a_48508_1159# a_48868_1256# 0.08717f
C15422 a_17844_24776# a_17844_23588# 0.05841f
C15423 _454_.D a_22620_27599# 0.24661f
C15424 a_22064_27912# a_23627_27967# 0.41635f
C15425 _340_.A2 VPWR 1.48858f
C15426 _416_.A1 _264_.B 0.19712f
C15427 a_63764_12232# a_64212_12232# 0.01328f
C15428 _452_.Q a_41536_17636# 0.00231f
C15429 a_28932_1636# a_29020_1592# 0.28563f
C15430 a_24988_1592# a_25436_1592# 0.01288f
C15431 a_37532_26247# a_37444_26344# 0.28563f
C15432 a_31396_21640# VPWR 0.20692f
C15433 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_58500_26344# 0.07348f
C15434 _281_.ZN a_51240_23340# 0.03877f
C15435 a_4740_29480# a_4940_27815# 0.00119f
C15436 _319_.A3 a_35968_20937# 0.00145f
C15437 a_54220_10567# a_54132_10664# 0.28563f
C15438 a_53348_1636# a_53212_1159# 0.00168f
C15439 a_49404_1592# a_49404_1159# 0.05841f
C15440 a_14148_2824# a_14148_1636# 0.05841f
C15441 a_10340_2824# a_10204_1592# 0.00154f
C15442 _452_.Q _325_.B 0.00272f
C15443 a_60852_28292# a_60492_28248# 0.08674f
C15444 _459_.Q VPWR 2.76735f
C15445 _355_.C a_27228_26247# 0.01136f
C15446 a_3620_22020# VPWR 0.22347f
C15447 _330_.A1 a_35988_18504# 0.00124f
C15448 a_65756_5863# VPWR 0.31505f
C15449 a_5388_8999# VPWR 0.35526f
C15450 a_21068_23544# VPWR 0.31547f
C15451 a_1828_18884# a_2276_18884# 0.01328f
C15452 a_9084_2727# VPWR 0.31143f
C15453 a_58924_13703# VPWR 0.29679f
C15454 a_24092_21543# a_24452_21640# 0.08707f
C15455 _334_.A1 a_36548_26724# 0.00124f
C15456 a_14596_29480# a_14708_28292# 0.02666f
C15457 _359_.B _402_.A1 0.00865f
C15458 _459_.CLK a_28556_29167# 0.0481f
C15459 _443_.D a_37444_26724# 0.01474f
C15460 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I a_55340_26680# 0.01025f
C15461 _324_.C a_57244_27815# 0.00408f
C15462 a_54020_11044# VPWR 0.20595f
C15463 a_50972_15704# a_51420_15704# 0.01288f
C15464 a_5052_26680# VPWR 0.33516f
C15465 a_24564_31048# _340_.A2 0.00321f
C15466 a_57132_23544# a_57580_23544# 0.0131f
C15467 _319_.ZN a_33052_19975# 0.00131f
C15468 a_62532_15748# a_62620_15704# 0.28563f
C15469 _319_.ZN a_34732_18407# 0.00134f
C15470 _438_.A2 a_37444_25156# 0.00168f
C15471 _336_.A2 a_28124_26680# 0.00417f
C15472 a_22352_25987# VPWR 0.51073f
C15473 a_28572_2727# a_28932_2824# 0.08717f
C15474 _416_.A1 a_44388_27912# 0.00982f
C15475 _431_.A3 a_38616_24328# 0.00765f
C15476 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN a_67772_24679# 0.00215f
C15477 a_16140_28248# VPWR 0.29679f
C15478 a_2724_23588# a_2812_23544# 0.28563f
C15479 a_1828_7908# a_1916_7864# 0.28563f
C15480 _455_.Q _351_.A2 0.31104f
C15481 _251_.A1 a_56036_28292# 0.00348f
C15482 a_2724_6340# a_2812_6296# 0.28563f
C15483 _461_.D VPWR 0.49965f
C15484 a_4516_3204# a_4604_3160# 0.28563f
C15485 a_3620_4772# a_3708_4728# 0.28563f
C15486 a_56348_14136# a_56460_13703# 0.02634f
C15487 a_19412_20452# a_19860_20452# 0.01328f
C15488 _412_.A1 a_51048_26680# 0.01282f
C15489 _399_.A1 _475_.Q 0.03682f
C15490 a_1020_30951# a_1380_31048# 0.08717f
C15491 a_53212_27815# a_53660_27815# 0.01255f
C15492 a_53704_23219# clk 0.00168f
C15493 _294_.A2 _362_.ZN 0.05144f
C15494 a_40644_29480# uo_out[1] 0.01597f
C15495 a_2812_1592# VPWR 0.30213f
C15496 _459_.CLK a_20980_25156# 0.00655f
C15497 _404_.A1 _403_.ZN 0.13654f
C15498 a_54468_12612# a_54556_12568# 0.28563f
C15499 a_58052_12612# a_58500_12612# 0.01328f
C15500 _324_.C a_41476_26344# 0.00313f
C15501 a_23084_30951# a_23108_29860# 0.0016f
C15502 _411_.A2 _282_.ZN 0.02915f
C15503 a_24900_24776# a_24788_23588# 0.02666f
C15504 a_36148_21976# a_36764_22512# 0.00478f
C15505 a_51420_1159# VPWR 0.3289f
C15506 a_4964_11044# a_5052_11000# 0.28563f
C15507 a_59932_1159# a_59844_1256# 0.28563f
C15508 a_50796_19001# VPWR 0.00272f
C15509 a_31708_1592# a_32380_1592# 0.00544f
C15510 _346_.A2 a_22992_27555# 0.02995f
C15511 _244_.Z a_60828_26680# 0.01278f
C15512 a_42236_27815# a_42596_27912# 0.0869f
C15513 _311_.A2 a_37472_24419# 0.00527f
C15514 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN 0.06719f
C15515 a_36404_19001# VPWR 0.00246f
C15516 a_50996_10664# a_51444_10664# 0.01328f
C15517 a_20060_1159# a_20508_1159# 0.0131f
C15518 a_64972_10567# a_65332_10664# 0.08717f
C15519 _384_.ZN a_48321_23208# 0.02366f
C15520 a_36076_18407# a_36100_17316# 0.0016f
C15521 a_60909_30600# _230_.I 0.0023f
C15522 a_21964_21976# VPWR 0.34431f
C15523 a_67996_21976# a_68020_20452# 0.00144f
C15524 _416_.A3 a_45696_20072# 0.02967f
C15525 _223_.I _371_.A1 0.2356f
C15526 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I a_51084_28248# 0.0283f
C15527 _287_.A1 _284_.ZN 0.00584f
C15528 _313_.ZN VPWR 0.79764f
C15529 a_31620_18884# a_31260_18840# 0.08717f
C15530 a_31484_2727# VPWR 0.31605f
C15531 a_52415_31220# _474_.CLK 0.00245f
C15532 a_52788_13800# VPWR 0.20862f
C15533 a_22660_21640# a_23108_21640# 0.01328f
C15534 _450_.D a_42996_18840# 0.00693f
C15535 _474_.CLK ui_in[7] 0.33557f
C15536 a_66428_15271# a_66876_15271# 0.01222f
C15537 a_41056_30669# _459_.CLK 0.00212f
C15538 a_8188_29816# VPWR 0.3582f
C15539 a_67684_11044# VPWR 0.21167f
C15540 a_1020_15271# a_932_15368# 0.28563f
C15541 _324_.B _419_.Z 0.01145f
C15542 a_19724_21976# a_19612_21543# 0.02634f
C15543 _352_.A2 a_31932_26247# 0.00202f
C15544 _246_.B2 a_60404_28292# 0.04555f
C15545 _437_.ZN a_36860_23111# 0.0091f
C15546 a_19164_23111# VPWR 0.33846f
C15547 _432_.ZN a_40656_23588# 0.00635f
C15548 _261_.ZN a_40004_23233# 0.01251f
C15549 a_2364_15271# a_2812_15271# 0.0131f
C15550 a_20308_27912# VPWR 0.20469f
C15551 _399_.A2 _324_.B 0.03755f
C15552 _285_.Z a_37584_29123# 0.00289f
C15553 a_64412_17272# a_64324_15748# 0.00151f
C15554 _324_.C _284_.A2 0.36132f
C15555 a_61524_23208# a_61972_23208# 0.01328f
C15556 a_39996_2727# a_39908_2824# 0.28563f
C15557 vgaringosc.workerclkbuff_notouch_.I a_44160_29123# 0.00146f
C15558 _355_.C _336_.A2 0.49956f
C15559 a_61836_16839# a_62196_16936# 0.08717f
C15560 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN 0.0506f
C15561 a_20084_23588# a_20532_23588# 0.01328f
C15562 a_16500_23588# a_16588_23544# 0.28563f
C15563 a_20868_1256# a_21316_1256# 0.01328f
C15564 a_65668_9476# a_65308_9432# 0.08717f
C15565 a_67012_9476# a_67460_9476# 0.01328f
C15566 a_64860_7864# a_65308_7864# 0.0131f
C15567 a_67012_7908# a_67100_7864# 0.28563f
C15568 a_5052_6296# a_4940_5863# 0.02634f
C15569 a_65756_6296# a_66204_6296# 0.0131f
C15570 a_67908_6340# a_67996_6296# 0.28563f
C15571 a_40196_31048# uo_out[3] 0.00265f
C15572 a_1380_25156# a_1468_25112# 0.28563f
C15573 a_67684_14180# a_67660_13703# 0.00172f
C15574 a_58028_18840# VPWR 0.3521f
C15575 a_66652_4728# a_67100_4728# 0.0131f
C15576 a_50188_13703# a_50636_13703# 0.01288f
C15577 a_67548_3160# a_67996_3160# 0.012f
C15578 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN 0.17717f
C15579 a_25012_20452# a_25100_20408# 0.28563f
C15580 _359_.B a_36656_29123# 0.01219f
C15581 a_39236_26344# a_39684_26344# 0.01328f
C15582 a_14908_30951# a_14820_31048# 0.28563f
C15583 a_11324_29383# a_11772_29383# 0.0131f
C15584 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I rst_n 0.00641f
C15585 _255_.I vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I 0.0015f
C15586 _416_.A1 a_44786_24120# 0.00499f
C15587 a_65308_17272# a_65420_16839# 0.02634f
C15588 a_16612_1636# VPWR 0.22423f
C15589 a_2812_30951# a_3260_30951# 0.0131f
C15590 a_68020_13800# a_68108_12135# 0.0027f
C15591 a_66228_20452# a_66092_19975# 0.00168f
C15592 _274_.ZN VPWR 0.21497f
C15593 a_40244_18180# _452_.D 0.00126f
C15594 _412_.A1 _381_.A2 0.00153f
C15595 _402_.A1 _424_.B1 0.00968f
C15596 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I vgaringosc.workerclkbuff_notouch_.I 0.06168f
C15597 a_41564_26247# _451_.Q 0.00541f
C15598 a_67460_9096# VPWR 0.20924f
C15599 a_45372_11000# a_45820_11000# 0.01288f
C15600 a_49316_11044# a_49404_11000# 0.28563f
C15601 a_66900_18504# a_66988_16839# 0.00151f
C15602 a_3172_18504# VPWR 0.20993f
C15603 a_65556_23588# a_65644_23544# 0.28563f
C15604 a_38652_1592# a_39100_1592# 0.01288f
C15605 a_36436_16936# a_36884_16936# 0.01328f
C15606 a_53548_24679# a_53996_24679# 0.01255f
C15607 a_932_26724# a_1380_26724# 0.01328f
C15608 a_40668_19975# _327_.Z 0.03396f
C15609 _459_.CLK a_23644_24679# 0.00813f
C15610 _359_.B _495_.I 0.05118f
C15611 _284_.ZN _293_.A2 1.95126f
C15612 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN 0.4361f
C15613 a_28556_29167# uo_out[7] 0.005f
C15614 a_65084_1592# a_65084_1159# 0.05841f
C15615 a_37408_18504# a_37980_17272# 0.00105f
C15616 _330_.ZN a_37532_17272# 0.00377f
C15617 _419_.A4 _473_.Q 0.52555f
C15618 _316_.ZN VPWR 0.76683f
C15619 _355_.C _346_.A2 0.11075f
C15620 a_47612_30951# a_48060_30951# 0.0131f
C15621 a_35728_29480# a_36284_29167# 0.8399f
C15622 a_2364_12568# VPWR 0.30029f
C15623 a_58588_21543# a_58500_21640# 0.28563f
C15624 _330_.A1 a_41572_18504# 0.00157f
C15625 a_53660_2727# VPWR 0.33981f
C15626 a_3620_26344# a_4068_26344# 0.01328f
C15627 a_17932_26247# a_18628_26344# 0.01227f
C15628 _452_.CLK a_38816_27555# 0.00161f
C15629 a_58588_26247# _251_.ZN 0.00582f
C15630 a_66900_16936# a_66876_15271# 0.00134f
C15631 a_63068_18407# a_62980_18504# 0.28563f
C15632 _384_.ZN _390_.ZN 0.36403f
C15633 _386_.ZN _402_.A1 0.02662f
C15634 a_23556_29860# VPWR 0.21403f
C15635 a_36860_15271# a_37220_15368# 0.08717f
C15636 a_38316_20408# _323_.A3 0.00236f
C15637 a_54668_10567# VPWR 0.31547f
C15638 _362_.B a_35728_29480# 0.01137f
C15639 a_26668_21976# a_26556_21543# 0.02634f
C15640 a_16500_23208# VPWR 0.20348f
C15641 _428_.Z clk 0.04369f
C15642 a_58539_30644# ui_in[4] 0.00145f
C15643 _294_.A2 _287_.A2 1.02855f
C15644 a_3172_28292# a_2812_28248# 0.08717f
C15645 a_57916_25112# vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN 0.00209f
C15646 a_3620_22020# a_3708_21976# 0.28563f
C15647 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I 0.14057f
C15648 a_50972_2727# a_51332_2824# 0.08717f
C15649 a_67012_17316# a_67100_17272# 0.28563f
C15650 a_47076_18504# a_47524_18504# 0.01328f
C15651 a_18740_25156# a_19188_25156# 0.01328f
C15652 a_15156_25156# a_15244_25112# 0.28563f
C15653 _451_.Q _433_.ZN 0.07532f
C15654 a_30388_20452# a_30836_20452# 0.01328f
C15655 a_61052_14136# a_61076_13800# 0.00172f
C15656 a_52900_26724# _412_.ZN 0.00467f
C15657 a_47164_13703# a_47076_13800# 0.28563f
C15658 a_14004_31048# uio_oe[1] 0.00329f
C15659 a_55140_20452# a_54780_20408# 0.0869f
C15660 a_24652_30951# _342_.ZN 0.00203f
C15661 a_22996_31048# _459_.CLK 0.00652f
C15662 a_33948_16839# a_33860_16936# 0.28563f
C15663 a_61500_11000# a_61412_9476# 0.00151f
C15664 a_30276_1636# VPWR 0.20348f
C15665 a_64636_12568# a_65084_12568# 0.01288f
C15666 _419_.A4 _475_.D 0.00789f
C15667 vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I 0.00322f
C15668 a_21740_29383# a_22188_29383# 0.01255f
C15669 _284_.B a_42784_25640# 0.00263f
C15670 a_1828_1636# a_2276_1636# 0.01328f
C15671 a_65756_26247# vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I 0.02009f
C15672 _452_.CLK a_45820_18840# 0.01452f
C15673 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN a_65668_26344# 0.00331f
C15674 a_55028_12232# a_55116_10567# 0.00151f
C15675 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN 0.00176f
C15676 a_45956_1636# a_45596_1592# 0.08707f
C15677 _362_.B a_35756_27216# 0.00322f
C15678 vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN 0.04023f
C15679 a_54892_23544# VPWR 0.32089f
C15680 _267_.A2 a_59572_29076# 0.43937f
C15681 _249_.A2 clk 0.0246f
C15682 _260_.A1 a_40656_23588# 0.01438f
C15683 a_54780_15704# a_54916_15368# 0.00168f
C15684 a_42236_1159# a_42908_1159# 0.00544f
C15685 a_53796_20452# a_54244_20452# 0.01328f
C15686 a_1380_27912# a_1380_26724# 0.05841f
C15687 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN a_58388_20452# 0.00129f
C15688 a_55340_24679# a_55252_24776# 0.28563f
C15689 a_17036_20408# VPWR 0.31143f
C15690 _427_.B1 a_52852_24372# 0.53347f
C15691 _474_.CLK _384_.A3 0.09872f
C15692 a_55812_12612# VPWR 0.20595f
C15693 a_66900_16936# a_67348_16936# 0.01328f
C15694 a_9980_29383# a_9892_29480# 0.28563f
C15695 a_46404_15368# a_46852_15368# 0.01328f
C15696 _342_.ZN a_25792_30301# 0.00666f
C15697 a_24864_29931# a_25420_30345# 0.8399f
C15698 a_48420_10664# VPWR 0.20924f
C15699 a_48284_15271# a_48196_15368# 0.28563f
C15700 a_56596_23588# VPWR 0.20907f
C15701 _267_.A1 a_56484_29480# 0.00142f
C15702 _370_.ZN a_25124_28776# 0.00347f
C15703 a_1020_4295# a_1380_4392# 0.08717f
C15704 a_36996_26724# a_37084_26680# 0.28563f
C15705 _260_.A1 a_42728_20452# 0.00147f
C15706 _287_.A1 _223_.ZN 0.08265f
C15707 a_37179_24831# a_37108_23588# 0.00126f
C15708 a_49852_15271# a_50300_15271# 0.0131f
C15709 _334_.A1 a_34084_28776# 0.28037f
C15710 a_63964_15271# VPWR 0.29679f
C15711 _459_.Q _370_.B 0.02066f
C15712 a_19328_28733# _378_.ZN 0.00114f
C15713 a_62396_2727# a_62308_2824# 0.28563f
C15714 a_20980_22020# a_21428_22020# 0.01328f
C15715 a_17396_22020# a_17484_21976# 0.28563f
C15716 _265_.ZN _451_.Q 0.00438f
C15717 a_67548_15704# VPWR 0.32971f
C15718 a_27004_27815# VPWR 0.35877f
C15719 a_31260_16839# a_31708_16839# 0.0131f
C15720 _436_.B a_40220_26247# 0.00806f
C15721 a_46716_30951# a_46628_31048# 0.28563f
C15722 a_42154_21236# a_42610_21812# 0.00165f
C15723 a_27812_23208# a_27900_21543# 0.00151f
C15724 _324_.B _416_.A2 0.00115f
C15725 a_27564_23544# a_28012_23544# 0.01222f
C15726 _365_.ZN uo_out[4] 0.00245f
C15727 a_66564_7908# VPWR 0.20631f
C15728 a_18404_1256# VPWR 0.20839f
C15729 a_43268_1256# a_43716_1256# 0.01328f
C15730 a_64412_4728# VPWR 0.3038f
C15731 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN a_57580_18840# 0.00472f
C15732 a_55004_14136# a_54916_12612# 0.00151f
C15733 a_4068_13800# a_4852_13800# 0.00276f
C15734 _272_.B1 a_57220_29861# 0.13363f
C15735 a_22300_2727# a_22748_2727# 0.0131f
C15736 a_9084_29383# VPWR 0.3289f
C15737 a_58028_13703# a_58388_13800# 0.08707f
C15738 a_57020_23111# vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN 0.00355f
C15739 _351_.A2 a_25108_27508# 0.00994f
C15740 _267_.A2 _257_.B 0.31898f
C15741 _397_.A1 _284_.B 0.79397f
C15742 a_43940_27912# a_43564_27209# 0.00189f
C15743 _330_.A1 a_43008_26795# 0.0372f
C15744 a_44812_16839# a_45172_16936# 0.08707f
C15745 a_50100_10664# a_49988_9476# 0.02666f
C15746 a_36412_1592# VPWR 0.3289f
C15747 _474_.CLK a_54824_22045# 0.16655f
C15748 _324_.C a_52452_24072# 0.0016f
C15749 a_3708_1159# a_3620_1256# 0.28563f
C15750 a_33860_16936# VPWR 0.21375f
C15751 _437_.A1 a_37644_23544# 0.0432f
C15752 a_60492_28248# VPWR 0.31552f
C15753 a_61948_12568# a_62060_12135# 0.02634f
C15754 _424_.A2 a_52452_21236# 0.0273f
C15755 a_37384_19624# VPWR 0.31792f
C15756 a_3620_29860# a_3708_29816# 0.28563f
C15757 a_7204_29860# a_7652_29860# 0.01328f
C15758 a_4604_17272# a_5052_17272# 0.01222f
C15759 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I 0.0586f
C15760 a_45148_30951# VPWR 0.31143f
C15761 a_48868_1636# a_48956_1592# 0.28563f
C15762 a_52452_1636# a_52900_1636# 0.01328f
C15763 a_59036_11000# a_59484_11000# 0.01288f
C15764 a_45820_11000# a_45820_10567# 0.05841f
C15765 a_49764_11044# a_49740_10567# 0.00172f
C15766 _301_.A1 _438_.ZN 0.03906f
C15767 _452_.CLK _447_.Q 0.06984f
C15768 a_60604_27815# a_61052_27815# 0.01255f
C15769 _370_.B _461_.D 0.28784f
C15770 a_1020_23111# a_1468_23111# 0.0131f
C15771 a_48508_18407# a_48420_18504# 0.28563f
C15772 a_66316_20408# a_66116_18884# 0.00119f
C15773 a_50324_18504# a_50412_16839# 0.00151f
C15774 _346_.ZN a_20756_26724# 0.00449f
C15775 a_43796_18559# VPWR 0.00246f
C15776 a_67012_18884# a_66652_18840# 0.0869f
C15777 a_16500_25156# VPWR 0.20348f
C15778 a_28012_20408# VPWR 0.31143f
C15779 a_15692_27815# a_16052_27912# 0.08717f
C15780 a_1380_27912# a_1828_27912# 0.01328f
C15781 _452_.CLK a_33584_22137# 0.001f
C15782 a_62396_12568# VPWR 0.31389f
C15783 a_23108_2824# a_23780_2824# 0.00347f
C15784 a_20308_26724# uio_out[7] 0.00146f
C15785 _451_.Q _261_.ZN 0.001f
C15786 hold2.Z _260_.A1 0.00193f
C15787 a_932_9096# a_932_7908# 0.05841f
C15788 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I 0.03402f
C15789 a_17396_21640# a_17396_20452# 0.05841f
C15790 a_43232_29480# VPWR 1.0975f
C15791 a_64436_16936# VPWR 0.2098f
C15792 _416_.A3 a_47047_21640# 0.00132f
C15793 a_43940_15368# VPWR 0.20348f
C15794 a_57380_16936# vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN 0.00326f
C15795 a_47388_15271# VPWR 0.29679f
C15796 a_4604_14136# a_5052_14136# 0.01222f
C15797 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62564_29032# 0.01858f
C15798 _349_.A4 a_25796_27912# 0.00133f
C15799 _455_.D a_21868_27208# 0.00881f
C15800 a_3708_16839# VPWR 0.33374f
C15801 a_64212_23208# vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN 0.0097f
C15802 _393_.ZN a_45484_28248# 0.01013f
C15803 a_40804_1256# VPWR 0.20382f
C15804 a_67548_3160# a_67548_2727# 0.05841f
C15805 a_1380_13800# a_1380_12612# 0.05841f
C15806 _397_.A2 _282_.ZN 0.00669f
C15807 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I a_59372_14136# 0.00251f
C15808 _229_.I ui_in[1] 0.05193f
C15809 _386_.A4 _402_.A1 0.02716f
C15810 _474_.CLK a_56684_23544# 0.00581f
C15811 a_14708_23208# a_14708_22020# 0.05841f
C15812 a_2364_17272# VPWR 0.30029f
C15813 a_50212_1636# VPWR 0.22509f
C15814 a_50300_12568# a_50212_11044# 0.00151f
C15815 a_14684_1159# a_15044_1256# 0.08717f
C15816 a_58164_16936# VPWR 0.26218f
C15817 a_58924_12135# a_59372_12135# 0.01288f
C15818 a_7876_29480# a_8548_29480# 0.00347f
C15819 a_29804_23544# a_29692_23111# 0.02634f
C15820 a_15492_1636# a_15940_1636# 0.01328f
C15821 a_11908_1636# a_11996_1592# 0.28563f
C15822 _395_.A1 _474_.Q 0.04371f
C15823 _252_.B _231_.ZN 0.00253f
C15824 a_57132_18407# VPWR 0.31795f
C15825 a_59226_25156# clk 0.00211f
C15826 a_36996_17316# a_36636_17272# 0.08707f
C15827 a_45060_31048# a_45508_31048# 0.01328f
C15828 a_20868_2824# VPWR 0.20815f
C15829 a_28124_1592# a_28124_1159# 0.05841f
C15830 _459_.Q _360_.ZN 0.03748f
C15831 _330_.A1 a_38752_26344# 0.00868f
C15832 a_66340_11044# a_66428_11000# 0.28563f
C15833 _459_.CLK a_20756_26724# 0.00683f
C15834 _424_.A1 a_52024_20083# 0.04463f
C15835 _452_.Q _441_.A2 0.50528f
C15836 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_64884_26724# 0.00434f
C15837 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_63092_26724# 0.0155f
C15838 a_54356_24776# VPWR 0.20348f
C15839 _285_.Z a_38584_28292# 0.04296f
C15840 a_21404_24679# a_21852_24679# 0.01288f
C15841 a_52900_26724# a_53908_26724# 0.00196f
C15842 a_3708_24679# a_3620_24776# 0.28563f
C15843 a_4156_19975# a_4940_19975# 0.00443f
C15844 a_64636_1159# a_65084_1159# 0.0131f
C15845 _250_.A2 a_62756_27912# 0.00181f
C15846 a_63180_26680# _245_.I1 0.00399f
C15847 a_1828_5960# a_2276_5960# 0.01328f
C15848 a_22188_29383# a_22548_29480# 0.0869f
C15849 a_2364_14136# VPWR 0.30029f
C15850 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.00165f
C15851 a_49316_2824# a_49316_1636# 0.05841f
C15852 a_2724_4392# a_3172_4392# 0.01328f
C15853 a_30812_18407# a_31260_18407# 0.0131f
C15854 _352_.A2 a_26548_24372# 0.02683f
C15855 a_57220_29861# VPWR 0.39227f
C15856 _452_.Q a_40416_18885# 0.01388f
C15857 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I a_58388_18884# 0.00409f
C15858 _384_.A3 _398_.C 0.23232f
C15859 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I 0.66091f
C15860 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN a_62172_18840# 0.00245f
C15861 a_56460_12135# VPWR 0.34525f
C15862 a_33948_15704# a_34396_15704# 0.01288f
C15863 a_5636_29480# VPWR 0.21011f
C15864 a_37892_15748# a_37980_15704# 0.28563f
C15865 _370_.ZN a_29835_28776# 0.00627f
C15866 a_62420_22020# a_62508_21976# 0.28563f
C15867 a_42820_31048# VPWR 0.25483f
C15868 _358_.A3 a_36636_26247# 0.00269f
C15869 a_19164_24679# VPWR 0.33846f
C15870 a_45232_25987# _402_.ZN 0.20799f
C15871 a_58116_30344# _246_.B2 0.00227f
C15872 _417_.A2 a_51332_24072# 0.53908f
C15873 _402_.A1 _407_.A1 0.01562f
C15874 a_43003_28409# a_43248_28777# 0.00232f
C15875 a_46156_25112# VPWR 0.3243f
C15876 a_31708_15704# VPWR 0.29679f
C15877 _311_.A2 _316_.A3 0.01022f
C15878 _324_.C vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I 0.08669f
C15879 a_4068_9476# a_4156_9432# 0.28563f
C15880 _381_.Z a_48820_28292# 0.01357f
C15881 a_30388_28776# _335_.ZN 1.37596f
C15882 a_49404_18407# a_50412_18407# 0.00323f
C15883 a_12548_31048# uio_oe[3] 0.12504f
C15884 a_27116_21976# a_27564_21976# 0.01288f
C15885 a_47164_18407# VPWR 0.31268f
C15886 a_53100_16839# a_53548_16839# 0.0131f
C15887 a_51556_14180# a_51196_14136# 0.08707f
C15888 _452_.CLK a_41432_17801# 0.00794f
C15889 a_50860_16839# VPWR 0.32024f
C15890 a_53012_16936# a_53124_15748# 0.02666f
C15891 a_49204_16936# a_49180_15704# 0.0016f
C15892 a_19328_28733# uio_out[6] 0.78773f
C15893 a_63204_1256# VPWR 0.20348f
C15894 a_65668_1256# a_66116_1256# 0.01328f
C15895 a_49652_13800# a_49764_12612# 0.02666f
C15896 a_44700_2727# a_45148_2727# 0.0131f
C15897 a_65780_13800# a_66228_13800# 0.01328f
C15898 a_56036_28292# a_55676_28248# 0.08663f
C15899 a_38676_20452# VPWR 0.20771f
C15900 vgaringosc.workerclkbuff_notouch_.I _392_.A2 0.0046f
C15901 _304_.B _438_.A2 0.19774f
C15902 a_55452_21543# vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.0367f
C15903 a_45172_17316# VPWR 0.20728f
C15904 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I 0.05574f
C15905 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I 0.10555f
C15906 a_56348_1592# VPWR 0.32925f
C15907 a_26108_1159# a_26020_1256# 0.28563f
C15908 a_62172_1592# a_62308_1256# 0.00168f
C15909 _397_.A1 a_52360_26355# 0.04659f
C15910 a_56012_12135# a_55924_12232# 0.28563f
C15911 a_2812_21543# VPWR 0.30213f
C15912 _268_.A2 _274_.A1 0.51328f
C15913 a_13340_29816# a_13788_29816# 0.01288f
C15914 _448_.Q a_38340_21327# 0.01227f
C15915 _452_.Q a_39772_19975# 0.0184f
C15916 a_3620_26344# a_3620_25156# 0.05841f
C15917 a_41048_17341# a_42460_17801# 0.00393f
C15918 a_44724_17316# a_44812_17272# 0.28563f
C15919 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.65337f
C15920 _230_.I a_59260_26680# 0.02434f
C15921 _397_.A2 a_47412_23588# 0.00244f
C15922 a_45820_10567# a_46268_10567# 0.0131f
C15923 a_58588_1592# a_59036_1592# 0.01288f
C15924 a_62532_1636# a_62620_1592# 0.28563f
C15925 a_43268_2824# VPWR 0.20511f
C15926 a_20060_23111# a_20420_23208# 0.08707f
C15927 a_31932_23111# a_32380_23111# 0.01288f
C15928 a_23644_24679# a_24004_24776# 0.08707f
C15929 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I 0.00407f
C15930 _459_.CLK _378_.I 0.00405f
C15931 a_46268_9432# VPWR 0.31143f
C15932 a_61052_27815# a_60964_27912# 0.28563f
C15933 a_16164_2824# a_16252_1159# 0.0027f
C15934 _294_.A2 a_35008_27533# 0.08987f
C15935 a_55812_14180# VPWR 0.20348f
C15936 _424_.B1 _218_.ZN 0.32685f
C15937 _267_.A1 a_55676_27815# 0.0051f
C15938 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I 0.00738f
C15939 a_36524_18407# a_36436_18504# 0.28563f
C15940 _284_.A2 a_44028_25156# 0.01071f
C15941 _390_.ZN a_51576_25896# 0.00402f
C15942 a_50548_12232# VPWR 0.2414f
C15943 a_41252_15748# a_40892_15704# 0.08707f
C15944 a_45508_2824# a_45956_2824# 0.01328f
C15945 a_57492_18884# a_57580_18840# 0.28563f
C15946 a_3708_20408# a_3708_19975# 0.05841f
C15947 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I a_56348_15271# 0.03293f
C15948 a_23556_24776# VPWR 0.20622f
C15949 a_54824_22045# a_55208_22505# 1.16391f
C15950 _395_.A1 _395_.A2 0.12883f
C15951 _416_.A1 a_41564_24679# 0.00119f
C15952 a_63336_29480# a_63524_29098# 0.00126f
C15953 a_43400_18909# a_43888_19204# 0.8399f
C15954 a_6172_2727# a_6084_2824# 0.28563f
C15955 a_32604_19975# a_32964_20072# 0.08717f
C15956 a_45372_15704# VPWR 0.29679f
C15957 _251_.A1 a_56816_26724# 0.00432f
C15958 a_48508_9432# a_49092_9476# 0.01675f
C15959 _384_.A3 a_51414_22504# 0.01166f
C15960 _384_.A1 _476_.Q 0.00171f
C15961 _384_.ZN _399_.A1 0.08162f
C15962 a_66988_19975# VPWR 0.32963f
C15963 _431_.A3 a_38852_25156# 0.01911f
C15964 hold2.Z _260_.A2 0.05694f
C15965 a_54916_14180# a_55004_14136# 0.28563f
C15966 a_58836_14180# a_59284_14180# 0.01328f
C15967 a_21068_25112# a_20980_23588# 0.00151f
C15968 _452_.CLK a_40668_26247# 0.00706f
C15969 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN a_65756_27815# 0.00365f
C15970 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I _250_.B 0.37882f
C15971 a_24304_26795# a_25232_27165# 1.16391f
C15972 _397_.A1 _474_.Q 0.00304f
C15973 a_8860_1592# a_8996_1256# 0.00168f
C15974 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN a_54892_16839# 0.03698f
C15975 _474_.CLK a_56148_24776# 0.00875f
C15976 _438_.A2 VPWR 1.3096f
C15977 _375_.Z VPWR 0.50153f
C15978 a_53212_17272# VPWR 0.31547f
C15979 a_6172_1159# VPWR 0.3289f
C15980 a_37084_1159# a_37444_1256# 0.08717f
C15981 a_50636_12135# a_50660_11044# 0.0016f
C15982 a_21628_1592# a_22076_1592# 0.01288f
C15983 a_66764_12135# a_67124_12232# 0.08717f
C15984 a_52788_12232# a_53236_12232# 0.01328f
C15985 _451_.Q _327_.Z 1.7915f
C15986 a_4852_4392# a_4964_3204# 0.02666f
C15987 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN a_56684_18407# 0.0072f
C15988 a_33724_21543# VPWR 0.35737f
C15989 vgaringosc.workerclkbuff_notouch_.I _416_.A1 0.52535f
C15990 a_49092_17316# a_48732_17272# 0.08707f
C15991 a_58500_26344# vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN 0.00294f
C15992 a_3260_10567# a_3172_10664# 0.28563f
C15993 a_65668_2824# VPWR 0.23752f
C15994 a_67236_1636# a_67324_1592# 0.28563f
C15995 _327_.A2 a_44724_17316# 0.00162f
C15996 _395_.A1 a_50196_22805# 0.08831f
C15997 a_31036_23111# a_30948_23208# 0.28563f
C15998 _452_.CLK a_33148_25641# 0.00275f
C15999 a_57244_9432# VPWR 0.31684f
C16000 a_2276_23588# VPWR 0.20634f
C16001 _455_.Q a_24860_27209# 0.00817f
C16002 a_64188_14136# VPWR 0.31479f
C16003 a_2276_6340# VPWR 0.20634f
C16004 a_3708_21543# a_4068_21640# 0.08717f
C16005 a_4068_3204# VPWR 0.2157f
C16006 _399_.ZN _324_.B 0.22315f
C16007 _324_.C _419_.A4 0.07697f
C16008 _459_.CLK a_32380_26247# 0.01501f
C16009 vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I 0.07218f
C16010 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN clk 0.03569f
C16011 a_47748_15748# a_48196_15748# 0.01328f
C16012 a_4516_11044# VPWR 0.20862f
C16013 a_11012_29860# a_10876_29383# 0.00168f
C16014 a_29176_25273# VPWR 0.00204f
C16015 a_50212_20452# VPWR 0.1439f
C16016 _256_.A2 a_59572_29076# 0.00129f
C16017 _330_.A1 a_36300_23544# 0.02924f
C16018 a_63964_19975# a_63876_20072# 0.28563f
C16019 _383_.A2 a_48820_28292# 0.0125f
C16020 a_30160_30301# a_30795_29977# 0.02112f
C16021 a_35232_24029# _312_.ZN 0.00127f
C16022 _355_.C _455_.D 0.04542f
C16023 a_22548_29480# a_22996_29480# 0.01328f
C16024 _313_.ZN _311_.Z 0.15902f
C16025 a_30724_18884# VPWR 0.22176f
C16026 a_60276_26724# VPWR 0.00419f
C16027 _296_.ZN a_38472_30169# 0.01326f
C16028 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN VPWR 0.969f
C16029 a_17148_2727# a_17508_2824# 0.08717f
C16030 _379_.A2 _346_.B 0.02227f
C16031 _416_.A1 a_52068_29480# 0.00268f
C16032 _260_.A1 _448_.Q 0.18763f
C16033 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN 0.00135f
C16034 a_54244_9476# a_54332_9432# 0.28563f
C16035 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I a_58924_17272# 0.00285f
C16036 _381_.Z _381_.A2 0.03984f
C16037 a_51868_17272# a_51780_15748# 0.00151f
C16038 _304_.B _475_.Q 0.03085f
C16039 _371_.A1 a_29575_28293# 0.00585f
C16040 a_2812_20408# a_3260_20408# 0.0131f
C16041 _230_.I a_63336_29480# 0.01022f
C16042 _452_.CLK a_33188_21640# 0.01459f
C16043 a_37408_18504# a_39264_18147# 0.02307f
C16044 _334_.A1 a_33776_29123# 0.04436f
C16045 a_51108_12612# a_51196_12568# 0.28563f
C16046 a_47164_12568# a_47612_12568# 0.01288f
C16047 a_67100_2727# a_67548_2727# 0.01222f
C16048 _386_.ZN _386_.A4 0.20748f
C16049 a_48508_1159# a_48420_1256# 0.28563f
C16050 a_22064_27912# a_22620_27599# 0.8399f
C16051 _454_.D a_22992_27555# 0.0057f
C16052 _349_.A4 _343_.A2 0.01143f
C16053 a_28572_1159# VPWR 0.29679f
C16054 a_67324_12568# a_67236_11044# 0.00151f
C16055 a_47524_12232# a_47524_11044# 0.05841f
C16056 a_28932_1636# a_28572_1592# 0.08707f
C16057 a_31484_30951# VPWR 0.32502f
C16058 a_57580_12135# a_57604_11044# 0.0016f
C16059 a_5300_7528# a_5388_5863# 0.0027f
C16060 _452_.Q a_41048_17341# 0.00399f
C16061 a_30948_21640# VPWR 0.20692f
C16062 a_40668_26247# a_41116_26247# 0.01222f
C16063 a_37084_26247# a_37444_26344# 0.08674f
C16064 a_53772_10567# a_54132_10664# 0.08707f
C16065 a_67660_10567# a_68108_10567# 0.0131f
C16066 a_60404_28292# a_60492_28248# 0.28563f
C16067 a_8636_1159# a_9084_1159# 0.0131f
C16068 _256_.A2 _257_.B 0.00824f
C16069 _407_.A1 _424_.B1 0.19069f
C16070 a_51240_19624# VPWR 0.51068f
C16071 a_29804_30951# VPWR 0.32592f
C16072 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN a_63313_28776# 0.00111f
C16073 a_29604_23208# a_30052_23208# 0.01328f
C16074 a_3172_22020# VPWR 0.20993f
C16075 a_33524_24776# a_34308_24776# 0.00276f
C16076 a_4940_8999# VPWR 0.31945f
C16077 a_20620_23544# VPWR 0.31547f
C16078 _334_.A1 a_36100_26724# 0.00383f
C16079 a_65308_5863# VPWR 0.30378f
C16080 a_2276_21640# a_2724_21640# 0.01328f
C16081 a_24092_21543# a_24004_21640# 0.28563f
C16082 a_8636_2727# VPWR 0.31605f
C16083 a_58476_13703# VPWR 0.32508f
C16084 a_38340_2824# a_38428_1159# 0.0027f
C16085 _397_.A1 _395_.A2 0.229f
C16086 _459_.CLK a_28928_29123# 0.01967f
C16087 _443_.D a_36996_26724# 0.00215f
C16088 a_36960_27912# a_37444_26724# 0.00263f
C16089 a_60964_27912# a_61412_27912# 0.01328f
C16090 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I a_54892_26680# 0.00115f
C16091 _324_.C a_56124_27815# 0.00398f
C16092 a_64412_29816# vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.00168f
C16093 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN 0.04868f
C16094 a_53572_11044# VPWR 0.20595f
C16095 _229_.I _324_.C 0.04772f
C16096 a_3260_21976# a_3260_21543# 0.05841f
C16097 a_47164_2727# a_47300_1636# 0.00154f
C16098 a_17148_29816# a_17148_29383# 0.05841f
C16099 a_4604_26680# VPWR 0.33016f
C16100 _397_.A1 a_46984_23588# 0.43787f
C16101 a_62532_15748# a_62172_15704# 0.08717f
C16102 a_65220_15748# a_65668_15748# 0.01328f
C16103 a_10540_30951# uio_oe[5] 0.00187f
C16104 _336_.A2 a_27676_26680# 0.00148f
C16105 a_28036_26724# a_28124_26680# 0.28563f
C16106 a_22059_26399# VPWR 0.37157f
C16107 a_61164_23111# a_61612_23111# 0.0131f
C16108 a_28572_2727# a_28484_2824# 0.28563f
C16109 _325_.ZN a_43664_17317# 0.08864f
C16110 _452_.CLK _451_.Q 0.05635f
C16111 a_59484_9432# a_59932_9432# 0.0131f
C16112 _455_.Q a_24900_27912# 0.11458f
C16113 a_15692_28248# VPWR 0.29679f
C16114 a_4516_23588# a_4964_23588# 0.01328f
C16115 a_2724_23588# a_2364_23544# 0.08717f
C16116 a_9444_1256# a_9892_1256# 0.01328f
C16117 a_1828_7908# a_1468_7864# 0.08717f
C16118 a_3620_7908# a_4068_7908# 0.01328f
C16119 a_1020_4728# a_1468_4728# 0.0131f
C16120 a_3620_4772# a_3260_4728# 0.08717f
C16121 _285_.Z uo_out[3] 0.06787f
C16122 a_2724_6340# a_2364_6296# 0.08717f
C16123 a_4516_6340# a_4964_6340# 0.01328f
C16124 _279_.Z a_48529_22460# 0.20523f
C16125 a_66428_14136# a_66876_14136# 0.01288f
C16126 a_1916_3160# a_2364_3160# 0.0131f
C16127 a_4516_3204# a_4156_3160# 0.08674f
C16128 a_5188_31048# a_5276_29383# 0.0027f
C16129 _475_.Q VPWR 1.83962f
C16130 a_66540_16839# a_66564_15748# 0.0016f
C16131 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_54444_26680# 0.0016f
C16132 a_1020_30951# a_932_31048# 0.28563f
C16133 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN _231_.I 0.74405f
C16134 a_62532_30736# _256_.A2 0.00414f
C16135 a_1020_12568# a_1020_12135# 0.05841f
C16136 a_57044_13800# a_57132_12135# 0.00151f
C16137 a_2364_1592# VPWR 0.30029f
C16138 a_40196_29480# uo_out[1] 0.01602f
C16139 a_54468_12612# a_54108_12568# 0.08707f
C16140 _459_.CLK a_20532_25156# 0.00645f
C16141 _459_.CLK _336_.Z 0.11f
C16142 a_36148_21976# a_36560_22512# 0.00705f
C16143 a_50972_1159# VPWR 0.33191f
C16144 a_59484_1159# a_59844_1256# 0.08717f
C16145 a_35428_1636# a_35876_1636# 0.01328f
C16146 a_2364_11000# a_2812_11000# 0.0131f
C16147 a_4964_11044# a_4604_11000# 0.08674f
C16148 a_33520_25597# a_34155_25273# 0.02112f
C16149 a_54580_12232# a_54468_11044# 0.02666f
C16150 _244_.Z a_59620_27208# 0.37046f
C16151 a_67436_16839# a_67884_16839# 0.012f
C16152 a_49840_19001# VPWR 0.0023f
C16153 _363_.Z _371_.A1 0.02595f
C16154 a_50300_20408# a_50748_20408# 0.01222f
C16155 _442_.ZN _444_.D 0.00744f
C16156 a_42236_27815# a_42148_27912# 0.28563f
C16157 a_64972_10567# a_64884_10664# 0.28563f
C16158 a_37532_25112# a_37472_24419# 0.0065f
C16159 _311_.A2 a_37179_24831# 0.0027f
C16160 _355_.C _454_.D 0.82693f
C16161 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN a_66787_30600# 0.00762f
C16162 a_21516_21976# VPWR 0.31589f
C16163 _223_.I a_30388_28776# 0.01995f
C16164 a_32964_18884# a_33412_18884# 0.01328f
C16165 _352_.ZN a_26756_24801# 0.03791f
C16166 a_33376_23659# VPWR 1.14541f
C16167 a_31172_18884# a_31260_18840# 0.28563f
C16168 a_52415_31220# a_52639_30644# 0.53809f
C16169 a_52340_13800# VPWR 0.20595f
C16170 a_30812_2727# VPWR 0.33981f
C16171 a_2812_26247# a_3260_26247# 0.0131f
C16172 a_52639_30644# ui_in[7] 0.01928f
C16173 a_7740_29816# VPWR 0.3289f
C16174 a_67236_11044# VPWR 0.20622f
C16175 a_18716_23111# VPWR 0.32683f
C16176 _352_.A2 a_30724_26020# 0.50398f
C16177 a_19860_27912# VPWR 0.20788f
C16178 _432_.ZN a_40452_23588# 0.00211f
C16179 _304_.B _402_.ZN 0.00984f
C16180 _242_.Z a_58588_26247# 0.00227f
C16181 _285_.Z a_37291_29535# 0.00314f
C16182 a_39548_2727# a_39908_2824# 0.08717f
C16183 a_61836_16839# a_61748_16936# 0.28563f
C16184 a_54692_18884# vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN 0.00339f
C16185 a_16500_23588# a_16140_23544# 0.08707f
C16186 a_3708_7864# a_3708_7431# 0.05841f
C16187 a_3172_25156# a_3620_25156# 0.01328f
C16188 a_65220_9476# a_65308_9432# 0.28563f
C16189 a_1380_25156# a_1020_25112# 0.08717f
C16190 a_67012_7908# a_66652_7864# 0.08717f
C16191 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.08287f
C16192 a_67908_6340# a_67548_6296# 0.08663f
C16193 a_39748_31048# uo_out[3] 0.00221f
C16194 a_57580_18840# VPWR 0.30535f
C16195 a_53212_14136# a_53236_13800# 0.00172f
C16196 a_64772_20072# a_64772_18884# 0.05841f
C16197 _324_.C rst_n 0.01323f
C16198 a_63740_14136# a_63852_13703# 0.02634f
C16199 a_22860_20408# a_23308_20408# 0.0131f
C16200 a_25012_20452# a_24652_20408# 0.08717f
C16201 _359_.B a_35728_29480# 0.03215f
C16202 a_14460_30951# a_14820_31048# 0.08674f
C16203 _424_.B2 a_51240_19624# 0.01288f
C16204 a_60940_28248# a_60740_26724# 0.00119f
C16205 a_64996_31048# rst_n 0.01765f
C16206 a_16028_1592# VPWR 0.35662f
C16207 _304_.B vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.32475f
C16208 a_51556_12612# a_51532_12135# 0.00172f
C16209 a_47612_12568# a_47612_12135# 0.05841f
C16210 a_60964_12612# a_61412_12612# 0.01328f
C16211 _260_.A2 _448_.Q 0.01414f
C16212 _386_.A4 a_47476_28292# 0.00193f
C16213 _332_.Z a_41572_18504# 0.01909f
C16214 a_41116_26247# _451_.Q 0.00284f
C16215 a_42168_22504# a_43600_22504# 0.01212f
C16216 a_67012_9096# VPWR 0.20348f
C16217 a_65556_23588# a_65196_23544# 0.08674f
C16218 a_49316_11044# a_48956_11000# 0.08707f
C16219 a_61524_12232# a_61412_11044# 0.02666f
C16220 a_2724_18504# VPWR 0.20782f
C16221 _324_.C vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN 0.01417f
C16222 _245_.Z clk 0.00353f
C16223 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN 0.76304f
C16224 _256_.A2 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I 0.05283f
C16225 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN VPWR 0.81502f
C16226 a_67236_1636# a_67100_1159# 0.00168f
C16227 a_30812_1159# a_31484_1159# 0.00544f
C16228 _330_.ZN a_37084_17272# 0.00118f
C16229 a_28928_29123# uo_out[7] 0.00484f
C16230 a_61524_10664# a_61972_10664# 0.01328f
C16231 _362_.B _359_.ZN 0.00849f
C16232 a_28036_2824# a_28036_1636# 0.05841f
C16233 a_23556_24776# a_23644_23111# 0.00151f
C16234 _371_.A3 _336_.Z 0.12149f
C16235 a_33152_22091# VPWR 1.13484f
C16236 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I a_55700_25156# 0.0016f
C16237 _349_.A4 a_24952_29032# 0.42096f
C16238 _416_.A1 a_38628_25156# 0.01454f
C16239 a_35728_29480# a_36656_29123# 1.16391f
C16240 a_1916_12568# VPWR 0.297f
C16241 a_33188_21640# a_33636_21640# 0.01328f
C16242 a_53212_2727# VPWR 0.31143f
C16243 a_62620_18407# a_62980_18504# 0.08717f
C16244 a_17932_26247# a_17844_26344# 0.28563f
C16245 _452_.CLK a_38523_27967# 0.00219f
C16246 a_34980_15368# a_35428_15368# 0.01328f
C16247 a_23108_29860# VPWR 0.12051f
C16248 _460_.Q a_35292_26247# 0.02828f
C16249 a_54220_10567# VPWR 0.31547f
C16250 a_40220_26247# _261_.ZN 0.00329f
C16251 a_36860_15271# a_36772_15368# 0.28563f
C16252 a_16052_23208# VPWR 0.20348f
C16253 a_31920_29480# a_32800_29167# 0.00306f
C16254 a_38428_15271# a_38876_15271# 0.0131f
C16255 _268_.A2 a_52292_29480# 0.00652f
C16256 a_50084_24328# clk 0.0245f
C16257 a_43444_19668# a_43668_19668# 0.01436f
C16258 a_48776_20204# a_49448_20072# 0.00478f
C16259 a_2724_28292# a_2812_28248# 0.28563f
C16260 _402_.ZN VPWR 0.37259f
C16261 a_1020_21976# a_1468_21976# 0.0131f
C16262 a_50972_2727# a_50884_2824# 0.28563f
C16263 a_3620_22020# a_3260_21976# 0.08717f
C16264 a_62620_17272# a_63068_17272# 0.0131f
C16265 a_67012_17316# a_66652_17272# 0.0869f
C16266 a_66652_7431# a_67100_7431# 0.0131f
C16267 a_22996_23588# a_23444_23588# 0.01328f
C16268 a_65756_8999# a_66204_8999# 0.0131f
C16269 a_31844_1256# a_32292_1256# 0.01328f
C16270 a_61860_30736# ui_in[3] 0.00378f
C16271 a_15156_25156# a_14796_25112# 0.08707f
C16272 a_46716_13703# a_47076_13800# 0.08717f
C16273 a_60716_13703# a_61164_13703# 0.01288f
C16274 a_51196_14136# a_51108_12612# 0.00151f
C16275 a_10876_2727# a_11324_2727# 0.0131f
C16276 a_1468_18840# a_1468_18407# 0.05841f
C16277 _474_.CLK a_52884_18884# 0.00132f
C16278 _229_.I _252_.ZN 0.06167f
C16279 a_54692_20452# a_54780_20408# 0.28563f
C16280 _324_.C _381_.A2 0.91159f
C16281 a_33500_16839# a_33860_16936# 0.08717f
C16282 _465_.D a_19248_29977# 0.00167f
C16283 a_3172_10664# a_3172_9476# 0.05841f
C16284 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I VPWR 1.23485f
C16285 a_22548_29480# uio_out[4] 0.00311f
C16286 a_29828_1636# VPWR 0.20348f
C16287 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN a_64860_19975# 0.00584f
C16288 a_14908_30951# a_15460_31048# 0.01375f
C16289 _419_.A4 a_47271_21640# 0.02001f
C16290 a_54556_12568# a_54668_12135# 0.02634f
C16291 a_58500_12612# a_58476_12135# 0.00172f
C16292 _402_.A1 _424_.A2 0.34306f
C16293 a_65220_18504# a_66004_18504# 0.00276f
C16294 a_65756_26247# a_65668_26344# 0.28563f
C16295 a_55812_11044# a_56260_11044# 0.01328f
C16296 a_4068_15368# a_4068_14180# 0.05841f
C16297 _398_.C _402_.B 0.05171f
C16298 a_13788_1592# a_13788_1159# 0.05841f
C16299 a_41564_1592# a_42012_1592# 0.01288f
C16300 a_45508_1636# a_45596_1592# 0.28563f
C16301 a_46964_16936# a_47412_16936# 0.01328f
C16302 a_63180_26680# vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN 0.03293f
C16303 _267_.A2 a_59348_29076# 0.00571f
C16304 _411_.A2 a_49172_27508# 0.00718f
C16305 a_54444_23544# VPWR 0.29714f
C16306 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_57168_26724# 0.00528f
C16307 _246_.B2 a_60740_26724# 0.00103f
C16308 _452_.Q _331_.ZN 0.01069f
C16309 a_51240_23340# _475_.Q 0.02416f
C16310 a_54892_24679# a_55252_24776# 0.08674f
C16311 a_16588_20408# VPWR 0.31143f
C16312 a_48308_23588# _324_.B 0.00268f
C16313 _474_.CLK a_52900_26724# 0.00345f
C16314 a_55364_12612# VPWR 0.20595f
C16315 _352_.A2 _337_.ZN 0.59561f
C16316 a_11684_2824# a_12356_2824# 0.00347f
C16317 _251_.A1 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN 0.66038f
C16318 a_19328_28733# a_18096_27165# 0.00141f
C16319 a_9532_29383# a_9892_29480# 0.08717f
C16320 a_31484_30951# _370_.B 0.00629f
C16321 _444_.D a_36048_24831# 0.00247f
C16322 a_30812_15704# a_30812_15271# 0.05841f
C16323 a_34756_15748# a_34620_15271# 0.00168f
C16324 a_24864_29931# a_25792_30301# 1.16391f
C16325 a_19372_30345# a_19716_29977# 0.00275f
C16326 a_47972_10664# VPWR 0.20348f
C16327 a_24876_21976# a_24900_21640# 0.00172f
C16328 a_47836_15271# a_48196_15368# 0.08717f
C16329 a_56148_23588# VPWR 0.20348f
C16330 a_36996_26724# a_36636_26680# 0.0869f
C16331 _260_.A1 a_42460_20452# 0.0013f
C16332 _371_.A2 _371_.A1 0.23966f
C16333 _334_.A1 a_33720_28776# 0.00128f
C16334 a_63516_15271# VPWR 0.29679f
C16335 a_19328_28733# a_17472_28363# 0.02366f
C16336 a_19035_28409# _378_.ZN 0.03473f
C16337 a_17396_22020# a_17036_21976# 0.08707f
C16338 a_67100_15704# VPWR 0.32971f
C16339 a_26556_27815# VPWR 0.32202f
C16340 a_61948_2727# a_62308_2824# 0.08717f
C16341 a_46044_30951# a_46628_31048# 0.01675f
C16342 a_58388_17316# a_58252_16839# 0.00168f
C16343 a_65444_15368# a_65892_15368# 0.01328f
C16344 a_38340_21327# a_38548_21327# 0.00334f
C16345 a_58164_18504# vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I 0.00122f
C16346 uio_out[0] uo_out[7] 0.06783f
C16347 a_17956_1256# VPWR 0.2067f
C16348 a_66116_7908# VPWR 0.23643f
C16349 a_67908_4772# VPWR 0.21437f
C16350 a_21516_25112# a_21964_25112# 0.012f
C16351 a_8636_29383# VPWR 0.33315f
C16352 a_58028_13703# a_57940_13800# 0.28563f
C16353 a_35504_18955# a_35628_18407# 0.00156f
C16354 _355_.B a_28891_25273# 0.00261f
C16355 a_53908_16936# a_54108_15271# 0.00119f
C16356 a_44812_16839# a_44724_16936# 0.28563f
C16357 VPWR uio_in[2] 0.00217f
C16358 _267_.A2 a_52756_29076# 0.03685f
C16359 a_43492_27912# a_43564_27209# 0.00175f
C16360 a_43940_27912# a_43936_27165# 0.00375f
C16361 a_44388_27912# a_43008_26795# 0.00999f
C16362 _324_.C a_51988_24072# 0.00491f
C16363 a_35964_1592# VPWR 0.3289f
C16364 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN a_55900_15271# 0.001f
C16365 a_3260_1159# a_3620_1256# 0.08717f
C16366 a_33412_16936# VPWR 0.20644f
C16367 a_4604_1592# a_5052_1592# 0.01288f
C16368 a_36836_20072# VPWR 0.00667f
C16369 a_65444_12612# a_65420_12135# 0.00172f
C16370 a_47612_12135# a_48060_12135# 0.0131f
C16371 _424_.A2 a_52081_21236# 0.0023f
C16372 _437_.A1 a_37196_23544# 0.00184f
C16373 a_16140_25112# a_16140_24679# 0.05841f
C16374 a_20084_25156# a_20060_24679# 0.00172f
C16375 a_3620_29860# a_3260_29816# 0.08707f
C16376 a_65780_12232# a_65868_10567# 0.00151f
C16377 a_44700_30951# VPWR 0.31143f
C16378 a_45284_15368# a_45284_14180# 0.05841f
C16379 a_40040_17675# a_40916_16936# 0.00102f
C16380 a_48868_1636# a_48508_1592# 0.08707f
C16381 _452_.D a_42896_18504# 0.00114f
C16382 _416_.A1 a_46476_20937# 0.06383f
C16383 _421_.A1 _419_.Z 0.05606f
C16384 a_46940_15271# a_47076_14180# 0.00154f
C16385 a_1020_24679# a_1468_24679# 0.0131f
C16386 a_48060_18407# a_48420_18504# 0.08717f
C16387 a_53212_1159# a_53660_1159# 0.0131f
C16388 a_17396_27912# a_16796_27209# 0.01033f
C16389 a_39684_20072# a_40132_20072# 0.01328f
C16390 a_66564_18884# a_66652_18840# 0.28563f
C16391 a_62172_18840# a_62620_18840# 0.0131f
C16392 a_16052_25156# VPWR 0.20348f
C16393 a_27564_20408# VPWR 0.31712f
C16394 a_15692_27815# a_15604_27912# 0.28563f
C16395 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN 0.03353f
C16396 a_30724_15748# a_31172_15748# 0.01328f
C16397 a_61948_12568# VPWR 0.31389f
C16398 a_19860_26724# uio_out[7] 0.03469f
C16399 vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I a_66228_20452# 0.00125f
C16400 a_41700_15748# a_41564_15271# 0.00168f
C16401 a_52360_26355# a_53772_26031# 0.00393f
C16402 _260_.A1 a_41664_22020# 0.00293f
C16403 a_36524_16839# a_36548_15748# 0.0016f
C16404 a_63988_16936# VPWR 0.20703f
C16405 a_58140_26680# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.02997f
C16406 _304_.B a_46068_25156# 0.00491f
C16407 a_23834_28292# VPWR 0.01449f
C16408 _274_.A1 a_56572_29383# 0.0056f
C16409 a_43492_15368# VPWR 0.20348f
C16410 _378_.ZN uio_out[7] 0.36081f
C16411 a_23892_22020# a_24340_22020# 0.01328f
C16412 a_46940_15271# VPWR 0.29679f
C16413 _294_.A2 _365_.ZN 0.95788f
C16414 a_41900_16839# a_42572_16839# 0.00544f
C16415 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN 0.14852f
C16416 a_3260_16839# VPWR 0.30487f
C16417 a_63764_23208# vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN 0.03524f
C16418 a_40356_1256# VPWR 0.20348f
C16419 a_54244_1256# a_54692_1256# 0.01328f
C16420 a_33276_2727# a_33724_2727# 0.0131f
C16421 a_54580_13800# a_55028_13800# 0.01328f
C16422 a_52428_13703# a_52452_12612# 0.0016f
C16423 _350_.A1 uo_out[6] 0.44833f
C16424 a_37532_17272# a_37420_16839# 0.02634f
C16425 _474_.CLK a_56236_23544# 0.01027f
C16426 a_1916_17272# VPWR 0.297f
C16427 _433_.ZN _441_.A2 0.36288f
C16428 a_14684_1159# a_14596_1256# 0.28563f
C16429 a_57380_16936# VPWR 0.15769f
C16430 vgaringosc.workerclkbuff_notouch_.I a_45012_29816# 0.03232f
C16431 a_57044_10664# a_57156_9476# 0.02666f
C16432 a_49764_1636# VPWR 0.20967f
C16433 a_5388_12135# a_5300_12232# 0.28563f
C16434 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN 0.00109f
C16435 a_11908_1636# a_11548_1592# 0.08707f
C16436 a_56684_18407# VPWR 0.33321f
C16437 a_10116_29860# a_10564_29860# 0.01328f
C16438 _386_.ZN a_47600_27912# 0.00835f
C16439 a_32604_17272# a_33052_17272# 0.01288f
C16440 a_36548_17316# a_36636_17272# 0.28563f
C16441 a_20420_2824# VPWR 0.20815f
C16442 a_55228_1592# a_55812_1636# 0.01675f
C16443 _459_.CLK a_20308_26724# 0.02152f
C16444 _459_.Q a_32380_26247# 0.04833f
C16445 a_66340_11044# a_65980_11000# 0.08707f
C16446 a_62396_11000# a_62844_11000# 0.01288f
C16447 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62644_26724# 0.01276f
C16448 a_53908_24776# VPWR 0.20524f
C16449 _416_.A1 _437_.A1 0.12052f
C16450 a_20956_23111# a_21404_23111# 0.01288f
C16451 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN 0.00244f
C16452 a_3260_24679# a_3620_24776# 0.08717f
C16453 _311_.A2 _448_.Q 0.00342f
C16454 a_52900_26724# a_52988_26680# 0.28563f
C16455 a_62732_26680# _245_.I1 0.00505f
C16456 a_1916_14136# VPWR 0.297f
C16457 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I a_56404_27208# 0.00162f
C16458 _434_.ZN a_39536_23588# 0.00175f
C16459 _230_.I _243_.ZN 0.10618f
C16460 a_4740_2824# a_4828_1159# 0.0027f
C16461 a_22188_29383# a_22100_29480# 0.28563f
C16462 a_56596_29861# VPWR 0.54333f
C16463 _352_.A2 a_27924_24776# 0.00978f
C16464 _448_.Q a_37067_19001# 0.00931f
C16465 a_37892_15748# a_37532_15704# 0.08663f
C16466 a_56012_12135# VPWR 0.31547f
C16467 a_5188_29480# VPWR 0.20885f
C16468 a_34084_2824# a_34532_2824# 0.01328f
C16469 a_41922_31073# VPWR 0.01259f
C16470 _358_.A3 a_36188_26247# 0.00572f
C16471 _352_.ZN a_27140_26344# 0.07238f
C16472 a_18716_24679# VPWR 0.32683f
C16473 a_44744_26355# _402_.ZN 0.27276f
C16474 a_58116_30344# a_57220_29861# 0.00915f
C16475 _255_.I a_59744_30352# 0.00188f
C16476 _399_.A2 a_48908_24080# 0.00593f
C16477 _281_.ZN _279_.Z 0.07208f
C16478 a_24452_21640# a_24564_20452# 0.02666f
C16479 a_43468_16839# a_43492_15748# 0.0016f
C16480 a_46068_25156# VPWR 0.22618f
C16481 a_33476_27912# VPWR 0.0154f
C16482 a_31260_15704# VPWR 0.29679f
C16483 _350_.A1 uo_out[5] 0.12131f
C16484 _324_.C a_56484_29480# 0.00569f
C16485 _424_.B1 _424_.A2 2.16362f
C16486 _337_.ZN _223_.ZN 0.0468f
C16487 _381_.Z a_48596_28292# 0.00131f
C16488 _304_.B _384_.ZN 0.02446f
C16489 a_1468_9432# a_1916_9432# 0.0131f
C16490 a_4068_9476# a_3708_9432# 0.08717f
C16491 a_11548_30951# uio_oe[3] 0.00925f
C16492 _452_.CLK _319_.A2 0.30992f
C16493 a_47164_14136# a_47612_14136# 0.01288f
C16494 a_51108_14180# a_51196_14136# 0.28563f
C16495 _452_.CLK a_41536_17636# 0.00895f
C16496 a_46716_18407# VPWR 0.32774f
C16497 a_19035_28409# uio_out[6] 0.00473f
C16498 a_50412_16839# VPWR 0.364f
C16499 a_62756_1256# VPWR 0.20348f
C16500 _384_.A1 a_53300_23047# 0.00864f
C16501 a_59372_13703# a_59396_12612# 0.0016f
C16502 a_55588_28292# a_55676_28248# 0.28563f
C16503 _475_.Q a_52434_22504# 0.007f
C16504 a_38228_20452# VPWR 0.12615f
C16505 _452_.CLK _325_.B 0.35968f
C16506 a_44724_17316# VPWR 0.20692f
C16507 a_55900_1592# VPWR 0.33352f
C16508 a_64212_10664# a_64324_9476# 0.02666f
C16509 a_25660_1159# a_26020_1256# 0.08717f
C16510 a_55564_12135# a_55924_12232# 0.08707f
C16511 a_53212_12568# a_53124_11044# 0.00151f
C16512 _412_.B2 _412_.ZN 0.00113f
C16513 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_55956_25940# 0.0893f
C16514 a_1828_12232# a_2276_12232# 0.01328f
C16515 a_18404_1636# a_18852_1636# 0.01328f
C16516 _448_.Q a_37444_21640# 0.00956f
C16517 a_2364_21543# VPWR 0.30029f
C16518 _452_.Q a_39324_19975# 0.00592f
C16519 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I 0.00372f
C16520 a_41048_17341# a_41968_17801# 0.00306f
C16521 a_44724_17316# a_44364_17272# 0.0869f
C16522 a_9308_29816# uio_oe[5] 0.00276f
C16523 _336_.A2 a_30388_23588# 0.00154f
C16524 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I a_56404_27208# 0.04325f
C16525 a_56036_27912# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.00383f
C16526 _230_.I a_58140_26680# 0.00338f
C16527 a_42820_2824# VPWR 0.2556f
C16528 a_62532_1636# a_62172_1592# 0.08707f
C16529 _397_.A2 a_47172_23588# 0.0039f
C16530 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I 0.82576f
C16531 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN 0.06152f
C16532 a_14708_24776# a_15156_24776# 0.01328f
C16533 a_20060_23111# a_19972_23208# 0.28563f
C16534 a_23644_24679# a_23556_24776# 0.28563f
C16535 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN a_59260_21976# 0.0046f
C16536 a_45820_9432# VPWR 0.31143f
C16537 a_60604_27815# a_60964_27912# 0.0869f
C16538 a_55364_14180# VPWR 0.20348f
C16539 a_36076_18407# a_36436_18504# 0.08663f
C16540 _393_.ZN a_46772_29977# 0.00247f
C16541 a_4740_31048# a_4604_29816# 0.00154f
C16542 _371_.ZN _350_.A2 0.01839f
C16543 _350_.A1 _373_.A2 0.59677f
C16544 a_50100_12232# VPWR 0.21427f
C16545 a_40804_15748# a_40892_15704# 0.28563f
C16546 a_44388_15748# a_44836_15748# 0.01328f
C16547 _316_.A3 a_36996_21640# 0.00641f
C16548 _421_.A1 _416_.A2 0.25827f
C16549 a_23108_24776# VPWR 0.20622f
C16550 _470_.Q _284_.A2 0.33648f
C16551 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_55252_26724# 0.00202f
C16552 vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN 0.01026f
C16553 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN 0.0386f
C16554 a_54824_22045# a_55312_22340# 0.8399f
C16555 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I a_55900_15271# 0.00473f
C16556 _261_.ZN _441_.A2 0.11098f
C16557 a_31844_21640# a_31732_20452# 0.02666f
C16558 a_30052_21640# a_30028_20408# 0.0016f
C16559 a_5724_2727# a_6084_2824# 0.08717f
C16560 a_50412_16839# a_50436_15748# 0.0016f
C16561 _442_.ZN _436_.ZN 0.10835f
C16562 _231_.ZN a_59397_26344# 0.04055f
C16563 a_32604_19975# a_32516_20072# 0.28563f
C16564 a_44924_15704# VPWR 0.29679f
C16565 _384_.ZN VPWR 0.83772f
C16566 _384_.A3 a_51220_22504# 0.01223f
C16567 a_41476_26344# _260_.A2 0.00392f
C16568 a_66540_19975# VPWR 0.33132f
C16569 a_1916_14136# a_1916_13703# 0.05841f
C16570 _459_.Q _336_.Z 1.21488f
C16571 a_54916_14180# a_54556_14136# 0.08717f
C16572 _452_.CLK a_40220_26247# 0.00716f
C16573 _444_.D _437_.ZN 0.00575f
C16574 uio_out[6] uio_out[7] 0.03426f
C16575 _358_.A3 a_33188_25940# 0.51374f
C16576 a_66316_13703# a_66340_12612# 0.0016f
C16577 a_4156_12568# a_4604_12568# 0.01222f
C16578 a_56372_13800# a_56260_12612# 0.02666f
C16579 a_55676_2727# a_56124_2727# 0.0131f
C16580 _424_.A2 a_52676_17316# 0.00155f
C16581 _474_.CLK a_55700_24776# 0.0497f
C16582 a_37980_26247# VPWR 0.34108f
C16583 a_52764_17272# VPWR 0.31547f
C16584 a_20191_29611# VPWR 0.00615f
C16585 a_17803_26841# a_18292_25156# 0.00225f
C16586 _327_.A2 a_46268_18407# 0.00133f
C16587 a_37084_1159# a_36996_1256# 0.28563f
C16588 a_1828_9096# a_1828_7908# 0.05841f
C16589 a_2724_7528# a_2724_6340# 0.05841f
C16590 a_5724_1159# VPWR 0.3289f
C16591 a_66764_12135# a_66676_12232# 0.28563f
C16592 a_3620_5960# a_3620_4772# 0.05841f
C16593 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN _248_.B1 0.00488f
C16594 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN 0.00789f
C16595 _451_.Q a_40668_19975# 0.01696f
C16596 a_33276_21543# VPWR 0.33094f
C16597 a_21052_26031# a_21428_25156# 0.00189f
C16598 a_52228_17316# a_52676_17316# 0.01328f
C16599 VPWR uo_out[4] 0.8734f
C16600 a_48644_17316# a_48732_17272# 0.28563f
C16601 a_64996_2824# VPWR 0.21436f
C16602 a_2812_10567# a_3172_10664# 0.08717f
C16603 a_56460_10567# a_57132_10567# 0.00544f
C16604 a_64636_1592# a_65084_1592# 0.0131f
C16605 a_67236_1636# a_66876_1592# 0.08674f
C16606 a_27228_26680# a_27228_26247# 0.05841f
C16607 _287_.A1 _459_.CLK 0.05459f
C16608 _438_.A2 a_39780_22805# 0.0196f
C16609 a_30588_23111# a_30948_23208# 0.08707f
C16610 _452_.CLK a_33520_25597# 0.00207f
C16611 a_18628_23208# a_19076_23208# 0.01328f
C16612 _388_.B a_44632_30206# 0.21723f
C16613 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I 0.00456f
C16614 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.05753f
C16615 a_1828_6340# VPWR 0.20348f
C16616 _455_.Q a_25232_27165# 0.01104f
C16617 a_1828_23588# VPWR 0.20348f
C16618 a_56796_9432# VPWR 0.31959f
C16619 a_63740_14136# VPWR 0.31389f
C16620 _399_.ZN a_47860_23208# 0.00397f
C16621 a_3708_21543# a_3620_21640# 0.28563f
C16622 a_3620_3204# VPWR 0.22347f
C16623 a_932_29480# a_932_28292# 0.05841f
C16624 a_24988_21543# a_25436_21543# 0.01288f
C16625 a_26916_2824# a_27004_1159# 0.0027f
C16626 a_63204_2824# a_63068_1592# 0.00154f
C16627 _424_.A2 _218_.ZN 0.09314f
C16628 _238_.ZN a_59572_29076# 0.07656f
C16629 _459_.CLK a_31932_26247# 0.04768f
C16630 a_38523_27967# a_38816_27555# 0.49319f
C16631 a_13364_31048# a_13340_29816# 0.0016f
C16632 _451_.Q _447_.Q 0.11827f
C16633 a_28228_25273# VPWR 0.00246f
C16634 a_4068_11044# VPWR 0.2157f
C16635 a_56484_2824# a_56932_2824# 0.01328f
C16636 _284_.A2 _260_.A2 0.00112f
C16637 a_49068_20408# VPWR 0.8101f
C16638 _284_.ZN _265_.ZN 0.07776f
C16639 a_63516_19975# a_63876_20072# 0.08717f
C16640 a_66652_18840# a_66540_18407# 0.02634f
C16641 a_52756_29076# vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.00127f
C16642 _383_.A2 a_48596_28292# 0.0122f
C16643 _428_.Z a_52452_24072# 0.02414f
C16644 _340_.A2 uio_out[0] 0.09955f
C16645 _313_.ZN a_34980_22895# 0.01057f
C16646 a_5052_18840# VPWR 0.33516f
C16647 _294_.ZN _371_.A1 0.1115f
C16648 _359_.B a_40264_30320# 0.00895f
C16649 _268_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I 0.04907f
C16650 a_59828_26724# VPWR 0.00636f
C16651 a_62284_26680# a_62732_26680# 0.01255f
C16652 a_17148_2727# a_17060_2824# 0.28563f
C16653 _416_.A1 a_51050_29480# 0.00593f
C16654 a_53460_24776# a_52920_22760# 0.00159f
C16655 a_54244_9476# a_53884_9432# 0.08717f
C16656 _274_.ZN _274_.A2 0.01643f
C16657 a_55588_9476# a_56036_9476# 0.01328f
C16658 a_62756_14180# a_63204_14180# 0.01328f
C16659 a_52452_14180# a_52428_13703# 0.00172f
C16660 a_48508_14136# a_48508_13703# 0.05841f
C16661 a_4964_20452# a_5052_20408# 0.28563f
C16662 _330_.ZN a_37964_18191# 0.22165f
C16663 a_37408_18504# a_38971_18559# 0.41635f
C16664 a_51108_12612# a_50748_12568# 0.08707f
C16665 _334_.A1 a_33483_29535# 0.03776f
C16666 _452_.CLK a_32740_21640# 0.00484f
C16667 a_63316_13800# a_63204_12612# 0.02666f
C16668 _438_.ZN a_40780_21543# 0.00362f
C16669 _384_.ZN _383_.ZN 0.04134f
C16670 _293_.A2 _459_.CLK 0.07964f
C16671 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN 0.00957f
C16672 _335_.ZN a_34084_28776# 1.66144f
C16673 a_17396_24776# a_17396_23588# 0.05841f
C16674 _452_.Q a_40132_20452# 0.04745f
C16675 a_22064_27912# a_22992_27555# 1.16391f
C16676 a_28124_1159# VPWR 0.29679f
C16677 _330_.A1 _403_.ZN 0.21653f
C16678 a_63316_12232# a_63764_12232# 0.01328f
C16679 a_48060_1159# a_48420_1256# 0.08717f
C16680 a_24540_1592# a_24988_1592# 0.01288f
C16681 a_28484_1636# a_28572_1592# 0.28563f
C16682 _257_.B _238_.ZN 0.3069f
C16683 _381_.A2 a_50724_24908# 0.00599f
C16684 a_30500_21640# VPWR 0.20692f
C16685 a_37084_26247# a_36996_26344# 0.28563f
C16686 a_38472_30169# a_37584_29123# 0.01356f
C16687 a_52900_1636# a_52764_1159# 0.00168f
C16688 a_48956_1592# a_48956_1159# 0.05841f
C16689 _275_.ZN _408_.ZN 0.00478f
C16690 a_53772_10567# a_53684_10664# 0.28563f
C16691 _438_.A2 a_39796_22504# 0.04047f
C16692 a_48776_20204# VPWR 0.29059f
C16693 a_13700_2824# a_13700_1636# 0.05841f
C16694 a_9892_2824# a_9756_1592# 0.00154f
C16695 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN 0.01409f
C16696 _247_.B _245_.Z 0.09978f
C16697 a_2724_22020# VPWR 0.20782f
C16698 a_20172_23544# VPWR 0.31547f
C16699 a_4156_8999# VPWR 0.3269f
C16700 a_58028_13703# VPWR 0.35236f
C16701 _270_.A2 ui_in[4] 0.00915f
C16702 a_1380_18884# a_1828_18884# 0.01328f
C16703 a_23644_21543# a_24004_21640# 0.08707f
C16704 a_7964_2727# VPWR 0.33981f
C16705 a_64860_5863# VPWR 0.30145f
C16706 _334_.A1 a_35140_26680# 0.00162f
C16707 _397_.Z clk 0.02671f
C16708 _459_.CLK a_28000_29480# 0.05639f
C16709 a_51791_30644# uio_in[0] 0.48586f
C16710 _351_.ZN a_24736_26841# 0.00242f
C16711 a_50524_15704# a_50972_15704# 0.01288f
C16712 a_17956_29860# _379_.Z 0.00564f
C16713 a_53124_11044# VPWR 0.2267f
C16714 a_44744_26355# a_46068_25156# 0.00179f
C16715 _325_.B a_43668_19668# 0.90178f
C16716 _474_.CLK _424_.ZN 0.04834f
C16717 a_4156_26680# VPWR 0.30552f
C16718 a_56684_23544# a_57132_23544# 0.0131f
C16719 a_62084_15748# a_62172_15704# 0.28563f
C16720 a_10092_30951# uio_oe[5] 0.00326f
C16721 a_28036_26724# a_27676_26680# 0.08663f
C16722 _436_.ZN _435_.ZN 0.38234f
C16723 _390_.ZN _404_.A1 0.0054f
C16724 a_21052_26031# VPWR 0.39897f
C16725 a_28124_2727# a_28484_2824# 0.08717f
C16726 a_2276_23588# a_2364_23544# 0.28563f
C16727 a_15244_28248# VPWR 0.29679f
C16728 a_2276_6340# a_2364_6296# 0.28563f
C16729 a_1380_7908# a_1468_7864# 0.28563f
C16730 a_3172_4772# a_3260_4728# 0.28563f
C16731 a_55900_14136# a_56012_13703# 0.02634f
C16732 a_4068_3204# a_4156_3160# 0.28563f
C16733 a_18964_20452# a_19412_20452# 0.01328f
C16734 _427_.B1 a_52660_21640# 0.00703f
C16735 _252_.B _247_.B 0.976f
C16736 a_52764_27815# a_53212_27815# 0.01255f
C16737 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_53996_26680# 0.0016f
C16738 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN a_57580_23544# 0.00799f
C16739 a_57492_23588# _231_.I 0.00493f
C16740 a_1916_1592# VPWR 0.297f
C16741 a_61860_30736# _256_.A2 0.002f
C16742 a_54020_12612# a_54108_12568# 0.28563f
C16743 a_57604_12612# a_58052_12612# 0.01328f
C16744 a_39748_29480# uo_out[1] 0.01799f
C16745 _459_.CLK a_20084_25156# 0.01384f
C16746 _287_.A1 uo_out[7] 0.02916f
C16747 _290_.ZN uo_out[6] 0.00129f
C16748 a_24452_24776# a_24340_23588# 0.02666f
C16749 a_59484_1159# a_59396_1256# 0.28563f
C16750 a_50524_1159# VPWR 0.37175f
C16751 a_4516_11044# a_4604_11000# 0.28563f
C16752 a_67908_18884# VPWR 0.21212f
C16753 a_32592_25227# a_34155_25273# 0.41635f
C16754 _363_.Z a_30388_28776# 0.0209f
C16755 a_41228_27815# a_42148_27912# 0.00795f
C16756 a_50548_10664# a_50996_10664# 0.01328f
C16757 _311_.A2 a_36172_24463# 0.00532f
C16758 a_64300_10567# a_64884_10664# 0.01675f
C16759 a_35628_18407# a_35652_17316# 0.0016f
C16760 a_19388_1159# a_20060_1159# 0.00544f
C16761 _355_.C a_22064_27912# 0.03617f
C16762 _474_.CLK vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN 0.00376f
C16763 a_21068_21976# VPWR 0.31589f
C16764 a_22212_21640# a_22660_21640# 0.01328f
C16765 a_31172_18884# a_30812_18840# 0.08717f
C16766 a_30364_2727# VPWR 0.31143f
C16767 a_51892_13800# VPWR 0.20595f
C16768 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN 0.00966f
C16769 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN 0.05849f
C16770 a_65980_15271# a_66428_15271# 0.01255f
C16771 _327_.Z a_40416_18885# 0.19464f
C16772 a_7292_29816# VPWR 0.3289f
C16773 a_52415_31220# ui_in[7] 0.00947f
C16774 a_66788_11044# VPWR 0.20622f
C16775 a_19276_21976# a_19164_21543# 0.02634f
C16776 a_17932_23111# VPWR 0.32173f
C16777 _359_.B _359_.ZN 0.14367f
C16778 _247_.ZN a_60068_27912# 0.00488f
C16779 a_1916_15271# a_2364_15271# 0.0131f
C16780 a_19412_27912# VPWR 0.2461f
C16781 _437_.A1 _431_.A3 0.58934f
C16782 _304_.B a_51576_25896# 0.0037f
C16783 a_63964_17272# a_63876_15748# 0.00151f
C16784 a_61076_23208# a_61524_23208# 0.01328f
C16785 _260_.A1 _450_.D 0.00218f
C16786 a_39548_2727# a_39460_2824# 0.28563f
C16787 _290_.ZN uo_out[5] 1.9187f
C16788 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I VPWR 0.73114f
C16789 a_61388_16839# a_61748_16936# 0.08717f
C16790 _255_.ZN _243_.A1 0.01862f
C16791 a_65220_9476# a_64860_9432# 0.08717f
C16792 a_66564_9476# a_67012_9476# 0.01328f
C16793 a_58388_20452# vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.00155f
C16794 a_19636_23588# a_20084_23588# 0.01328f
C16795 a_16052_23588# a_16140_23544# 0.28563f
C16796 a_932_25156# a_1020_25112# 0.28563f
C16797 a_65308_6296# a_65756_6296# 0.0131f
C16798 a_67460_6340# a_67548_6296# 0.28563f
C16799 a_64412_7864# a_64860_7864# 0.0131f
C16800 a_66564_7908# a_66652_7864# 0.28563f
C16801 a_20420_1256# a_20868_1256# 0.01328f
C16802 a_39300_31048# uo_out[3] 0.00247f
C16803 _293_.A2 uo_out[7] 0.01448f
C16804 a_54780_18840# VPWR 0.3272f
C16805 a_66204_4728# a_66652_4728# 0.0131f
C16806 _246_.B2 ui_in[2] 0.02814f
C16807 a_67236_14180# a_67212_13703# 0.00172f
C16808 a_24564_20452# a_24652_20408# 0.28563f
C16809 a_67100_3160# a_67548_3160# 0.0131f
C16810 a_49740_13703# a_50188_13703# 0.01288f
C16811 a_14460_30951# a_14372_31048# 0.28563f
C16812 a_10876_29383# a_11324_29383# 0.0131f
C16813 a_64860_17272# a_64972_16839# 0.02634f
C16814 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN a_60852_15748# 0.0356f
C16815 a_40692_21640# a_40668_20408# 0.0016f
C16816 a_67572_13800# a_67660_12135# 0.00151f
C16817 a_15580_1592# VPWR 0.29679f
C16818 a_2364_30951# a_2812_30951# 0.0131f
C16819 a_23920_27555# _351_.A2 0.00237f
C16820 _421_.A1 _399_.ZN 0.02834f
C16821 _268_.A2 vgaringosc.workerclkbuff_notouch_.I 0.04485f
C16822 _386_.A4 a_46804_28292# 0.00123f
C16823 a_16028_29816# a_16164_29480# 0.00168f
C16824 a_66452_18504# a_66540_16839# 0.00151f
C16825 a_42168_22504# a_43192_22504# 0.00951f
C16826 a_66564_9096# VPWR 0.20631f
C16827 a_65108_23588# a_65196_23544# 0.28563f
C16828 a_48868_11044# a_48956_11000# 0.28563f
C16829 a_35988_16936# a_36436_16936# 0.01328f
C16830 a_2276_18504# VPWR 0.20634f
C16831 a_38204_1592# a_38652_1592# 0.01288f
C16832 _336_.A2 a_24080_25227# 0.00124f
C16833 _324_.C a_64412_29816# 0.00308f
C16834 a_40220_19975# a_40668_19975# 0.012f
C16835 _268_.A2 a_53124_27912# 0.00169f
C16836 a_28000_29480# uo_out[7] 0.01091f
C16837 a_64636_1592# a_64636_1159# 0.05841f
C16838 _256_.A2 a_64324_29860# 0.0038f
C16839 _457_.D a_24512_25273# 0.00165f
C16840 a_44795_29535# a_45040_29167# 0.00232f
C16841 _436_.ZN _441_.ZN 0.7188f
C16842 a_5052_26680# a_4940_26247# 0.02634f
C16843 a_38644_19368# _330_.A2 0.38386f
C16844 a_47164_30951# a_47612_30951# 0.0131f
C16845 a_52764_2727# VPWR 0.31143f
C16846 a_1468_12568# VPWR 0.29679f
C16847 a_62620_18407# a_62532_18504# 0.28563f
C16848 a_17484_26247# a_17844_26344# 0.08717f
C16849 a_66452_16936# a_66428_15271# 0.00134f
C16850 a_3172_26344# a_3620_26344# 0.01328f
C16851 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I 0.72819f
C16852 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I 0.00228f
C16853 _452_.CLK a_37516_27599# 0.00996f
C16854 a_22560_30288# VPWR 0.4471f
C16855 a_53772_10567# VPWR 0.31547f
C16856 _460_.Q a_33396_26344# 0.00329f
C16857 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I VPWR 0.7394f
C16858 a_36412_15271# a_36772_15368# 0.08717f
C16859 a_15604_23208# VPWR 0.20348f
C16860 _268_.A2 a_52068_29480# 0.01847f
C16861 a_38336_18147# a_38316_16839# 0.00148f
C16862 a_4516_28292# a_4964_28292# 0.01328f
C16863 a_2724_28292# a_2364_28248# 0.08717f
C16864 a_51576_25896# VPWR 0.51401f
C16865 a_50524_2727# a_50884_2824# 0.08717f
C16866 a_3172_22020# a_3260_21976# 0.28563f
C16867 _435_.ZN _439_.ZN 0.01944f
C16868 a_66564_17316# a_66652_17272# 0.28563f
C16869 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN a_59620_23208# 0.00253f
C16870 _300_.A2 a_38876_19975# 0.00259f
C16871 _304_.B vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN 0.0128f
C16872 a_46628_18504# a_47076_18504# 0.01328f
C16873 a_14708_25156# a_14796_25112# 0.28563f
C16874 _375_.Z _378_.I 0.18361f
C16875 a_18292_25156# a_18740_25156# 0.01328f
C16876 a_60909_30600# ui_in[3] 0.50678f
C16877 a_41028_26344# _432_.ZN 0.00116f
C16878 a_46716_13703# a_46628_13800# 0.28563f
C16879 _474_.CLK a_52436_18884# 0.00185f
C16880 _474_.CLK vgaringosc.ro_inv4.inv_array_notouch_\[3\].I 0.037f
C16881 a_29940_20452# a_30388_20452# 0.01328f
C16882 _452_.CLK _441_.A2 0.10419f
C16883 a_54692_20452# a_54332_20408# 0.0869f
C16884 _229_.I a_60276_29032# 0.00199f
C16885 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I 0.00447f
C16886 a_33500_16839# a_33412_16936# 0.28563f
C16887 a_22996_31048# a_23108_29860# 0.02666f
C16888 a_61052_11000# a_60964_9476# 0.00151f
C16889 a_29380_1636# VPWR 0.20348f
C16890 _424_.B1 a_49988_21236# 0.44954f
C16891 a_64188_12568# a_64636_12568# 0.01288f
C16892 _419_.A4 a_47047_21640# 0.00185f
C16893 a_1380_1636# a_1828_1636# 0.01328f
C16894 a_59955_30600# ui_in[1] 0.00105f
C16895 _274_.A2 a_57220_29861# 0.00128f
C16896 _402_.A1 a_46198_27060# 0.0694f
C16897 a_64860_26247# a_65668_26344# 0.00965f
C16898 _398_.C a_46356_24072# 0.01094f
C16899 a_54580_12232# a_54668_10567# 0.00151f
C16900 a_45508_1636# a_45148_1592# 0.08707f
C16901 a_62732_26680# vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN 0.00473f
C16902 a_54420_21976# a_54768_22137# 0.00277f
C16903 _411_.A2 a_48988_27508# 0.00775f
C16904 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN a_60084_25640# 0.00492f
C16905 a_51540_23588# VPWR 0.00407f
C16906 a_48084_18884# a_48060_18407# 0.00172f
C16907 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_56816_26724# 0.00108f
C16908 a_56404_27208# a_57168_26724# 0.00399f
C16909 a_41788_1159# a_42236_1159# 0.0131f
C16910 _441_.A2 a_40316_23233# 0.01049f
C16911 a_932_27912# a_932_26724# 0.05841f
C16912 a_54332_15704# a_54468_15368# 0.00168f
C16913 _402_.A1 clkbuf_1_0__f_clk.I 0.16887f
C16914 _324_.C _325_.ZN 0.00101f
C16915 a_54892_24679# a_54804_24776# 0.28563f
C16916 a_16140_20408# VPWR 0.31143f
C16917 _349_.A4 _371_.A2 0.13893f
C16918 a_66452_16936# a_66900_16936# 0.01328f
C16919 a_54916_12612# VPWR 0.20595f
C16920 _395_.A1 _397_.A4 0.0926f
C16921 a_45956_15368# a_46404_15368# 0.01328f
C16922 a_9532_29383# a_9444_29480# 0.28563f
C16923 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN 0.0017f
C16924 input9.Z a_56348_30951# 0.01327f
C16925 _444_.D a_37472_24419# 0.01513f
C16926 a_47524_10664# VPWR 0.20348f
C16927 a_47836_15271# a_47748_15368# 0.28563f
C16928 _355_.B a_28012_24679# 0.00268f
C16929 a_55700_23588# VPWR 0.20348f
C16930 a_36548_26724# a_36636_26680# 0.28563f
C16931 _251_.A1 ui_in[0] 0.0492f
C16932 a_36172_24463# a_36660_23588# 0.01025f
C16933 _323_.A3 a_35504_18955# 0.00839f
C16934 a_63068_15271# VPWR 0.29679f
C16935 a_49180_15271# a_49852_15271# 0.00544f
C16936 a_19035_28409# a_17472_28363# 0.41622f
C16937 a_16948_22020# a_17036_21976# 0.28563f
C16938 a_20532_22020# a_20980_22020# 0.01328f
C16939 _419_.Z a_51620_19911# 0.00128f
C16940 _474_.Q _384_.A1 0.20123f
C16941 a_61948_2727# a_61860_2824# 0.28563f
C16942 a_25884_27815# VPWR 0.34652f
C16943 a_66652_15704# VPWR 0.32971f
C16944 a_30812_16839# a_31260_16839# 0.0131f
C16945 a_40780_21543# a_40692_21640# 0.28563f
C16946 a_42778_21812# a_42982_21730# 0.4995f
C16947 a_46044_30951# a_45956_31048# 0.28563f
C16948 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN VPWR 0.75343f
C16949 a_27364_23208# a_27452_21543# 0.00151f
C16950 a_65668_7908# VPWR 0.21209f
C16951 a_17508_1256# VPWR 0.20402f
C16952 a_27116_23544# a_27564_23544# 0.01255f
C16953 a_42820_1256# a_43268_1256# 0.01328f
C16954 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN 0.00673f
C16955 a_67460_4772# VPWR 0.20348f
C16956 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I 0.00859f
C16957 a_56572_23111# a_57020_23111# 0.012f
C16958 a_57580_13703# a_57940_13800# 0.08707f
C16959 a_54556_14136# a_54468_12612# 0.00151f
C16960 a_3620_13800# a_4068_13800# 0.01328f
C16961 a_7964_29383# VPWR 0.35803f
C16962 a_21852_2727# a_22300_2727# 0.0131f
C16963 a_63316_20452# a_63404_20408# 0.28563f
C16964 _330_.A1 a_38506_26724# 0.01351f
C16965 _417_.A2 a_51892_23340# 0.00984f
C16966 _399_.A2 a_48321_23208# 0.10952f
C16967 a_44364_16839# a_44724_16936# 0.08707f
C16968 a_49652_10664# a_49540_9476# 0.02666f
C16969 a_59820_10567# a_59844_9476# 0.0016f
C16970 a_3260_1159# a_3172_1256# 0.28563f
C16971 a_32964_16936# VPWR 0.20348f
C16972 a_35516_1592# VPWR 0.32932f
C16973 a_36612_20072# VPWR 0.01386f
C16974 a_21964_23544# a_21852_23111# 0.02634f
C16975 _424_.A2 a_51877_21236# 0.00248f
C16976 a_61500_12568# a_61612_12135# 0.02634f
C16977 a_8100_1636# a_8772_1636# 0.00347f
C16978 a_6756_29860# a_7204_29860# 0.01328f
C16979 a_3172_29860# a_3260_29816# 0.28563f
C16980 _324_.C _400_.ZN 0.31588f
C16981 _424_.A2 a_46794_25156# 0.00492f
C16982 a_40580_20452# _327_.Z 0.00109f
C16983 a_4156_17272# a_4604_17272# 0.01222f
C16984 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN a_65072_29860# 0.04688f
C16985 a_44252_30951# VPWR 0.31143f
C16986 a_49316_11044# a_49292_10567# 0.00172f
C16987 _362_.B _371_.A1 0.18907f
C16988 a_45372_11000# a_45372_10567# 0.05841f
C16989 _452_.CLK a_46180_18504# 0.00111f
C16990 a_58588_11000# a_59036_11000# 0.01288f
C16991 a_48420_1636# a_48508_1592# 0.28563f
C16992 a_52004_1636# a_52452_1636# 0.01328f
C16993 a_60156_27815# a_60604_27815# 0.01255f
C16994 _304_.B a_53460_24776# 0.00162f
C16995 _416_.A1 a_46848_20893# 0.02046f
C16996 _448_.Q a_38764_20408# 0.0052f
C16997 a_48060_18407# a_47972_18504# 0.28563f
C16998 a_17396_27912# a_17168_27165# 0.00186f
C16999 _470_.Q _419_.A4 0.00287f
C17000 a_20308_27912# a_20308_26724# 0.05841f
C17001 a_33776_29123# _335_.ZN 0.01034f
C17002 a_15604_25156# VPWR 0.20348f
C17003 _441_.ZN _439_.ZN 0.04362f
C17004 a_66564_18884# a_66204_18840# 0.0869f
C17005 a_67884_18407# VPWR 0.33379f
C17006 a_932_27912# a_1380_27912# 0.01328f
C17007 a_15244_27815# a_15604_27912# 0.08717f
C17008 a_27116_20408# VPWR 0.36297f
C17009 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I a_58836_17316# 0.00696f
C17010 a_61500_12568# VPWR 0.31389f
C17011 a_22660_2824# a_23108_2824# 0.01328f
C17012 _447_.Q _319_.A2 0.66534f
C17013 _337_.ZN a_30520_27508# 0.00188f
C17014 a_18096_27165# uio_out[7] 0.81831f
C17015 a_41028_26344# _260_.A1 0.00141f
C17016 _284_.ZN _452_.CLK 0.00711f
C17017 _317_.A2 a_37744_20452# 0.00869f
C17018 a_67548_8999# a_67460_9096# 0.28563f
C17019 _316_.ZN a_35268_21640# 0.00188f
C17020 _371_.A1 a_32628_26725# 0.00497f
C17021 a_16948_21640# a_16948_20452# 0.05841f
C17022 a_19320_28409# VPWR 0.00302f
C17023 a_45012_29816# a_45408_30345# 0.00232f
C17024 a_63540_16936# VPWR 0.20703f
C17025 _218_.ZN a_49988_21236# 0.26075f
C17026 a_43044_15368# VPWR 0.2117f
C17027 a_17472_28363# uio_out[7] 0.07132f
C17028 _294_.A2 a_35740_30951# 0.00202f
C17029 a_46492_15271# VPWR 0.29679f
C17030 a_4156_14136# a_4604_14136# 0.01222f
C17031 a_2812_16839# VPWR 0.30213f
C17032 a_45620_16936# a_45732_15748# 0.02666f
C17033 a_41812_16936# a_41788_15704# 0.0016f
C17034 a_39908_1256# VPWR 0.20348f
C17035 a_25012_31048# _342_.ZN 0.00225f
C17036 a_67100_3160# a_67100_2727# 0.05841f
C17037 a_932_13800# a_932_12612# 0.05841f
C17038 _358_.A2 VPWR 0.24102f
C17039 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN VPWR 0.83474f
C17040 _397_.A2 _421_.A1 0.40827f
C17041 _459_.Q _287_.A1 0.00109f
C17042 _474_.CLK a_55788_23544# 0.03242f
C17043 a_1468_17272# VPWR 0.29679f
C17044 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN 0.16849f
C17045 a_49316_1636# VPWR 0.20761f
C17046 _246_.B2 a_61297_30300# 0.18809f
C17047 vgaringosc.workerclkbuff_notouch_.I a_43916_29816# 0.02892f
C17048 a_54804_16936# VPWR 0.20782f
C17049 a_14236_1159# a_14596_1256# 0.08717f
C17050 a_4940_12135# a_5300_12232# 0.08674f
C17051 a_11460_1636# a_11548_1592# 0.28563f
C17052 a_15044_1636# a_15492_1636# 0.01328f
C17053 a_49852_12568# a_49764_11044# 0.00151f
C17054 a_7428_29480# a_7876_29480# 0.01328f
C17055 a_58476_12135# a_58924_12135# 0.01288f
C17056 a_29716_23588# a_29692_23111# 0.00172f
C17057 _386_.ZN a_47376_27912# 0.0063f
C17058 _416_.A1 a_43736_25896# 0.01855f
C17059 a_36548_17316# a_36188_17272# 0.08707f
C17060 a_44612_31048# a_45060_31048# 0.01328f
C17061 a_65892_11044# a_65980_11000# 0.28563f
C17062 a_31620_1636# a_31484_1159# 0.00168f
C17063 a_27676_1592# a_27676_1159# 0.05841f
C17064 _424_.A1 a_51620_19911# 0.00799f
C17065 _459_.CLK a_19860_26724# 0.01886f
C17066 _459_.Q a_31932_26247# 0.00271f
C17067 a_19972_2824# VPWR 0.22918f
C17068 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62196_26724# 0.01551f
C17069 a_53460_24776# VPWR 0.16303f
C17070 _395_.A2 _384_.A1 0.00682f
C17071 a_3260_24679# a_3172_24776# 0.28563f
C17072 _397_.A1 _397_.A4 0.06726f
C17073 a_20956_24679# a_21404_24679# 0.01288f
C17074 a_3708_19975# a_4156_19975# 0.0131f
C17075 a_62284_26680# _245_.I1 0.0061f
C17076 a_64188_1159# a_64636_1159# 0.0131f
C17077 _434_.ZN a_39332_23588# 0.02026f
C17078 a_48868_2824# a_48868_1636# 0.05841f
C17079 a_21740_29383# a_22100_29480# 0.0869f
C17080 a_1380_5960# a_1828_5960# 0.01328f
C17081 a_1468_14136# VPWR 0.29679f
C17082 a_2276_4392# a_2724_4392# 0.01328f
C17083 _355_.ZN VPWR 0.34754f
C17084 _352_.A2 a_26756_24801# 0.01674f
C17085 _304_.A1 a_42778_21812# 0.01638f
C17086 _229_.I a_62564_29032# 0.49164f
C17087 _459_.CLK _378_.ZN 0.01417f
C17088 _448_.Q a_37360_19325# 0.20874f
C17089 a_37444_15748# a_37532_15704# 0.28563f
C17090 a_51791_30644# _274_.ZN 0.00465f
C17091 a_33500_15704# a_33948_15704# 0.01288f
C17092 a_4740_29480# VPWR 0.22961f
C17093 a_55564_12135# VPWR 0.31547f
C17094 _378_.I a_19860_27912# 0.00158f
C17095 _251_.A1 _274_.A1 0.0016f
C17096 _358_.A3 a_35740_26247# 0.01497f
C17097 _287_.A1 _461_.D 0.01232f
C17098 _290_.ZN _460_.Q 0.05429f
C17099 a_27228_26247# _457_.D 0.00134f
C17100 a_57500_30344# a_57220_29861# 0.00126f
C17101 _352_.ZN a_26746_26344# 0.00927f
C17102 a_17932_24679# VPWR 0.32173f
C17103 a_23780_26344# a_24228_26344# 0.01328f
C17104 a_59332_29816# a_59948_30352# 0.00478f
C17105 _281_.ZN a_47297_25596# 0.01647f
C17106 a_44948_28292# a_45396_28292# 0.01328f
C17107 a_41642_25156# VPWR 0.0149f
C17108 a_30812_15704# VPWR 0.30073f
C17109 a_33028_27912# VPWR 0.01455f
C17110 _311_.A2 a_36560_22512# 0.0032f
C17111 a_48956_18407# a_49404_18407# 0.012f
C17112 a_3620_9476# a_3708_9432# 0.28563f
C17113 a_26668_21976# a_27116_21976# 0.01288f
C17114 hold2.Z _284_.B 0.10897f
C17115 _381_.Z a_47924_28292# 0.00593f
C17116 _303_.ZN a_43380_20452# 0.02059f
C17117 a_11091_30644# uio_oe[3] 0.00151f
C17118 _281_.A1 _427_.B2 0.57531f
C17119 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN 0.01877f
C17120 a_46268_18407# VPWR 0.32882f
C17121 a_51108_14180# a_50748_14136# 0.08707f
C17122 a_52652_16839# a_53100_16839# 0.0131f
C17123 _452_.CLK a_41048_17341# 0.02743f
C17124 _229_.I a_63092_26724# 0.002f
C17125 a_48756_16936# a_48732_15704# 0.0016f
C17126 a_52564_16936# a_52676_15748# 0.02666f
C17127 a_49740_16839# VPWR 0.35134f
C17128 a_64996_1256# a_65668_1256# 0.00347f
C17129 a_62308_1256# VPWR 0.20348f
C17130 _384_.A1 a_50196_22805# 0.01549f
C17131 a_65332_13800# a_65780_13800# 0.01328f
C17132 a_44252_2727# a_44700_2727# 0.0131f
C17133 a_49204_13800# a_49316_12612# 0.02666f
C17134 a_55588_28292# a_55228_28248# 0.08674f
C17135 _424_.B1 clkbuf_1_0__f_clk.I 0.01946f
C17136 a_44752_18147# a_45260_17272# 0.00136f
C17137 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I a_61164_23111# 0.00409f
C17138 _475_.Q a_52240_22504# 0.00731f
C17139 _421_.B a_47524_22021# 0.09337f
C17140 _304_.B clkload0.Z 0.00463f
C17141 a_44276_17316# VPWR 0.11759f
C17142 a_25660_1159# a_25572_1256# 0.28563f
C17143 a_61724_1592# a_61860_1256# 0.00168f
C17144 a_62980_1636# VPWR 0.2147f
C17145 _397_.A1 a_51956_26183# 0.03028f
C17146 a_55564_12135# a_55476_12232# 0.28563f
C17147 _355_.ZN a_28903_24776# 0.07669f
C17148 a_1916_21543# VPWR 0.297f
C17149 a_12892_29816# a_13340_29816# 0.01288f
C17150 _452_.Q a_38876_19975# 0.00281f
C17151 a_3172_26344# a_3172_25156# 0.05841f
C17152 _336_.A2 a_29804_23544# 0.00179f
C17153 _336_.A1 a_29716_23588# 0.00182f
C17154 a_45820_15704# a_45732_14180# 0.0027f
C17155 a_44276_17316# a_44364_17272# 0.28563f
C17156 a_41536_17636# a_41432_17801# 0.10745f
C17157 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN a_59708_23111# 0.00284f
C17158 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I a_55252_26724# 0.00916f
C17159 a_55588_27912# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.00656f
C17160 a_58836_18884# vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I 0.00197f
C17161 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN a_58924_18840# 0.02703f
C17162 a_45372_10567# a_45820_10567# 0.0131f
C17163 a_42148_2824# VPWR 0.22175f
C17164 _416_.A1 _417_.A2 0.1461f
C17165 a_38564_1636# a_38428_1159# 0.00168f
C17166 a_34620_1592# a_34620_1159# 0.05841f
C17167 a_58140_1592# a_58588_1592# 0.01288f
C17168 a_62084_1636# a_62172_1592# 0.28563f
C17169 a_31484_23111# a_31932_23111# 0.01288f
C17170 a_19612_23111# a_19972_23208# 0.08707f
C17171 _330_.A1 _319_.A3 0.43385f
C17172 a_23196_24679# a_23556_24776# 0.08707f
C17173 a_45372_9432# VPWR 0.31538f
C17174 a_60604_27815# a_60516_27912# 0.28563f
C17175 a_4940_21543# a_5388_21543# 0.01222f
C17176 a_54916_14180# VPWR 0.20348f
C17177 a_36076_18407# a_35988_18504# 0.28563f
C17178 _267_.A1 a_53660_27815# 0.00126f
C17179 _397_.A2 _409_.ZN 0.07236f
C17180 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN _249_.A2 0.16497f
C17181 _439_.ZN _437_.ZN 0.32126f
C17182 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I 0.87086f
C17183 _362_.B a_34700_28776# 0.0013f
C17184 a_49652_12232# VPWR 0.21158f
C17185 a_40804_15748# a_40444_15704# 0.08707f
C17186 a_45060_2824# a_45508_2824# 0.01328f
C17187 _421_.A1 a_47860_21640# 0.14499f
C17188 _316_.A3 a_36548_21640# 0.00641f
C17189 a_59955_30600# _324_.C 0.009f
C17190 _402_.A1 a_43003_28409# 0.02931f
C17191 _474_.CLK _412_.B2 0.11798f
C17192 a_3260_20408# a_3260_19975# 0.05841f
C17193 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_54804_26724# 0.02723f
C17194 a_22660_24776# VPWR 0.20622f
C17195 _294_.A2 a_31396_26724# 0.01138f
C17196 a_42996_18840# a_43784_19369# 0.02112f
C17197 a_5724_2727# a_5636_2824# 0.28563f
C17198 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_63764_23588# 0.00313f
C17199 a_44476_15704# VPWR 0.29679f
C17200 a_32156_19975# a_32516_20072# 0.08717f
C17201 a_21652_29480# a_21628_28248# 0.0016f
C17202 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN 0.00254f
C17203 a_48060_9432# a_48508_9432# 0.0131f
C17204 _474_.Q clk 0.06889f
C17205 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I a_57156_27912# 0.0023f
C17206 a_66092_19975# VPWR 0.3734f
C17207 _452_.CLK a_39772_26247# 0.00629f
C17208 a_54468_14180# a_54556_14136# 0.28563f
C17209 a_15580_29383# a_15604_28292# 0.0016f
C17210 a_20620_25112# a_20532_23588# 0.00151f
C17211 _265_.ZN _470_.D 0.00568f
C17212 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.30902f
C17213 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_61940_29076# 0.01136f
C17214 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN a_63721_28776# 0.00745f
C17215 _474_.CLK a_55252_24776# 0.01743f
C17216 clkload0.Z VPWR 0.34482f
C17217 a_37532_26247# VPWR 0.29679f
C17218 a_52316_17272# VPWR 0.31547f
C17219 _336_.A2 _457_.D 0.02958f
C17220 _327_.A2 a_45820_18407# 0.009f
C17221 a_5276_1159# VPWR 0.3289f
C17222 a_36636_1159# a_36996_1256# 0.08717f
C17223 a_50188_12135# a_50212_11044# 0.0016f
C17224 a_21180_1592# a_21628_1592# 0.01288f
C17225 a_66316_12135# a_66676_12232# 0.08717f
C17226 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN 0.00103f
C17227 a_52340_12232# a_52788_12232# 0.01328f
C17228 _451_.Q a_40220_19975# 0.04206f
C17229 a_32828_21543# VPWR 0.3215f
C17230 _397_.A2 a_48988_27508# 0.00244f
C17231 _441_.ZN _303_.ZN 0.47943f
C17232 a_20496_26344# a_21876_25156# 0.00999f
C17233 a_21424_25987# a_21428_25156# 0.00254f
C17234 a_21052_26031# a_20980_25156# 0.00175f
C17235 a_48644_17316# a_48284_17272# 0.08707f
C17236 _448_.Q a_44028_22020# 0.0011f
C17237 a_2812_10567# a_2724_10664# 0.28563f
C17238 a_66788_1636# a_66876_1592# 0.28563f
C17239 a_64548_2824# VPWR 0.20655f
C17240 a_30588_23111# a_30500_23208# 0.28563f
C17241 _388_.B a_43828_29860# 0.01534f
C17242 _452_.CLK a_32592_25227# 0.00499f
C17243 a_25348_24776# a_25796_24776# 0.01328f
C17244 a_3260_21543# a_3620_21640# 0.08717f
C17245 _327_.Z _331_.ZN 0.60298f
C17246 a_59844_9476# VPWR 0.21241f
C17247 a_1380_23588# VPWR 0.20348f
C17248 a_1380_6340# VPWR 0.20348f
C17249 a_3172_3204# VPWR 0.20993f
C17250 _238_.ZN a_59348_29076# 0.00167f
C17251 a_63292_14136# VPWR 0.31389f
C17252 _459_.CLK a_30724_26020# 0.00503f
C17253 _411_.A2 a_51883_27508# 0.00987f
C17254 a_47300_15748# a_47748_15748# 0.01328f
C17255 a_3620_11044# VPWR 0.22347f
C17256 a_10564_29860# a_10428_29383# 0.00168f
C17257 _284_.ZN a_41440_28363# 0.04434f
C17258 _229_.I _250_.B 0.18497f
C17259 a_63516_19975# a_63428_20072# 0.28563f
C17260 _427_.A2 _384_.A1 0.25703f
C17261 _386_.A4 a_47376_27912# 0.00451f
C17262 a_30160_30301# a_29788_30345# 0.10745f
C17263 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN 0.00766f
C17264 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I a_57156_27912# 0.02057f
C17265 a_22100_29480# a_22548_29480# 0.01328f
C17266 _294_.ZN a_30388_28776# 0.02975f
C17267 a_4604_18840# VPWR 0.33016f
C17268 a_57168_26724# VPWR 0.01056f
C17269 _313_.ZN a_34586_23208# 0.00488f
C17270 a_16700_2727# a_17060_2824# 0.08717f
C17271 a_25652_31048# _340_.ZN 0.00101f
C17272 a_44744_26355# a_46156_26031# 0.00393f
C17273 _454_.Q _346_.A2 0.19501f
C17274 a_53796_9476# a_53884_9432# 0.28563f
C17275 a_51420_17272# a_51332_15748# 0.00151f
C17276 _470_.Q _381_.A2 0.00707f
C17277 a_2364_20408# a_2812_20408# 0.0131f
C17278 a_4964_20452# a_4604_20408# 0.08674f
C17279 _251_.ZN a_59652_25640# 0.02319f
C17280 _424_.A1 a_54040_22366# 0.00415f
C17281 _452_.CLK a_32292_21640# 0.002f
C17282 _330_.ZN a_38336_18147# 0.01413f
C17283 a_37408_18504# a_37964_18191# 0.8399f
C17284 a_66652_2727# a_67100_2727# 0.01255f
C17285 a_46716_12568# a_47164_12568# 0.01288f
C17286 a_50660_12612# a_50748_12568# 0.28563f
C17287 _438_.ZN a_40332_21543# 0.00635f
C17288 _452_.Q a_39684_20452# 0.01062f
C17289 a_27676_1159# VPWR 0.30414f
C17290 a_48060_1159# a_47972_1256# 0.28563f
C17291 a_4852_7528# a_4940_5863# 0.00151f
C17292 a_57132_12135# a_57156_11044# 0.0016f
C17293 _294_.A2 VPWR 2.79508f
C17294 a_66876_12568# a_66788_11044# 0.00151f
C17295 a_47076_12232# a_47076_11044# 0.05841f
C17296 _381_.A2 a_50464_24908# 0.00727f
C17297 a_28484_1636# a_28124_1592# 0.08707f
C17298 a_40220_26247# a_40668_26247# 0.01255f
C17299 a_36636_26247# a_36996_26344# 0.08674f
C17300 _422_.ZN a_52512_19715# 0.00127f
C17301 a_30052_21640# VPWR 0.20641f
C17302 _319_.A3 a_35723_20569# 0.0592f
C17303 a_53324_10567# a_53684_10664# 0.08707f
C17304 a_67212_10567# a_67660_10567# 0.0131f
C17305 a_7964_1159# a_8636_1159# 0.00544f
C17306 _285_.Z _402_.A1 0.24247f
C17307 a_47552_19715# VPWR 0.51815f
C17308 a_2276_22020# VPWR 0.20634f
C17309 _395_.A2 clk 0.02533f
C17310 a_31803_24831# a_32048_24463# 0.00232f
C17311 a_29156_23208# a_29604_23208# 0.01328f
C17312 _416_.A1 _267_.A2 0.00605f
C17313 a_19724_23544# VPWR 0.32344f
C17314 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN 0.62866f
C17315 a_64412_5863# VPWR 0.3038f
C17316 a_3708_8999# VPWR 0.33374f
C17317 a_37892_2824# a_37980_1159# 0.0027f
C17318 a_23644_21543# a_23556_21640# 0.28563f
C17319 a_1828_21640# a_2276_21640# 0.01328f
C17320 _409_.ZN _330_.A1 0.40052f
C17321 a_7516_2727# VPWR 0.31143f
C17322 a_57580_13703# VPWR 0.32122f
C17323 _459_.CLK a_26970_29480# 0.00269f
C17324 a_60516_27912# a_60964_27912# 0.01328f
C17325 a_46984_23588# clk 0.00393f
C17326 a_52540_11000# VPWR 0.34431f
C17327 a_16700_29816# a_16700_29383# 0.05841f
C17328 a_2812_21976# a_2812_21543# 0.05841f
C17329 a_46716_2727# a_46852_1636# 0.00154f
C17330 a_67460_2824# a_67908_2824# 0.01328f
C17331 _325_.B a_43444_19668# 0.00189f
C17332 a_3708_26680# VPWR 0.33374f
C17333 vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN clk 0.00105f
C17334 a_33636_23208# a_33708_22505# 0.00175f
C17335 _398_.C _412_.B2 0.02967f
C17336 a_61388_15704# a_62172_15704# 0.00443f
C17337 a_64772_15748# a_65220_15748# 0.01328f
C17338 a_33164_20408# a_33052_19975# 0.02634f
C17339 a_9635_30644# uio_oe[5] 0.04236f
C17340 _371_.A3 a_30724_26020# 0.00182f
C17341 a_21424_25987# VPWR 0.18741f
C17342 a_27588_26724# a_27676_26680# 0.28563f
C17343 a_28124_2727# a_28036_2824# 0.28563f
C17344 _435_.A3 _325_.A1 0.00116f
C17345 a_59260_21976# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I 0.08702f
C17346 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I VPWR 1.06346f
C17347 _439_.ZN a_41488_24072# 0.02235f
C17348 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN a_61972_20452# 0.00205f
C17349 a_14796_28248# VPWR 0.30073f
C17350 a_1380_7908# a_1020_7864# 0.08717f
C17351 a_3172_7908# a_3620_7908# 0.01328f
C17352 a_59036_9432# a_59484_9432# 0.0131f
C17353 a_4068_23588# a_4516_23588# 0.01328f
C17354 a_8996_1256# a_9444_1256# 0.01328f
C17355 a_2276_23588# a_1916_23544# 0.08717f
C17356 a_2276_6340# a_1916_6296# 0.08717f
C17357 a_12916_31048# a_13364_31048# 0.01328f
C17358 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN _245_.I1 0.7364f
C17359 _474_.Q _416_.A3 0.0502f
C17360 _279_.Z _475_.Q 0.12808f
C17361 a_4068_6340# a_4516_6340# 0.01328f
C17362 a_65980_14136# a_66428_14136# 0.01288f
C17363 a_4068_3204# a_3708_3160# 0.08717f
C17364 a_1468_3160# a_1916_3160# 0.0131f
C17365 a_3172_4772# a_2812_4728# 0.08717f
C17366 a_66092_16839# a_66116_15748# 0.0016f
C17367 a_4740_31048# a_4828_29383# 0.0027f
C17368 a_60909_30600# _256_.A2 0.00215f
C17369 a_57492_23588# a_57580_23544# 0.28563f
C17370 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN a_57132_23544# 0.00142f
C17371 a_1468_1592# VPWR 0.29679f
C17372 a_39300_29480# uo_out[1] 0.00421f
C17373 a_54020_12612# a_53660_12568# 0.08707f
C17374 _459_.CLK a_19636_25156# 0.00252f
C17375 a_56372_13800# a_56460_12135# 0.00151f
C17376 _452_.CLK _331_.ZN 0.01642f
C17377 _416_.A2 a_47724_18840# 0.00642f
C17378 a_34715_22137# _316_.A3 0.03712f
C17379 a_59036_1159# a_59396_1256# 0.08717f
C17380 _436_.B uo_out[7] 0.00292f
C17381 a_54132_12232# a_54020_11044# 0.02666f
C17382 a_49852_1159# VPWR 0.33324f
C17383 a_4516_11044# a_4156_11000# 0.08674f
C17384 a_1916_11000# a_2364_11000# 0.0131f
C17385 a_67460_18884# VPWR 0.20692f
C17386 a_32592_25227# a_34448_25597# 0.02307f
C17387 a_33520_25597# a_33148_25641# 0.10745f
C17388 a_66988_16839# a_67436_16839# 0.01255f
C17389 a_34980_1636# a_35428_1636# 0.01328f
C17390 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN a_64860_26247# 0.00108f
C17391 _359_.B _285_.Z 0.06385f
C17392 a_45416_29885# _397_.A1 0.004f
C17393 _311_.A2 a_36544_24419# 0.00511f
C17394 a_64300_10567# a_64212_10664# 0.28563f
C17395 _346_.A2 a_23284_26724# 0.02028f
C17396 _272_.A2 _258_.ZN 0.00232f
C17397 _359_.B a_44476_27815# 0.00122f
C17398 _459_.CLK _337_.ZN 0.05319f
C17399 a_60909_30600# a_61029_31220# 0.00165f
C17400 a_20620_21976# VPWR 0.31589f
C17401 a_32268_23544# VPWR 0.32796f
C17402 a_30724_18884# a_30812_18840# 0.28563f
C17403 a_29916_2727# VPWR 0.31143f
C17404 a_51444_13800# VPWR 0.20595f
C17405 a_32516_18884# a_32964_18884# 0.01328f
C17406 _459_.Q a_34308_26344# 0.00732f
C17407 a_2364_26247# a_2812_26247# 0.0131f
C17408 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN 0.00449f
C17409 _267_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN 0.04559f
C17410 _399_.A2 _399_.A1 0.82446f
C17411 a_6844_29816# VPWR 0.3289f
C17412 a_66340_11044# VPWR 0.2154f
C17413 _251_.A1 _250_.ZN 0.41458f
C17414 _324_.B a_44038_21236# 0.02712f
C17415 _416_.A1 a_44736_26031# 0.00128f
C17416 a_53660_2727# a_53796_1636# 0.00154f
C17417 a_17484_23111# VPWR 0.29719f
C17418 _304_.A1 _301_.A1 0.70589f
C17419 _447_.Q _441_.A2 0.95181f
C17420 _247_.ZN a_59172_27912# 0.12599f
C17421 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I a_67908_22020# 0.01186f
C17422 a_17844_27912# VPWR 0.21272f
C17423 _437_.A1 a_38752_26344# 0.01003f
C17424 _399_.ZN a_48321_23208# 0.53153f
C17425 _260_.A1 a_41776_20072# 0.00106f
C17426 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I 0.00213f
C17427 _370_.ZN a_29664_29977# 0.00242f
C17428 a_25124_28776# _371_.A2 1.66226f
C17429 a_39100_2727# a_39460_2824# 0.08717f
C17430 a_56036_28292# VPWR 0.20836f
C17431 _355_.C a_27140_26724# 0.00153f
C17432 a_54244_18884# a_54692_18884# 0.01328f
C17433 a_61388_16839# a_61300_16936# 0.28563f
C17434 a_66564_7908# a_66204_7864# 0.08717f
C17435 a_16052_23588# a_15692_23544# 0.08707f
C17436 a_3260_7864# a_3260_7431# 0.05841f
C17437 a_64772_9476# a_64860_9432# 0.28563f
C17438 a_4156_6296# a_4156_5863# 0.05841f
C17439 a_67460_6340# a_67100_6296# 0.08717f
C17440 a_2724_25156# a_3172_25156# 0.01328f
C17441 a_63292_14136# a_63404_13703# 0.02634f
C17442 a_54332_18840# VPWR 0.32052f
C17443 a_62148_29505# _250_.C 0.03406f
C17444 a_64324_20072# a_64324_18884# 0.05841f
C17445 a_22412_20408# a_22860_20408# 0.0131f
C17446 a_24564_20452# a_24204_20408# 0.08717f
C17447 _390_.ZN _411_.A2 0.05389f
C17448 a_14004_31048# a_14372_31048# 0.02601f
C17449 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN VPWR 0.77069f
C17450 a_15132_1592# VPWR 0.29679f
C17451 a_60380_12568# a_60964_12612# 0.01675f
C17452 a_23920_27555# a_24900_27912# 0.00211f
C17453 a_23627_27967# _351_.A2 0.00125f
C17454 a_51108_12612# a_51084_12135# 0.00172f
C17455 a_47164_12568# a_47164_12135# 0.05841f
C17456 a_49764_31048# vgaringosc.workerclkbuff_notouch_.I 0.00648f
C17457 _386_.A4 a_46580_28292# 0.00109f
C17458 _359_.B a_32820_29535# 0.00127f
C17459 a_42168_22504# a_42784_22504# 0.00951f
C17460 _275_.ZN _324_.C 0.05365f
C17461 a_61076_12232# a_60964_11044# 0.02666f
C17462 a_66116_9096# VPWR 0.23643f
C17463 _351_.ZN VPWR 0.53799f
C17464 a_932_4772# VPWR 0.22176f
C17465 a_48868_11044# a_48508_11000# 0.08707f
C17466 a_1828_18504# VPWR 0.20348f
C17467 a_65108_23588# a_64748_23544# 0.08674f
C17468 a_26160_27165# a_25643_25273# 0.00122f
C17469 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I 0.00618f
C17470 a_61076_10664# a_61524_10664# 0.01328f
C17471 a_67741_30600# vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.03313f
C17472 a_30364_1159# a_30812_1159# 0.0131f
C17473 a_66788_1636# a_66652_1159# 0.00168f
C17474 a_23108_24776# a_23196_23111# 0.00151f
C17475 a_27588_2824# a_27588_1636# 0.05841f
C17476 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN rst_n 0.00542f
C17477 _324_.B _325_.A2 0.03098f
C17478 _395_.A3 a_50732_23233# 0.00836f
C17479 a_32268_21976# VPWR 0.32364f
C17480 a_40780_27815# a_39536_26795# 0.00102f
C17481 a_39268_18840# _330_.A2 0.02985f
C17482 a_32740_21640# a_33188_21640# 0.01328f
C17483 a_1020_12568# VPWR 0.30073f
C17484 _421_.A1 a_47483_20569# 0.00979f
C17485 a_52316_2727# VPWR 0.31143f
C17486 a_17484_26247# a_17396_26344# 0.28563f
C17487 _452_.CLK a_37888_27555# 0.00613f
C17488 a_62172_18407# a_62532_18504# 0.08717f
C17489 a_34532_15368# a_34980_15368# 0.01328f
C17490 a_20672_30301# VPWR 1.03095f
C17491 _337_.A3 VPWR 2.43876f
C17492 a_36412_15271# a_36324_15368# 0.28563f
C17493 _337_.ZN _371_.A3 0.34895f
C17494 a_53324_10567# VPWR 0.31547f
C17495 a_56036_27912# VPWR 0.20734f
C17496 a_25772_21976# a_25884_21543# 0.02634f
C17497 a_29716_22020# a_29692_21543# 0.00172f
C17498 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN 0.03075f
C17499 a_15156_23208# VPWR 0.20348f
C17500 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN 0.63827f
C17501 a_37756_15271# a_38428_15271# 0.00544f
C17502 _439_.ZN a_40880_23588# 0.0015f
C17503 a_2276_28292# a_2364_28248# 0.28563f
C17504 _274_.A1 a_55676_28248# 0.00156f
C17505 _268_.A2 _272_.A2 0.24741f
C17506 a_3172_22020# a_2812_21976# 0.08717f
C17507 a_50120_26476# VPWR 0.34986f
C17508 a_50524_2727# a_50436_2824# 0.28563f
C17509 a_62172_17272# a_62620_17272# 0.0131f
C17510 a_66564_17316# a_66204_17272# 0.0869f
C17511 _281_.ZN a_51618_22504# 0.00119f
C17512 a_4852_16936# a_4964_15748# 0.02666f
C17513 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN a_59172_23208# 0.00601f
C17514 a_65308_8999# a_65756_8999# 0.0131f
C17515 a_22548_23588# a_22996_23588# 0.01328f
C17516 a_31396_1256# a_31844_1256# 0.01328f
C17517 a_60285_30600# ui_in[3] 0.09407f
C17518 a_67100_5863# a_67548_5863# 0.0131f
C17519 a_66204_7431# a_66652_7431# 0.0131f
C17520 a_1020_18840# a_1020_18407# 0.05841f
C17521 a_10428_2727# a_10876_2727# 0.0131f
C17522 _474_.CLK a_54000_30344# 0.00206f
C17523 a_50748_14136# a_50660_12612# 0.00151f
C17524 a_60268_13703# a_60716_13703# 0.01288f
C17525 a_46268_13703# a_46628_13800# 0.08717f
C17526 a_67796_18504# a_67908_17316# 0.02666f
C17527 a_54244_20452# a_54332_20408# 0.28563f
C17528 _402_.A1 _412_.A1 0.10821f
C17529 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN 0.00258f
C17530 a_62308_26344# _245_.I1 0.02934f
C17531 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_65108_23588# 0.00101f
C17532 a_33052_16839# a_33412_16936# 0.08717f
C17533 a_2724_10664# a_2724_9476# 0.05841f
C17534 _355_.C _379_.Z 0.05725f
C17535 a_28932_1636# VPWR 0.20348f
C17536 uio_oe[7] uio_oe[6] 0.05393f
C17537 a_58052_12612# a_58028_12135# 0.00172f
C17538 a_54108_12568# a_54220_12135# 0.02634f
C17539 a_53616_29480# VPWR 0.01626f
C17540 a_14460_30951# a_14908_30951# 0.01222f
C17541 a_67684_12612# a_67772_12568# 0.28563f
C17542 _388_.B _383_.A2 0.28226f
C17543 _337_.ZN uo_out[7] 0.02646f
C17544 a_64772_18504# a_65220_18504# 0.01328f
C17545 _274_.A2 a_56596_29861# 0.13237f
C17546 a_38523_27967# a_38768_27599# 0.00232f
C17547 a_3620_15368# a_3620_14180# 0.05841f
C17548 a_46516_16936# a_46964_16936# 0.01328f
C17549 a_13340_1592# a_13340_1159# 0.05841f
C17550 a_41116_1592# a_41564_1592# 0.01288f
C17551 a_45060_1636# a_45148_1592# 0.28563f
C17552 a_55364_11044# a_55812_11044# 0.01328f
C17553 _284_.ZN _447_.Q 0.00417f
C17554 a_49764_23588# VPWR 0.01045f
C17555 _424_.A1 a_54556_21543# 0.00255f
C17556 _411_.A2 a_48580_27508# 0.00181f
C17557 a_14796_26680# a_15244_26680# 0.01222f
C17558 a_56404_27208# a_56816_26724# 0.00736f
C17559 a_34532_2824# a_34532_1636# 0.05841f
C17560 _441_.A2 a_40004_23233# 0.01491f
C17561 a_54444_24679# a_54804_24776# 0.0869f
C17562 a_15692_20408# VPWR 0.31143f
C17563 a_62503_28293# a_63105_28293# 0.07676f
C17564 a_54468_12612# VPWR 0.20595f
C17565 _268_.A2 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN 0.04825f
C17566 _355_.B a_28756_25940# 0.00233f
C17567 _363_.Z a_34084_28776# 0.00424f
C17568 a_11236_2824# a_11684_2824# 0.01328f
C17569 _359_.B _371_.A1 0.04562f
C17570 a_7628_30951# uio_oe[7] 0.00187f
C17571 a_9084_29383# a_9444_29480# 0.08717f
C17572 _294_.A2 _370_.B 0.08314f
C17573 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _276_.A2 0.01292f
C17574 _444_.D a_37179_24831# 0.01312f
C17575 _304_.A1 a_42252_20936# 0.17207f
C17576 a_47076_10664# VPWR 0.20348f
C17577 a_47388_15271# a_47748_15368# 0.08717f
C17578 a_24428_21976# a_24452_21640# 0.00172f
C17579 a_55252_23588# VPWR 0.20348f
C17580 a_36548_26724# a_36188_26680# 0.0869f
C17581 _260_.A1 a_44491_20936# 0.00943f
C17582 a_35616_24776# a_37108_23588# 0.00103f
C17583 a_62620_15271# VPWR 0.29679f
C17584 _241_.Z a_58052_26724# 0.06889f
C17585 _229_.I _245_.Z 0.00164f
C17586 _373_.A2 _373_.ZN 0.39292f
C17587 _419_.Z a_49448_20072# 0.00172f
C17588 a_61276_2727# a_61860_2824# 0.01675f
C17589 a_66204_15704# VPWR 0.35041f
C17590 a_16948_22020# a_16588_21976# 0.08707f
C17591 a_64996_15368# a_65444_15368# 0.01328f
C17592 a_21044_27508# VPWR 0.80432f
C17593 _424_.A2 hold1.Z 0.0175f
C17594 a_42154_21236# a_42982_21730# 0.00135f
C17595 a_40332_21543# a_40692_21640# 0.08674f
C17596 a_45596_30951# a_45956_31048# 0.08717f
C17597 _304_.B a_50308_26476# 0.00147f
C17598 a_47732_22504# _421_.B 0.00948f
C17599 a_65220_7908# VPWR 0.20921f
C17600 a_21068_25112# a_21516_25112# 0.01288f
C17601 a_17060_1256# VPWR 0.20348f
C17602 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN 0.0923f
C17603 _452_.CLK _470_.D 0.00123f
C17604 a_67012_4772# VPWR 0.20348f
C17605 a_7516_29383# VPWR 0.32932f
C17606 a_57580_13703# a_57492_13800# 0.28563f
C17607 a_59652_25640# vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I 0.00118f
C17608 _304_.B _404_.A1 0.16131f
C17609 a_5052_17272# a_4940_16839# 0.02634f
C17610 a_43492_27912# a_43008_26795# 0.00263f
C17611 a_44364_16839# a_44276_16936# 0.28563f
C17612 a_35068_1592# VPWR 0.35496f
C17613 a_47388_1592# a_47524_1256# 0.00168f
C17614 a_2812_1159# a_3172_1256# 0.08717f
C17615 _424_.A2 a_49988_21236# 0.36305f
C17616 a_32516_16936# VPWR 0.20348f
C17617 a_47164_12135# a_47612_12135# 0.0131f
C17618 a_64996_12612# a_64972_12135# 0.00172f
C17619 a_4156_1592# a_4604_1592# 0.01288f
C17620 a_8100_1636# a_8188_1592# 0.28563f
C17621 _355_.C a_28054_30196# 0.44398f
C17622 a_3172_29860# a_2812_29816# 0.08707f
C17623 a_15692_25112# a_15692_24679# 0.05841f
C17624 a_19636_25156# a_19612_24679# 0.00172f
C17625 a_43804_30951# VPWR 0.31143f
C17626 a_48420_1636# a_48060_1592# 0.08707f
C17627 a_65332_12232# a_65420_10567# 0.00151f
C17628 _452_.CLK a_45732_18504# 0.00334f
C17629 _304_.B a_53076_24776# 0.00159f
C17630 _311_.A2 a_33724_23111# 0.00137f
C17631 a_46492_15271# a_46628_14180# 0.00154f
C17632 _416_.A1 a_45920_20523# 0.08867f
C17633 a_37844_29860# uo_out[2] 0.01617f
C17634 a_47612_18407# a_47972_18504# 0.08717f
C17635 _448_.Q a_38316_20408# 0.04486f
C17636 a_52764_1159# a_53212_1159# 0.0131f
C17637 a_39236_20072# a_39684_20072# 0.01328f
C17638 _229_.I _252_.B 0.41158f
C17639 a_16948_27912# a_17168_27165# 0.00585f
C17640 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN _248_.B1 0.03719f
C17641 a_67436_18407# VPWR 0.31389f
C17642 a_66116_18884# a_66204_18840# 0.28563f
C17643 _388_.B _324_.C 0.00161f
C17644 a_15156_25156# VPWR 0.20348f
C17645 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I a_58388_17316# 0.00166f
C17646 a_26668_20408# VPWR 0.32016f
C17647 a_15244_27815# a_15156_27912# 0.28563f
C17648 _342_.ZN VPWR 0.45887f
C17649 a_61052_12568# VPWR 0.3185f
C17650 _470_.D a_45577_27509# 0.00207f
C17651 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN a_58836_14180# 0.05215f
C17652 a_40580_26344# _260_.A1 0.03508f
C17653 _424_.B1 _408_.ZN 0.05508f
C17654 a_17803_26841# uio_out[7] 0.01919f
C17655 a_41252_15748# a_41116_15271# 0.00168f
C17656 a_67100_8999# a_67460_9096# 0.08717f
C17657 _316_.ZN a_35044_21640# 0.00654f
C17658 _438_.A2 _441_.B 0.00748f
C17659 a_36076_16839# a_36100_15748# 0.0016f
C17660 a_25436_21543# a_25460_20452# 0.0016f
C17661 a_40644_29480# VPWR 0.01475f
C17662 a_63092_16936# VPWR 0.20703f
C17663 a_18372_28409# VPWR 0.00262f
C17664 a_42596_15368# VPWR 0.23666f
C17665 _300_.A2 a_38676_20452# 0.02529f
C17666 a_23444_22020# a_23892_22020# 0.01328f
C17667 a_41452_16839# a_41900_16839# 0.012f
C17668 a_46044_15271# VPWR 0.33486f
C17669 a_50308_26476# VPWR 0.01026f
C17670 a_2364_16839# VPWR 0.30029f
C17671 a_53572_1256# a_54244_1256# 0.00347f
C17672 a_39460_1256# VPWR 0.20348f
C17673 a_25012_31048# a_24864_29931# 0.00179f
C17674 a_24564_31048# _342_.ZN 0.00164f
C17675 a_29828_26344# VPWR 0.61198f
C17676 a_32828_2727# a_33276_2727# 0.0131f
C17677 a_51980_13703# a_52004_12612# 0.0016f
C17678 a_54132_13800# a_54580_13800# 0.01328f
C17679 _404_.A1 VPWR 1.06751f
C17680 a_37084_17272# a_36972_16839# 0.02634f
C17681 _474_.CLK a_55340_23544# 0.02977f
C17682 a_1020_17272# VPWR 0.30073f
C17683 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN a_54804_16936# 0.0037f
C17684 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN 0.64164f
C17685 _355_.C a_28891_25273# 0.00438f
C17686 a_48868_1636# VPWR 0.2062f
C17687 a_14236_1159# a_14148_1256# 0.28563f
C17688 a_54356_16936# VPWR 0.20637f
C17689 a_4940_12135# a_4852_12232# 0.28563f
C17690 a_11460_1636# a_11100_1592# 0.08707f
C17691 _386_.ZN a_47172_27912# 0.00183f
C17692 a_9668_29860# a_10116_29860# 0.01328f
C17693 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I 0.01363f
C17694 a_32156_17272# a_32604_17272# 0.01288f
C17695 a_36100_17316# a_36188_17272# 0.28563f
C17696 _459_.Q a_30724_26020# 0.27702f
C17697 a_65892_11044# a_65532_11000# 0.08707f
C17698 a_61948_11000# a_62396_11000# 0.01288f
C17699 a_19300_2824# VPWR 0.24564f
C17700 _459_.CLK a_18096_27165# 0.0736f
C17701 a_30795_29977# uo_out[7] 0.00247f
C17702 a_54780_1592# a_55228_1592# 0.012f
C17703 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_61748_26724# 0.00541f
C17704 a_53076_24776# VPWR 0.00405f
C17705 a_59620_23208# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I 0.00565f
C17706 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I 0.00266f
C17707 a_20508_23111# a_20956_23111# 0.01288f
C17708 a_2812_24679# a_3172_24776# 0.08717f
C17709 _342_.ZN a_25296_29977# 0.00271f
C17710 a_52920_22760# _424_.A1 0.00209f
C17711 a_62284_26680# a_62308_26344# 0.00172f
C17712 a_21740_29383# a_21652_29480# 0.28563f
C17713 _459_.CLK _265_.ZN 0.00195f
C17714 a_1020_14136# VPWR 0.30073f
C17715 _474_.CLK a_57044_23588# 0.00183f
C17716 a_27328_25227# VPWR 1.11408f
C17717 _352_.A2 a_25796_24776# 0.01034f
C17718 _304_.A1 a_42154_21236# 0.06526f
C17719 _355_.C _373_.A2 0.10116f
C17720 _459_.CLK a_17472_28363# 0.0177f
C17721 _378_.I a_19412_27912# 0.06666f
C17722 _226_.ZN a_41440_23208# 0.00199f
C17723 a_4068_29480# VPWR 0.22189f
C17724 a_55116_12135# VPWR 0.31547f
C17725 a_37444_15748# a_37084_15704# 0.08707f
C17726 a_33636_2824# a_34084_2824# 0.01328f
C17727 _424_.B1 _412_.A1 0.19878f
C17728 _358_.A3 a_35292_26247# 0.04684f
C17729 a_17484_24679# VPWR 0.29719f
C17730 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN VPWR 0.88009f
C17731 a_59332_29816# a_59744_30352# 0.00705f
C17732 a_43020_16839# a_43044_15748# 0.0016f
C17733 a_24004_21640# a_24116_20452# 0.02666f
C17734 a_40468_25157# VPWR 0.6686f
C17735 a_37892_15748# VPWR 0.21241f
C17736 a_32580_27912# VPWR 0.01438f
C17737 _311_.A2 a_38576_22504# 0.30862f
C17738 _381_.Z a_47700_28292# 0.01297f
C17739 a_1020_9432# a_1468_9432# 0.0131f
C17740 a_3620_9476# a_3260_9432# 0.08717f
C17741 _397_.A2 _390_.ZN 0.81538f
C17742 _303_.ZN a_43156_20452# 0.01509f
C17743 a_46716_14136# a_47164_14136# 0.01288f
C17744 a_50660_14180# a_50748_14136# 0.28563f
C17745 a_45820_18407# VPWR 0.29687f
C17746 _229_.I a_62644_26724# 0.00103f
C17747 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I 0.07319f
C17748 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I a_54692_18884# 0.00206f
C17749 a_49292_16839# VPWR 0.32013f
C17750 _251_.A1 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.0689f
C17751 a_61860_1256# VPWR 0.22423f
C17752 a_28124_30600# uio_out[1] 0.00268f
C17753 a_55140_28292# a_55228_28248# 0.28563f
C17754 a_58924_13703# a_58948_12612# 0.0016f
C17755 _386_.ZN _412_.A1 0.0015f
C17756 a_35040_20937# VPWR 0.00124f
C17757 _475_.Q a_52036_22504# 0.0083f
C17758 _304_.B a_48384_26724# 0.00877f
C17759 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I 0.00502f
C17760 _340_.A2 a_26970_29480# 0.00112f
C17761 a_40644_17272# VPWR 0.35892f
C17762 a_63764_10664# a_63740_9432# 0.0016f
C17763 a_25212_1159# a_25572_1256# 0.08717f
C17764 a_1380_12232# a_1828_12232# 0.01328f
C17765 a_55116_12135# a_55476_12232# 0.08707f
C17766 a_62532_1636# VPWR 0.2085f
C17767 a_17956_1636# a_18404_1636# 0.01328f
C17768 a_1468_21543# VPWR 0.29679f
C17769 a_41048_17341# a_41432_17801# 1.16391f
C17770 _336_.A1 a_28820_24072# 0.39821f
C17771 a_54780_20408# a_54692_18884# 0.00151f
C17772 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN a_58476_18840# 0.00122f
C17773 _451_.Q _441_.A2 0.01845f
C17774 _383_.ZN _404_.A1 0.00906f
C17775 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I a_54804_26724# 0.002f
C17776 a_62084_1636# a_61724_1592# 0.08707f
C17777 a_41700_2824# VPWR 0.21295f
C17778 a_58063_30644# ui_in[4] 0.47495f
C17779 a_19612_23111# a_19524_23208# 0.28563f
C17780 a_23196_24679# a_23108_24776# 0.28563f
C17781 _330_.A1 a_37532_21543# 0.00116f
C17782 a_48420_9476# VPWR 0.20968f
C17783 a_60156_27815# a_60516_27912# 0.0869f
C17784 a_54468_14180# VPWR 0.20348f
C17785 a_4852_18504# a_5300_18504# 0.01328f
C17786 a_35628_18407# a_35988_18504# 0.0869f
C17787 _451_.Q a_40416_18885# 0.13105f
C17788 a_37644_23544# _437_.ZN 0.03072f
C17789 _435_.A3 hold2.I 0.00398f
C17790 a_49204_12232# VPWR 0.23105f
C17791 a_40356_15748# a_40444_15704# 0.28563f
C17792 a_43940_15748# a_44388_15748# 0.01328f
C17793 _284_.A2 _284_.B 0.11399f
C17794 _381_.A2 a_50084_24328# 0.47044f
C17795 _402_.A1 a_43296_28733# 0.03562f
C17796 a_22212_24776# VPWR 0.20862f
C17797 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_54356_26724# 0.03181f
C17798 a_31396_21640# a_31284_20452# 0.02666f
C17799 a_5276_2727# a_5636_2824# 0.08717f
C17800 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN a_57940_20452# 0.03185f
C17801 a_32156_19975# a_32068_20072# 0.28563f
C17802 a_44028_15704# VPWR 0.29679f
C17803 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_63316_23588# 0.05469f
C17804 _402_.A1 _473_.Q 0.01815f
C17805 _384_.ZN _279_.Z 0.26926f
C17806 a_46198_27060# _424_.A2 0.76464f
C17807 _324_.B _302_.Z 0.42847f
C17808 a_65308_19975# VPWR 0.34487f
C17809 _452_.CLK a_39324_26247# 0.00866f
C17810 a_54468_14180# a_54108_14136# 0.08717f
C17811 a_1468_14136# a_1468_13703# 0.05841f
C17812 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I a_64972_26680# 0.02922f
C17813 a_24864_29931# uio_out[2] 0.0034f
C17814 _274_.A3 a_53660_27815# 0.00192f
C17815 a_65868_13703# a_65892_12612# 0.0016f
C17816 a_55228_2727# a_55676_2727# 0.0131f
C17817 a_55924_13800# a_55812_12612# 0.02666f
C17818 a_3708_12568# a_4156_12568# 0.0131f
C17819 _424_.A2 clkbuf_1_0__f_clk.I 0.15102f
C17820 a_31732_25156# _459_.D 0.00422f
C17821 vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN 0.65059f
C17822 _474_.CLK a_54804_24776# 0.00791f
C17823 a_48384_26724# VPWR 0.99377f
C17824 a_37084_26247# VPWR 0.29679f
C17825 a_19140_29612# VPWR 0.0104f
C17826 a_51868_17272# VPWR 0.31547f
C17827 a_1380_9096# a_1380_7908# 0.05841f
C17828 a_4828_1159# VPWR 0.33352f
C17829 a_36636_1159# a_36548_1256# 0.28563f
C17830 _327_.A2 a_44752_18147# 0.1945f
C17831 _459_.Q _337_.ZN 0.16007f
C17832 a_66316_12135# a_66228_12232# 0.28563f
C17833 a_2276_7528# a_2276_6340# 0.05841f
C17834 a_3172_5960# a_3172_4772# 0.05841f
C17835 _451_.Q a_39772_19975# 0.0012f
C17836 _397_.A2 a_48580_27508# 0.00226f
C17837 a_4068_4392# a_4068_3204# 0.05841f
C17838 _346_.B uio_out[5] 0.00177f
C17839 a_32380_21543# VPWR 0.31547f
C17840 a_48196_17316# a_48284_17272# 0.28563f
C17841 a_51780_17316# a_52228_17316# 0.01328f
C17842 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN VPWR 0.73877f
C17843 a_2364_10567# a_2724_10664# 0.08717f
C17844 a_56012_10567# a_56460_10567# 0.012f
C17845 _399_.ZN _399_.A1 0.20418f
C17846 a_64100_2824# VPWR 0.20363f
C17847 a_66788_1636# a_66428_1592# 0.08717f
C17848 a_64188_1592# a_64636_1592# 0.0131f
C17849 _424_.B1 a_51912_20452# 0.00177f
C17850 _272_.A2 _241_.I0 0.00224f
C17851 a_17844_23208# a_18628_23208# 0.00276f
C17852 a_30140_23111# a_30500_23208# 0.08707f
C17853 _281_.ZN a_51240_20452# 0.00171f
C17854 a_59396_9476# VPWR 0.20622f
C17855 a_932_23588# VPWR 0.22176f
C17856 a_62756_2824# a_62620_1592# 0.00154f
C17857 a_26468_2824# a_26556_1159# 0.0027f
C17858 a_24540_21543# a_24988_21543# 0.01288f
C17859 a_62844_14136# VPWR 0.31389f
C17860 a_38788_20072# _330_.A2 0.00191f
C17861 a_39684_20072# a_39268_18840# 0.00238f
C17862 a_2724_3204# VPWR 0.20782f
C17863 a_3260_21543# a_3172_21640# 0.28563f
C17864 _304_.B _435_.A3 0.69363f
C17865 _251_.A1 _230_.I 0.48807f
C17866 _459_.CLK a_27588_26344# 0.03397f
C17867 _474_.CLK _281_.ZN 0.01137f
C17868 _352_.A2 _352_.ZN 0.9017f
C17869 a_12916_31048# a_12892_29816# 0.0016f
C17870 a_3172_11044# VPWR 0.20993f
C17871 a_56036_2824# a_56484_2824# 0.01328f
C17872 _359_.B a_43296_28733# 0.00404f
C17873 a_51332_24072# _384_.A1 0.00563f
C17874 a_63068_19975# a_63428_20072# 0.08717f
C17875 a_66204_18840# a_66092_18407# 0.02634f
C17876 _386_.A4 a_47172_27912# 0.02111f
C17877 _243_.B2 a_58656_27912# 0.00246f
C17878 a_4156_18840# VPWR 0.30552f
C17879 _359_.B a_43828_29860# 0.00252f
C17880 a_44038_21236# a_44290_21236# 0.00184f
C17881 a_56816_26724# VPWR 0.00667f
C17882 a_61836_26680# a_62284_26680# 0.01255f
C17883 a_16700_2727# a_16612_2824# 0.28563f
C17884 _284_.ZN _451_.Q 0.01614f
C17885 a_55140_9476# a_55588_9476# 0.01328f
C17886 a_53796_9476# a_53436_9432# 0.08717f
C17887 _246_.B2 _247_.ZN 0.02009f
C17888 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN VPWR 0.74228f
C17889 _350_.A1 uo_out[2] 0.06089f
C17890 a_48060_14136# a_48060_13703# 0.05841f
C17891 a_52004_14180# a_51980_13703# 0.00172f
C17892 a_62308_14180# a_62756_14180# 0.01328f
C17893 a_4516_20452# a_4604_20408# 0.28563f
C17894 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN a_61188_20072# 0.00636f
C17895 a_62868_13800# a_62756_12612# 0.02666f
C17896 _229_.I vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN 0.32485f
C17897 a_37408_18504# a_38336_18147# 1.16391f
C17898 a_50660_12612# a_50300_12568# 0.08707f
C17899 _275_.ZN a_51457_29861# 0.17673f
C17900 _335_.ZN a_33312_28776# 0.00342f
C17901 a_16948_24776# a_16948_23588# 0.05841f
C17902 a_47612_1159# a_47972_1256# 0.08717f
C17903 _407_.A1 _408_.ZN 0.18156f
C17904 a_27004_1159# VPWR 0.39029f
C17905 a_62868_12232# a_63316_12232# 0.01328f
C17906 a_28036_1636# a_28124_1592# 0.28563f
C17907 a_29604_21640# VPWR 0.20896f
C17908 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_56368_26344# 0.00145f
C17909 a_36636_26247# a_36548_26344# 0.28563f
C17910 _363_.Z a_36100_26724# 0.00329f
C17911 _454_.D a_23284_26724# 0.0018f
C17912 a_53324_10567# a_53236_10664# 0.28563f
C17913 _319_.A3 a_36016_20893# 0.02494f
C17914 a_52452_1636# a_52316_1159# 0.00168f
C17915 a_48508_1592# a_48508_1159# 0.05841f
C17916 a_25420_30345# _340_.ZN 0.00545f
C17917 a_13252_2824# a_13252_1636# 0.05841f
C17918 a_9444_2824# a_9308_1592# 0.00154f
C17919 a_47259_20127# VPWR 0.36713f
C17920 a_1828_22020# VPWR 0.20348f
C17921 _392_.A2 _395_.A1 0.08678f
C17922 _402_.A1 a_44028_27815# 0.01697f
C17923 a_33076_24776# a_33524_24776# 0.01328f
C17924 _304_.B _419_.Z 0.02138f
C17925 a_43008_26795# a_43736_25896# 0.00131f
C17926 a_3260_8999# VPWR 0.30487f
C17927 a_19276_23544# VPWR 0.35601f
C17928 _334_.A1 a_34348_27208# 0.00146f
C17929 a_5388_5863# VPWR 0.35526f
C17930 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.00132f
C17931 a_22352_25987# a_22300_24679# 0.00173f
C17932 a_23196_21543# a_23556_21640# 0.08707f
C17933 a_932_18884# a_1380_18884# 0.01328f
C17934 _435_.A3 VPWR 0.98416f
C17935 a_7068_2727# VPWR 0.31143f
C17936 a_57132_13703# VPWR 0.32388f
C17937 a_52092_11000# VPWR 0.31589f
C17938 a_50076_15704# a_50524_15704# 0.01288f
C17939 a_4964_22020# a_4940_21543# 0.00172f
C17940 _416_.A1 a_52073_30344# 0.00201f
C17941 a_56236_23544# a_56684_23544# 0.0131f
C17942 a_3260_26680# VPWR 0.30487f
C17943 _276_.A2 _416_.A1 0.40829f
C17944 _268_.A1 _274_.ZN 0.51394f
C17945 a_9084_30951# uio_oe[5] 0.00469f
C17946 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I 0.00519f
C17947 a_27588_26724# a_27228_26680# 0.08674f
C17948 _402_.A1 _381_.Z 0.83462f
C17949 _267_.A2 _243_.ZN 0.00122f
C17950 a_20496_26344# VPWR 1.10385f
C17951 a_27676_2727# a_28036_2824# 0.08717f
C17952 a_63316_20452# VPWR 0.19856f
C17953 _304_.B a_55588_28292# 0.00209f
C17954 _311_.A2 a_39536_23588# 0.00125f
C17955 _474_.CLK a_53660_17272# 0.00111f
C17956 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN a_61524_20452# 0.03125f
C17957 a_48708_29816# _383_.A2 0.00375f
C17958 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN a_62308_26344# 0.00491f
C17959 a_62396_26247# _245_.I1 0.06481f
C17960 a_1828_23588# a_1916_23544# 0.28563f
C17961 a_16500_28292# VPWR 0.20815f
C17962 a_2724_4772# a_2812_4728# 0.28563f
C17963 a_1828_6340# a_1916_6296# 0.28563f
C17964 _419_.A4 _397_.Z 0.00135f
C17965 a_55452_14136# a_55564_13703# 0.02634f
C17966 a_3620_3204# a_3708_3160# 0.28563f
C17967 a_18516_20452# a_18964_20452# 0.01328f
C17968 a_57492_23588# a_57132_23544# 0.08717f
C17969 a_52316_27815# a_52764_27815# 0.01255f
C17970 a_1020_1592# VPWR 0.30073f
C17971 a_57156_12612# a_57604_12612# 0.01328f
C17972 a_53572_12612# a_53660_12568# 0.28563f
C17973 _470_.Q _400_.ZN 0.13534f
C17974 _459_.CLK a_19188_25156# 0.00114f
C17975 _258_.I _255_.ZN 0.129f
C17976 _451_.Q a_40580_20452# 0.02998f
C17977 a_24004_24776# a_23892_23588# 0.02666f
C17978 a_5300_18504# a_5388_16839# 0.0027f
C17979 _371_.A2 _336_.A1 0.01726f
C17980 a_49404_1159# VPWR 0.30187f
C17981 a_35008_22461# _316_.A3 0.03442f
C17982 a_39884_27815# uo_out[7] 0.00521f
C17983 a_59036_1159# a_58948_1256# 0.28563f
C17984 _313_.ZN a_33808_23705# 0.00247f
C17985 a_32592_25227# a_33148_25641# 0.8399f
C17986 _438_.A2 _452_.Q 0.05521f
C17987 a_4068_11044# a_4156_11000# 0.28563f
C17988 _459_.Q a_30795_29977# 0.00261f
C17989 a_67012_18884# VPWR 0.20637f
C17990 a_41228_27815# a_41140_27912# 0.28563f
C17991 a_50660_20452# a_51240_20452# 0.00566f
C17992 a_63852_10567# a_64212_10664# 0.08663f
C17993 _311_.A2 a_35616_24776# 0.00911f
C17994 a_50100_10664# a_50548_10664# 0.01328f
C17995 a_35180_18407# a_35204_17316# 0.0016f
C17996 a_18940_1159# a_19388_1159# 0.0131f
C17997 _346_.A2 a_23060_26724# 0.00176f
C17998 _359_.B a_44028_27815# 0.0017f
C17999 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN rst_n 0.00127f
C18000 a_20172_21976# VPWR 0.31589f
C18001 _419_.Z VPWR 1.32267f
C18002 vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I VPWR 0.7761f
C18003 a_61300_15748# a_62084_15748# 0.00276f
C18004 a_34396_21543# a_34308_21640# 0.28563f
C18005 a_31820_23544# VPWR 0.31389f
C18006 a_65072_29860# vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN 0.01698f
C18007 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN _248_.B1 0.6071f
C18008 a_21764_21640# a_22212_21640# 0.01328f
C18009 a_50996_13800# VPWR 0.2093f
C18010 a_29468_2727# VPWR 0.31143f
C18011 _398_.C _281_.ZN 0.36668f
C18012 a_65532_15271# a_65980_15271# 0.01255f
C18013 _399_.A2 VPWR 0.41727f
C18014 _450_.D a_42392_19243# 0.01958f
C18015 _416_.A1 _395_.A1 0.00331f
C18016 a_6396_29816# VPWR 0.3289f
C18017 a_65892_11044# VPWR 0.23512f
C18018 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN _274_.A2 0.11779f
C18019 _324_.B a_43814_21236# 0.00144f
C18020 a_18828_21976# a_18716_21543# 0.02634f
C18021 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I 0.01507f
C18022 _230_.I a_58020_27508# 0.00412f
C18023 _304_.A1 a_37408_23208# 0.00288f
C18024 _304_.B a_55588_27912# 0.00114f
C18025 a_17036_23111# VPWR 0.29679f
C18026 a_42161_24776# _441_.A2 0.00273f
C18027 a_64660_23208# vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I 0.00112f
C18028 a_17396_27912# VPWR 0.20504f
C18029 _260_.A1 _438_.ZN 0.00119f
C18030 a_1468_15271# a_1916_15271# 0.0131f
C18031 _437_.A1 a_37892_26344# 0.01768f
C18032 a_25124_28776# a_26954_28776# 0.00879f
C18033 a_63516_17272# a_63428_15748# 0.00151f
C18034 a_39100_2727# a_39012_2824# 0.28563f
C18035 a_55588_28292# VPWR 0.20348f
C18036 _355_.C a_25867_26841# 0.0289f
C18037 a_19188_23588# a_19636_23588# 0.01328f
C18038 a_15604_23588# a_15692_23544# 0.28563f
C18039 a_58028_20408# a_58476_20408# 0.01222f
C18040 a_19972_1256# a_20420_1256# 0.01328f
C18041 a_64772_9476# a_64412_9432# 0.08717f
C18042 a_66116_9476# a_66564_9476# 0.01328f
C18043 a_66116_7908# a_66204_7864# 0.28563f
C18044 a_5052_4728# a_4940_4295# 0.02634f
C18045 a_65756_4728# a_66204_4728# 0.0131f
C18046 a_67908_4772# a_67996_4728# 0.28563f
C18047 a_64860_6296# a_65308_6296# 0.0131f
C18048 a_67012_6340# a_67100_6296# 0.28563f
C18049 _267_.A2 _258_.ZN 0.0416f
C18050 a_49292_13703# a_49740_13703# 0.01288f
C18051 a_66652_3160# a_67100_3160# 0.0131f
C18052 a_66788_14180# a_66764_13703# 0.00172f
C18053 a_24116_20452# a_24204_20408# 0.28563f
C18054 a_13452_30951# a_14372_31048# 0.00375f
C18055 a_14004_31048# a_13364_31048# 0.00782f
C18056 a_10428_29383# a_10876_29383# 0.0131f
C18057 a_64412_17272# a_64524_16839# 0.02634f
C18058 a_40244_21640# a_40220_20408# 0.0016f
C18059 a_14684_1592# VPWR 0.29679f
C18060 _416_.A1 _442_.ZN 0.59485f
C18061 a_67124_13800# a_67212_12135# 0.00151f
C18062 a_1916_30951# a_2364_30951# 0.0131f
C18063 _274_.A3 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN 0.01316f
C18064 a_49316_31048# vgaringosc.workerclkbuff_notouch_.I 0.00649f
C18065 a_31803_24831# a_32180_23588# 0.0306f
C18066 a_42168_22504# a_42376_22504# 0.00748f
C18067 _244_.Z a_61836_25515# 0.00218f
C18068 a_65668_9096# VPWR 0.21209f
C18069 a_24304_26795# VPWR 1.11491f
C18070 a_67460_5960# VPWR 0.20924f
C18071 a_64660_23588# a_64748_23544# 0.28563f
C18072 a_52004_11044# a_52452_11044# 0.01328f
C18073 a_66004_18504# a_66092_16839# 0.00151f
C18074 a_48420_11044# a_48508_11000# 0.28563f
C18075 a_35540_16936# a_35988_16936# 0.01328f
C18076 a_37756_1592# a_38204_1592# 0.01288f
C18077 a_1380_18504# VPWR 0.20348f
C18078 a_39772_19975# a_40220_19975# 0.01255f
C18079 _441_.A3 _325_.A1 0.00216f
C18080 _355_.B a_28596_26725# 0.11576f
C18081 a_67117_30600# vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.00987f
C18082 a_64188_1592# a_64188_1159# 0.05841f
C18083 a_62508_21976# vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I 0.02646f
C18084 a_65084_30951# rst_n 0.00758f
C18085 a_31820_21976# VPWR 0.31389f
C18086 a_26427_29977# _373_.ZN 0.00351f
C18087 a_46716_30951# a_47164_30951# 0.0131f
C18088 a_39268_18840# a_38644_19368# 0.00587f
C18089 a_4964_12612# VPWR 0.21167f
C18090 _421_.A1 a_47776_20893# 0.00189f
C18091 a_51868_2727# VPWR 0.31143f
C18092 a_2724_26344# a_3172_26344# 0.01328f
C18093 a_62172_18407# a_62084_18504# 0.28563f
C18094 a_17036_26247# a_17396_26344# 0.08717f
C18095 a_66004_16936# a_65980_15271# 0.00134f
C18096 _383_.A2 _402_.A1 0.61786f
C18097 a_20379_29977# VPWR 0.51398f
C18098 a_52876_10567# VPWR 0.33016f
C18099 a_35964_15271# a_36324_15368# 0.08717f
C18100 a_54780_20408# a_55228_20408# 0.01255f
C18101 _447_.Q a_39324_19975# 0.02793f
C18102 a_14708_23208# VPWR 0.22176f
C18103 a_55588_27912# VPWR 0.20844f
C18104 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I a_65668_23208# 0.00569f
C18105 a_47259_20127# a_47504_19759# 0.00232f
C18106 _274_.A1 a_55228_28248# 0.00278f
C18107 _439_.ZN a_40656_23588# 0.00446f
C18108 a_4068_28292# a_4516_28292# 0.01328f
C18109 a_2276_28292# a_1916_28248# 0.08717f
C18110 a_49852_2727# a_50436_2824# 0.01675f
C18111 a_2724_22020# a_2812_21976# 0.28563f
C18112 _424_.A1 a_52652_18407# 0.02054f
C18113 a_66116_17316# a_66204_17272# 0.28563f
C18114 _448_.Q _301_.Z 0.05173f
C18115 _424_.A1 VPWR 1.206f
C18116 a_46180_18504# a_46628_18504# 0.01328f
C18117 a_17844_25156# a_18292_25156# 0.01328f
C18118 a_46268_13703# a_46180_13800# 0.28563f
C18119 _474_.CLK a_53796_30344# 0.00194f
C18120 a_29356_20408# a_29940_20452# 0.01675f
C18121 a_61860_26344# _245_.I1 0.00309f
C18122 a_54244_20452# a_53884_20408# 0.0869f
C18123 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_64660_23588# 0.00188f
C18124 a_33052_16839# a_32964_16936# 0.28563f
C18125 _355_.C a_17148_29383# 0.04948f
C18126 _395_.A2 _284_.A2 0.31527f
C18127 a_22548_31048# a_22560_30288# 0.01402f
C18128 input9.Z _272_.B1 0.00459f
C18129 _218_.ZN _473_.Q 0.00478f
C18130 _419_.Z _424_.B2 0.33339f
C18131 a_28484_1636# VPWR 0.20348f
C18132 a_53412_29480# VPWR 0.00559f
C18133 a_63740_12568# a_64188_12568# 0.01288f
C18134 a_67684_12612# a_67324_12568# 0.08707f
C18135 _264_.B _305_.A2 0.0037f
C18136 a_54132_12232# a_54220_10567# 0.00151f
C18137 a_45060_1636# a_44700_1592# 0.08707f
C18138 a_62284_26680# a_62396_26247# 0.02634f
C18139 _362_.B a_36548_26724# 0.00489f
C18140 a_60940_28248# a_61052_27815# 0.02634f
C18141 _424_.A1 a_54108_21543# 0.00522f
C18142 a_49316_23588# VPWR 0.00471f
C18143 a_15156_26724# a_15244_26680# 0.28563f
C18144 _411_.A2 a_48376_27508# 0.00122f
C18145 a_47636_18884# a_47612_18407# 0.00172f
C18146 _268_.A2 _267_.A2 0.58217f
C18147 a_59652_25640# vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I 0.01344f
C18148 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN a_60212_25156# 0.03424f
C18149 a_41340_1159# a_41788_1159# 0.0131f
C18150 _381_.Z _424_.B1 0.04392f
C18151 _416_.A1 _397_.A1 0.77532f
C18152 _459_.CLK a_31088_30301# 0.00252f
C18153 a_54444_24679# a_54356_24776# 0.28563f
C18154 a_15244_20408# VPWR 0.31143f
C18155 _304_.B input9.Z 0.0632f
C18156 _336_.Z _358_.A2 0.75375f
C18157 a_66004_16936# a_66452_16936# 0.01328f
C18158 _268_.A2 a_53212_29816# 0.2518f
C18159 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I a_51665_30344# 0.004f
C18160 a_54020_12612# VPWR 0.20595f
C18161 _359_.B _383_.A2 0.00893f
C18162 a_9084_29383# a_8996_29480# 0.28563f
C18163 a_7180_30951# uio_oe[7] 0.00326f
C18164 vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN a_67124_20452# 0.00135f
C18165 a_45284_15368# a_45956_15368# 0.00347f
C18166 _444_.D a_36172_24463# 0.22938f
C18167 _424_.B1 a_51540_24776# 0.00638f
C18168 a_46628_10664# VPWR 0.20348f
C18169 a_47388_15271# a_47300_15368# 0.28563f
C18170 a_54804_23588# VPWR 0.20348f
C18171 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN a_52756_29076# 0.01361f
C18172 a_67548_2727# a_67684_1636# 0.00154f
C18173 _324_.C vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN 0.02732f
C18174 a_44276_20072# _325_.ZN 0.00159f
C18175 _245_.I1 a_62404_25156# 0.00122f
C18176 a_36100_26724# a_36188_26680# 0.28563f
C18177 _416_.A2 VPWR 0.45564f
C18178 a_62172_15271# VPWR 0.29679f
C18179 a_48732_15271# a_49180_15271# 0.0131f
C18180 _241_.Z a_56964_26724# 0.23666f
C18181 _386_.ZN _381_.Z 0.13431f
C18182 _229_.I a_59172_26724# 0.00141f
C18183 a_16500_22020# a_16588_21976# 0.28563f
C18184 a_20084_22020# a_20532_22020# 0.01328f
C18185 a_65756_15704# VPWR 0.34793f
C18186 a_23912_27967# VPWR 0.00204f
C18187 a_61276_2727# a_61188_2824# 0.28563f
C18188 a_57492_17316# a_57468_16839# 0.00172f
C18189 _324_.C _402_.A1 0.38502f
C18190 a_45596_30951# a_45508_31048# 0.28563f
C18191 _474_.CLK _274_.ZN 0.42894f
C18192 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN a_64772_26344# 0.02376f
C18193 a_42154_21236# a_42778_21812# 0.10711f
C18194 a_40332_21543# a_40244_21640# 0.28563f
C18195 a_26916_23208# a_27004_21543# 0.00151f
C18196 a_26668_23544# a_27116_23544# 0.01255f
C18197 a_42148_1256# a_42820_1256# 0.00347f
C18198 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN a_59172_23588# 0.00238f
C18199 a_16612_1256# VPWR 0.20348f
C18200 a_64772_7908# VPWR 0.20727f
C18201 a_66564_4772# VPWR 0.20631f
C18202 _287_.A1 uo_out[4] 1.64301f
C18203 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN a_58388_18884# 0.00102f
C18204 a_7068_29383# VPWR 0.32932f
C18205 a_21404_2727# a_21852_2727# 0.0131f
C18206 a_57132_13703# a_57492_13800# 0.08707f
C18207 a_3172_13800# a_3620_13800# 0.01328f
C18208 a_54108_14136# a_54020_12612# 0.00151f
C18209 _336_.Z _355_.ZN 0.40816f
C18210 _355_.B a_28256_25597# 0.01119f
C18211 a_56124_23111# a_56572_23111# 0.01222f
C18212 a_61972_20452# a_62060_20408# 0.28563f
C18213 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I a_61164_20408# 0.00581f
C18214 a_43916_16839# a_44276_16936# 0.08707f
C18215 clkbuf_1_0__f_clk.I hold1.Z 0.03391f
C18216 a_34620_1592# VPWR 0.31011f
C18217 a_2812_1159# a_2724_1256# 0.28563f
C18218 a_59372_10567# a_59396_9476# 0.0016f
C18219 a_49204_10664# a_49092_9476# 0.02666f
C18220 a_32068_16936# VPWR 0.20348f
C18221 a_8100_1636# a_7740_1592# 0.08663f
C18222 a_61052_12568# a_61164_12135# 0.02634f
C18223 a_5052_12568# a_4964_11044# 0.00151f
C18224 _324_.C _243_.A1 0.00589f
C18225 _355_.C a_26427_29977# 0.00167f
C18226 a_21516_23544# a_21404_23111# 0.02634f
C18227 _375_.Z uio_out[6] 0.13131f
C18228 a_2724_29860# a_2812_29816# 0.28563f
C18229 a_6308_29860# a_6756_29860# 0.01328f
C18230 a_3708_17272# a_4156_17272# 0.0131f
C18231 a_58140_11000# a_58588_11000# 0.01288f
C18232 a_43356_30951# VPWR 0.31143f
C18233 a_51556_1636# a_52004_1636# 0.01328f
C18234 a_47972_1636# a_48060_1592# 0.28563f
C18235 _419_.A4 _284_.B 0.14682f
C18236 a_37396_29860# uo_out[2] 0.01651f
C18237 _424_.A2 a_53436_18840# 0.00648f
C18238 _451_.Q _331_.ZN 0.27178f
C18239 a_47612_18407# a_47524_18504# 0.28563f
C18240 a_49316_18504# a_49292_16839# 0.00131f
C18241 a_16948_27912# a_16240_26795# 0.00758f
C18242 a_19860_27912# a_19860_26724# 0.05841f
C18243 _330_.A1 _325_.A1 0.53278f
C18244 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN 0.00127f
C18245 a_32476_29167# _335_.ZN 0.0101f
C18246 a_66116_18884# a_65756_18840# 0.0869f
C18247 a_66988_18407# VPWR 0.31389f
C18248 _319_.A3 _325_.A2 0.18271f
C18249 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN VPWR 0.95403f
C18250 a_14708_25156# VPWR 0.22176f
C18251 a_14796_27815# a_15156_27912# 0.08717f
C18252 a_26220_20408# VPWR 0.32182f
C18253 input9.Z VPWR 0.65168f
C18254 _424_.A1 _424_.B2 0.24467f
C18255 a_24864_29931# VPWR 1.11253f
C18256 _402_.B a_46352_22021# 0.01248f
C18257 a_67684_12612# VPWR 0.21167f
C18258 a_22212_2824# a_22660_2824# 0.01328f
C18259 _447_.Q a_40132_20452# 0.0015f
C18260 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN a_57604_14180# 0.00676f
C18261 _304_.A1 a_42168_22504# 0.01683f
C18262 a_55700_24776# a_56148_24776# 0.01328f
C18263 a_932_9476# VPWR 0.22176f
C18264 a_67100_8999# a_67012_9096# 0.28563f
C18265 a_932_7528# a_932_6340# 0.05841f
C18266 _316_.ZN a_34308_21640# 0.03142f
C18267 a_16500_21640# a_16500_20452# 0.05841f
C18268 a_62644_16936# VPWR 0.20703f
C18269 a_55340_26680# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.00207f
C18270 vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN a_56684_18407# 0.00615f
C18271 _355_.C a_28012_24679# 0.03893f
C18272 a_40196_29480# VPWR 0.01455f
C18273 _300_.A2 a_38228_20452# 0.01196f
C18274 a_42148_15368# VPWR 0.23123f
C18275 _359_.B _324_.C 0.00879f
C18276 a_45372_15271# VPWR 0.32517f
C18277 a_16796_27209# a_17140_26841# 0.00275f
C18278 a_3708_14136# a_4156_14136# 0.0131f
C18279 a_49212_26369# VPWR 0.00941f
C18280 a_41364_16936# a_41340_15704# 0.0016f
C18281 a_45172_16936# a_45284_15748# 0.02666f
C18282 a_1916_16839# VPWR 0.297f
C18283 _437_.A1 uo_out[1] 0.00453f
C18284 a_39012_1256# VPWR 0.22423f
C18285 a_68108_13703# a_68020_13800# 0.28563f
C18286 a_66652_3160# a_66652_2727# 0.05841f
C18287 _474_.CLK a_54892_23544# 0.00744f
C18288 _355_.C a_29184_25597# 0.004f
C18289 a_54892_16839# a_54804_16936# 0.28563f
C18290 a_4964_17316# VPWR 0.21167f
C18291 _294_.A2 a_32380_26247# 0.00294f
C18292 a_13788_1159# a_14148_1256# 0.08717f
C18293 a_53908_16936# VPWR 0.20932f
C18294 a_48420_1636# VPWR 0.20348f
C18295 a_49404_12568# a_49316_11044# 0.00151f
C18296 a_6980_29480# a_7428_29480# 0.01328f
C18297 a_58028_12135# a_58476_12135# 0.01288f
C18298 a_4156_12135# a_4852_12232# 0.01227f
C18299 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I 0.06245f
C18300 a_11012_1636# a_11100_1592# 0.28563f
C18301 a_14596_1636# a_15044_1636# 0.01328f
C18302 a_28820_24072# a_29244_23111# 0.01957f
C18303 a_36100_17316# a_35740_17272# 0.08707f
C18304 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN clk 0.05085f
C18305 a_44164_31048# a_44612_31048# 0.01328f
C18306 _304_.B _411_.A2 0.10984f
C18307 a_65444_11044# a_65532_11000# 0.28563f
C18308 a_18852_2824# VPWR 0.21061f
C18309 a_31088_30301# uo_out[7] 0.00193f
C18310 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN a_63180_26680# 0.01675f
C18311 _459_.CLK a_17803_26841# 0.04514f
C18312 a_59172_23208# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I 0.00163f
C18313 a_2812_24679# a_2724_24776# 0.28563f
C18314 _330_.A1 _327_.A2 0.04086f
C18315 a_20508_24679# a_20956_24679# 0.01288f
C18316 _234_.ZN a_41228_27815# 0.00189f
C18317 a_63740_1159# a_64188_1159# 0.0131f
C18318 a_3260_19975# a_3708_19975# 0.0131f
C18319 a_1828_4392# a_2276_4392# 0.01328f
C18320 _459_.CLK a_41440_28363# 0.01376f
C18321 a_4964_14180# VPWR 0.21167f
C18322 _474_.CLK a_56596_23588# 0.00456f
C18323 a_48420_2824# a_48420_1636# 0.05841f
C18324 a_4940_18407# a_5388_18407# 0.01222f
C18325 _260_.A1 a_40692_21640# 0.00722f
C18326 a_36996_15748# a_37084_15704# 0.28563f
C18327 a_3620_29480# VPWR 0.22347f
C18328 a_33052_15704# a_33500_15704# 0.01288f
C18329 a_54668_12135# VPWR 0.31547f
C18330 _378_.I a_17844_27912# 0.00104f
C18331 _325_.A1 _226_.ZN 1.30671f
C18332 _383_.A2 _386_.ZN 0.03869f
C18333 _358_.A3 a_33396_26344# 0.00187f
C18334 a_23332_26344# a_23780_26344# 0.01328f
C18335 a_17036_24679# VPWR 0.29679f
C18336 _416_.A1 _441_.ZN 0.17537f
C18337 a_40084_25156# VPWR 0.00664f
C18338 a_32132_27912# VPWR 0.01679f
C18339 a_37444_15748# VPWR 0.20622f
C18340 a_48776_20204# a_48888_19243# 0.00259f
C18341 a_3172_9476# a_3260_9432# 0.28563f
C18342 a_26220_21976# a_26668_21976# 0.01288f
C18343 a_48508_18407# a_48956_18407# 0.0131f
C18344 _476_.Q _427_.B2 0.04093f
C18345 _397_.A2 a_48141_29480# 0.00642f
C18346 a_52204_16839# a_52652_16839# 0.0131f
C18347 a_50660_14180# a_50300_14136# 0.08707f
C18348 _303_.ZN a_42728_20452# 0.02291f
C18349 a_52116_16936# a_52228_15748# 0.02666f
C18350 a_48308_16936# a_48284_15704# 0.0016f
C18351 a_44752_18147# VPWR 0.5127f
C18352 _229_.I a_62196_26724# 0.00201f
C18353 _251_.A1 a_56516_26344# 0.30233f
C18354 a_48844_16839# VPWR 0.31857f
C18355 a_20853_30644# uio_out[5] 0.00957f
C18356 _300_.ZN _325_.A1 0.07509f
C18357 a_27668_31048# uio_out[1] 0.08996f
C18358 a_61188_1256# VPWR 0.20968f
C18359 a_64548_1256# a_64996_1256# 0.01328f
C18360 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN 0.63757f
C18361 a_44459_18559# a_44812_17272# 0.00158f
C18362 a_43804_2727# a_44252_2727# 0.0131f
C18363 a_64884_13800# a_65332_13800# 0.01328f
C18364 _475_.Q a_51618_22504# 0.0043f
C18365 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN 0.10606f
C18366 a_39324_17272# VPWR 0.32802f
C18367 _416_.A2 a_47504_19759# 0.00103f
C18368 a_62084_1636# VPWR 0.2085f
C18369 a_25212_1159# a_25124_1256# 0.28563f
C18370 a_55116_12135# a_55028_12232# 0.28563f
C18371 _409_.ZN a_51084_28248# 0.00379f
C18372 _325_.A1 a_44459_18559# 0.00133f
C18373 a_12444_29816# a_12892_29816# 0.01288f
C18374 a_2724_26344# a_2724_25156# 0.05841f
C18375 a_1020_21543# VPWR 0.30073f
C18376 a_41048_17341# a_41536_17636# 0.8399f
C18377 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I clk 0.03932f
C18378 _336_.A1 a_28460_23544# 0.0547f
C18379 _336_.A2 a_29716_23588# 0.00482f
C18380 _411_.A2 VPWR 2.13216f
C18381 a_41252_2824# VPWR 0.2113f
C18382 _386_.A4 _381_.Z 0.45736f
C18383 a_38116_1636# a_37980_1159# 0.00168f
C18384 a_34172_1592# a_34172_1159# 0.05841f
C18385 a_57692_1592# a_58140_1592# 0.01288f
C18386 a_61636_1636# a_61724_1592# 0.28563f
C18387 _294_.ZN a_33776_29123# 0.05474f
C18388 a_31036_23111# a_31484_23111# 0.01288f
C18389 a_19164_23111# a_19524_23208# 0.08707f
C18390 a_22748_24679# a_23108_24776# 0.08707f
C18391 _330_.A1 a_37084_21543# 0.00224f
C18392 a_47972_9476# VPWR 0.20348f
C18393 a_20672_30301# _378_.I 0.00571f
C18394 a_4156_21543# a_4940_21543# 0.00443f
C18395 _343_.A2 _346_.A2 0.11498f
C18396 a_54020_14180# VPWR 0.20348f
C18397 a_60156_27815# a_60068_27912# 0.28563f
C18398 _267_.A1 a_52764_27815# 0.02209f
C18399 _324_.C _424_.B1 0.5006f
C18400 a_35628_18407# a_35540_18504# 0.28563f
C18401 _442_.ZN _431_.A3 0.103f
C18402 a_37196_23544# _437_.ZN 0.01161f
C18403 VPWR ui_in[5] 0.00108f
C18404 _362_.B a_34084_28776# 0.09687f
C18405 _226_.ZN _327_.A2 0.35289f
C18406 a_48420_12232# VPWR 0.20924f
C18407 a_40356_15748# a_39996_15704# 0.08707f
C18408 a_44612_2824# a_45060_2824# 0.01328f
C18409 _267_.ZN a_52292_29480# 0.01909f
C18410 _402_.A1 a_41996_28777# 0.0182f
C18411 _424_.A2 _412_.A1 0.04727f
C18412 a_2812_20408# a_2812_19975# 0.05841f
C18413 a_55140_15748# a_55004_15271# 0.00168f
C18414 a_21764_24776# VPWR 0.20595f
C18415 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_53908_26724# 0.00234f
C18416 a_42996_18840# a_43400_18909# 0.41635f
C18417 _355_.C _346_.B 0.60089f
C18418 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN ui_in[0] 0.00669f
C18419 a_5276_2727# a_5188_2824# 0.28563f
C18420 _454_.Q a_22064_27912# 0.00497f
C18421 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_62196_23588# 0.00751f
C18422 a_38472_30169# _402_.A1 0.00175f
C18423 a_62396_26247# vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN 0.00747f
C18424 a_43580_15704# VPWR 0.29679f
C18425 a_31708_19975# a_32068_20072# 0.08717f
C18426 _250_.A2 a_63105_28293# 0.26368f
C18427 vgaringosc.workerclkbuff_notouch_.I _409_.ZN 0.01417f
C18428 a_47612_9432# a_48060_9432# 0.0131f
C18429 _324_.C _386_.ZN 0.00314f
C18430 a_64860_19975# VPWR 0.33125f
C18431 _304_.A1 a_42996_18840# 0.00148f
C18432 a_52639_30644# uio_in[0] 0.00353f
C18433 a_15132_29383# a_15156_28292# 0.0016f
C18434 a_57156_14180# a_57604_14180# 0.01328f
C18435 a_54020_14180# a_54108_14136# 0.28563f
C18436 a_20172_25112# a_20084_23588# 0.00151f
C18437 _381_.Z _407_.A1 0.01262f
C18438 _268_.A2 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.01398f
C18439 _452_.CLK a_34396_21543# 0.01088f
C18440 _474_.CLK a_54356_24776# 0.0054f
C18441 a_44856_26841# VPWR 0.00204f
C18442 _416_.A1 _389_.ZN 0.04955f
C18443 a_53660_17272# a_53548_16839# 0.02634f
C18444 a_30476_25112# _459_.D 0.09094f
C18445 a_36636_26247# VPWR 0.29679f
C18446 a_51420_17272# VPWR 0.31547f
C18447 _327_.A2 a_44459_18559# 0.02032f
C18448 a_18264_29480# VPWR 0.6182f
C18449 a_51892_12232# a_52340_12232# 0.01328f
C18450 a_36188_1159# a_36548_1256# 0.08717f
C18451 a_4156_1159# VPWR 0.3339f
C18452 a_65868_12135# a_66228_12232# 0.08717f
C18453 a_49740_12135# a_49764_11044# 0.0016f
C18454 a_20732_1592# a_21180_1592# 0.01288f
C18455 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN 0.05837f
C18456 _451_.Q a_39324_19975# 0.0044f
C18457 a_31932_21543# VPWR 0.31547f
C18458 a_48196_17316# a_47836_17272# 0.08707f
C18459 a_20496_26344# a_20980_25156# 0.00263f
C18460 _419_.A4 _474_.Q 1.16338f
C18461 a_52900_15368# a_52876_13703# 0.00144f
C18462 _399_.ZN VPWR 1.12166f
C18463 a_63652_2824# VPWR 0.20348f
C18464 a_2364_10567# a_2276_10664# 0.28563f
C18465 a_66340_1636# a_66428_1592# 0.28563f
C18466 a_30140_23111# a_30052_23208# 0.28563f
C18467 a_24900_24776# a_25348_24776# 0.01328f
C18468 a_67684_24776# VPWR 0.20076f
C18469 a_58948_9476# VPWR 0.20622f
C18470 a_62396_14136# VPWR 0.31389f
C18471 a_2812_21543# a_3172_21640# 0.08717f
C18472 a_2276_3204# VPWR 0.20634f
C18473 a_39236_20072# a_39268_18840# 0.02001f
C18474 a_38788_20072# a_38644_19368# 0.0014f
C18475 _459_.CLK a_27140_26344# 0.02727f
C18476 _355_.C a_28372_23588# 0.01962f
C18477 a_37888_27555# a_38523_27967# 0.02112f
C18478 _411_.A2 a_50068_27508# 0.01066f
C18479 _285_.Z a_40264_30320# 0.50199f
C18480 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I 0.00145f
C18481 a_2724_11044# VPWR 0.20782f
C18482 a_46852_15748# a_47300_15748# 0.01328f
C18483 a_10116_29860# a_9980_29383# 0.00168f
C18484 _229_.I a_61940_29076# 0.07787f
C18485 a_63068_19975# a_62980_20072# 0.28563f
C18486 _427_.A2 a_52452_24072# 0.48718f
C18487 _430_.ZN VPWR 0.64027f
C18488 a_21652_29480# a_22100_29480# 0.01328f
C18489 a_3708_18840# VPWR 0.33374f
C18490 _359_.B a_38472_30169# 0.0037f
C18491 a_16252_2727# a_16612_2824# 0.08717f
C18492 _381_.A2 _284_.B 1.0904f
C18493 a_16700_29816# uio_oe[0] 0.00697f
C18494 a_53348_9476# a_53436_9432# 0.28563f
C18495 a_65556_23588# VPWR 0.21619f
C18496 a_50972_17272# a_50884_15748# 0.00151f
C18497 a_4516_20452# a_4156_20408# 0.08674f
C18498 a_1916_20408# a_2364_20408# 0.0131f
C18499 _448_.Q _330_.ZN 0.00182f
C18500 _304_.A1 _317_.A2 0.00644f
C18501 a_66204_2727# a_66652_2727# 0.01255f
C18502 a_46268_12568# a_46716_12568# 0.01288f
C18503 a_50212_12612# a_50300_12568# 0.28563f
C18504 _334_.A1 a_31920_29480# 0.00405f
C18505 _383_.A2 _386_.A4 0.05557f
C18506 _335_.ZN a_32904_28776# 0.00259f
C18507 a_46628_12232# a_46628_11044# 0.05841f
C18508 a_26556_1159# VPWR 0.33679f
C18509 a_66428_12568# a_66340_11044# 0.00151f
C18510 a_47612_1159# a_47524_1256# 0.28563f
C18511 a_28036_1636# a_27676_1592# 0.08707f
C18512 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I 0.65223f
C18513 a_5300_5960# a_5388_4295# 0.0027f
C18514 a_29156_21640# VPWR 0.20614f
C18515 a_39772_26247# a_40220_26247# 0.01255f
C18516 a_36188_26247# a_36548_26344# 0.0869f
C18517 a_52360_26355# a_53280_26031# 0.00306f
C18518 _454_.D a_23060_26724# 0.00621f
C18519 _363_.Z a_35140_26680# 0.21133f
C18520 a_7516_1159# a_7964_1159# 0.0131f
C18521 a_66764_10567# a_67212_10567# 0.0131f
C18522 _319_.A3 a_34716_20937# 0.00101f
C18523 a_52876_10567# a_53236_10664# 0.08707f
C18524 a_46252_19759# VPWR 0.39698f
C18525 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN 0.03444f
C18526 a_25792_30301# _340_.ZN 0.00195f
C18527 a_28708_23208# a_29156_23208# 0.01328f
C18528 a_1380_22020# VPWR 0.20348f
C18529 _402_.A1 a_43580_27815# 0.03634f
C18530 a_41099_26841# _435_.A3 0.00113f
C18531 a_18828_23544# VPWR 0.32368f
C18532 a_2812_8999# VPWR 0.30213f
C18533 _334_.A1 a_33940_27208# 0.00365f
C18534 a_6620_2727# VPWR 0.31143f
C18535 a_56460_13703# VPWR 0.34572f
C18536 _431_.A3 _435_.ZN 0.00116f
C18537 a_37444_2824# a_37532_1159# 0.0027f
C18538 a_23196_21543# a_23108_21640# 0.28563f
C18539 a_4940_5863# VPWR 0.31945f
C18540 a_1380_21640# a_1828_21640# 0.01328f
C18541 _424_.A2 a_42168_22504# 0.01432f
C18542 _437_.A1 a_38506_26724# 0.00639f
C18543 a_60068_27912# a_60516_27912# 0.01328f
C18544 _317_.A2 _448_.D 0.00328f
C18545 a_51644_11000# VPWR 0.31589f
C18546 _230_.I _255_.I 0.1065f
C18547 a_53572_15748# a_54244_15748# 0.00347f
C18548 a_2364_21976# a_2364_21543# 0.05841f
C18549 a_67012_2824# a_67460_2824# 0.01328f
C18550 a_2812_26680# VPWR 0.30213f
C18551 a_64324_15748# a_64772_15748# 0.01328f
C18552 a_32716_20408# a_32604_19975# 0.02634f
C18553 _384_.A3 _412_.B2 0.20819f
C18554 a_8627_30644# uio_oe[5] 0.00126f
C18555 a_27140_26724# a_27228_26680# 0.28563f
C18556 a_24952_29032# _346_.A2 0.00117f
C18557 a_19524_26344# VPWR 0.23653f
C18558 a_27676_2727# a_27588_2824# 0.28563f
C18559 a_61972_20452# VPWR 0.20547f
C18560 _274_.A2 a_53616_29480# 0.01823f
C18561 _304_.B a_55140_28292# 0.03234f
C18562 _246_.B2 _251_.ZN 0.01044f
C18563 a_1828_23588# a_1468_23544# 0.08717f
C18564 a_3620_23588# a_4068_23588# 0.01328f
C18565 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN a_61076_20452# 0.00409f
C18566 a_58588_9432# a_59036_9432# 0.0131f
C18567 a_16052_28292# VPWR 0.2061f
C18568 _474_.CLK a_53212_17272# 0.00111f
C18569 a_3620_6340# a_4068_6340# 0.01328f
C18570 a_8548_1256# a_8996_1256# 0.01328f
C18571 a_1828_6340# a_1468_6296# 0.08717f
C18572 a_2724_7908# a_3172_7908# 0.01328f
C18573 a_62396_26247# a_62308_26344# 0.28563f
C18574 a_61948_26247# _245_.I1 0.0037f
C18575 a_2724_4772# a_2364_4728# 0.08717f
C18576 a_4516_4772# a_4964_4772# 0.01328f
C18577 a_32268_21976# a_32180_20452# 0.00151f
C18578 a_1020_3160# a_1468_3160# 0.0131f
C18579 a_3620_3204# a_3260_3160# 0.08717f
C18580 a_46356_24072# _402_.B 0.59735f
C18581 _419_.A4 a_46984_23588# 0.04865f
C18582 a_65532_14136# a_65980_14136# 0.01288f
C18583 a_57044_23588# a_57132_23544# 0.28563f
C18584 a_8100_1636# VPWR 0.21493f
C18585 a_63616_31128# _229_.I 0.02469f
C18586 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I 0.12762f
C18587 a_55924_13800# a_56012_12135# 0.00151f
C18588 a_53572_12612# a_53212_12568# 0.08707f
C18589 _459_.CLK a_18740_25156# 0.00249f
C18590 _451_.Q a_40132_20452# 0.00986f
C18591 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN 0.04319f
C18592 _304_.B _397_.A2 0.03457f
C18593 a_44571_26841# _284_.A2 0.01412f
C18594 _305_.A2 a_44038_21236# 0.02323f
C18595 a_48956_1159# VPWR 0.30013f
C18596 _304_.A1 _434_.ZN 0.20137f
C18597 a_58588_1159# a_58948_1256# 0.08717f
C18598 a_33708_22505# _316_.A3 0.00187f
C18599 _337_.A3 _336_.Z 0.00105f
C18600 a_1468_11000# a_1916_11000# 0.0131f
C18601 a_4068_11044# a_3708_11000# 0.08717f
C18602 a_53684_12232# a_53572_11044# 0.02666f
C18603 a_34532_1636# a_34980_1636# 0.01328f
C18604 a_66540_16839# a_66988_16839# 0.01255f
C18605 a_32592_25227# a_33520_25597# 1.16391f
C18606 a_66564_18884# VPWR 0.20919f
C18607 _424_.B1 _281_.A1 0.14674f
C18608 _267_.A1 _258_.I 0.00204f
C18609 a_50660_20452# a_50748_20408# 0.28563f
C18610 _452_.CLK _313_.ZN 0.18905f
C18611 a_40780_27815# a_41140_27912# 0.08674f
C18612 a_64412_29816# a_63952_29480# 0.0011f
C18613 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I 0.0029f
C18614 a_63852_10567# a_63764_10664# 0.28563f
C18615 _275_.A2 a_52292_29480# 0.00206f
C18616 _324_.C _386_.A4 0.00388f
C18617 _331_.ZN a_41536_17636# 0.00393f
C18618 a_19724_21976# VPWR 0.32386f
C18619 a_61300_15748# a_61388_15704# 0.28563f
C18620 a_44270_21790# VPWR 0.00418f
C18621 a_31372_23544# VPWR 0.31389f
C18622 a_29020_2727# VPWR 0.31143f
C18623 a_32068_18884# a_32516_18884# 0.01328f
C18624 a_50548_13800# VPWR 0.2414f
C18625 a_33724_21543# a_34308_21640# 0.01675f
C18626 a_1916_26247# a_2364_26247# 0.0131f
C18627 _398_.C a_46156_25112# 0.04783f
C18628 a_5948_29816# VPWR 0.32916f
C18629 _450_.D a_41188_18840# 0.03203f
C18630 _359_.B a_25124_28776# 0.00146f
C18631 a_65444_11044# VPWR 0.21306f
C18632 _268_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.00142f
C18633 a_53212_2727# a_53348_1636# 0.00154f
C18634 a_16588_23111# VPWR 0.29679f
C18635 _304_.A1 a_36772_23208# 0.05258f
C18636 _304_.B a_55140_27912# 0.00336f
C18637 _223_.I a_32292_26344# 0.00282f
C18638 a_16948_27912# VPWR 0.20418f
C18639 _437_.A1 a_37444_26344# 0.00446f
C18640 _399_.ZN a_51240_23340# 0.00177f
C18641 _417_.A2 _324_.B 0.14437f
C18642 a_47972_31048# _397_.A2 0.00304f
C18643 a_25124_28776# a_26750_28776# 0.01107f
C18644 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN 0.85428f
C18645 a_38428_2727# a_39012_2824# 0.01675f
C18646 a_55140_28292# VPWR 0.20015f
C18647 _355_.C a_26160_27165# 0.08368f
C18648 a_41160_29083# a_41228_27815# 0.00115f
C18649 a_53436_18840# a_54244_18884# 0.00965f
C18650 a_64324_9476# a_64412_9432# 0.28563f
C18651 a_15604_23588# a_15244_23544# 0.08707f
C18652 a_3708_6296# a_3708_5863# 0.05841f
C18653 a_2276_25156# a_2724_25156# 0.01328f
C18654 a_67012_6340# a_66652_6296# 0.08717f
C18655 a_66116_7908# a_65756_7864# 0.08717f
C18656 _267_.A2 a_56572_29383# 0.01227f
C18657 a_2812_7864# a_2812_7431# 0.05841f
C18658 a_63876_20072# a_63876_18884# 0.05841f
C18659 a_67908_4772# a_67548_4728# 0.08663f
C18660 a_62844_14136# a_62956_13703# 0.02634f
C18661 a_24116_20452# a_23756_20408# 0.08717f
C18662 _441_.A3 VPWR 1.43429f
C18663 _448_.Q _303_.ZN 0.02674f
C18664 a_51240_20452# a_51240_19624# 0.00496f
C18665 _294_.ZN a_33720_28776# 0.00144f
C18666 a_13452_30951# a_13364_31048# 0.28563f
C18667 _284_.ZN _441_.A2 0.00479f
C18668 _416_.A1 a_39536_26795# 0.00172f
C18669 a_42154_21236# a_42252_20936# 0.0014f
C18670 a_14236_1592# VPWR 0.29679f
C18671 a_50660_12612# a_50636_12135# 0.00172f
C18672 a_46716_12568# a_46716_12135# 0.05841f
C18673 a_59932_12568# a_60380_12568# 0.012f
C18674 _431_.A3 _441_.ZN 0.18141f
C18675 a_22064_27912# a_22452_27599# 0.00393f
C18676 _285_.Z a_40196_31048# 0.00121f
C18677 _474_.CLK a_51240_19624# 0.00421f
C18678 _424_.ZN a_52884_18884# 0.01167f
C18679 _397_.A2 VPWR 2.8558f
C18680 a_37408_18504# a_38288_18191# 0.00306f
C18681 a_48868_31048# vgaringosc.workerclkbuff_notouch_.I 0.00647f
C18682 a_31803_24831# a_31732_23588# 0.00126f
C18683 a_59260_26680# vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN 0.00155f
C18684 a_65220_9096# VPWR 0.20921f
C18685 a_67012_5960# VPWR 0.20348f
C18686 a_64660_23588# a_64300_23544# 0.0869f
C18687 a_48420_11044# a_48060_11000# 0.08707f
C18688 a_932_18504# VPWR 0.22176f
C18689 a_21600_26725# VPWR 0.63929f
C18690 a_34084_28776# a_35914_28776# 0.00879f
C18691 _251_.A1 _272_.A2 0.57745f
C18692 _452_.CLK _316_.ZN 0.36063f
C18693 _459_.CLK a_21404_24679# 0.00239f
C18694 a_55228_20408# a_55252_20072# 0.00172f
C18695 a_60628_10664# a_61076_10664# 0.01328f
C18696 a_66340_1636# a_66204_1159# 0.00168f
C18697 a_29916_1159# a_30364_1159# 0.0131f
C18698 _251_.A1 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN 0.00169f
C18699 vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I 0.01737f
C18700 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I 0.01861f
C18701 a_22660_24776# a_22748_23111# 0.00151f
C18702 _350_.A1 uo_out[1] 0.00272f
C18703 a_63616_31128# rst_n 0.02625f
C18704 a_4156_26680# a_4156_26247# 0.05841f
C18705 _251_.A1 _244_.Z 0.3468f
C18706 a_31372_21976# VPWR 0.31389f
C18707 _424_.A2 _473_.Q 0.66157f
C18708 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.9187f
C18709 a_26720_30301# _373_.ZN 0.00104f
C18710 _287_.A1 a_33028_27912# 0.00145f
C18711 a_51420_2727# VPWR 0.31143f
C18712 a_32292_21640# a_32740_21640# 0.01328f
C18713 _421_.A1 a_46476_20937# 0.00193f
C18714 a_17036_26247# a_16948_26344# 0.28563f
C18715 a_4516_12612# VPWR 0.20862f
C18716 a_61724_18407# a_62084_18504# 0.08717f
C18717 _369_.ZN a_29680_26724# 0.02375f
C18718 a_33860_15368# a_34532_15368# 0.00347f
C18719 a_18044_29816# VPWR 0.33647f
C18720 a_52428_10567# VPWR 0.31389f
C18721 _455_.Q VPWR 1.7783f
C18722 a_29268_22020# a_29244_21543# 0.00172f
C18723 a_55140_27912# VPWR 0.19737f
C18724 a_25324_21976# a_25436_21543# 0.02634f
C18725 _438_.A2 _261_.ZN 0.35205f
C18726 a_35964_15271# a_35876_15368# 0.28563f
C18727 a_5300_23208# VPWR 0.21406f
C18728 a_65644_23544# a_65668_23208# 0.00172f
C18729 _459_.D a_30588_23111# 0.00179f
C18730 a_37308_15271# a_37756_15271# 0.0131f
C18731 a_48776_20204# a_48964_20204# 0.00257f
C18732 _439_.ZN a_40452_23588# 0.00159f
C18733 a_60401_30300# _250_.ZN 0.00343f
C18734 a_1828_28292# a_1916_28248# 0.28563f
C18735 a_49852_2727# a_49764_2824# 0.28563f
C18736 a_2724_22020# a_2364_21976# 0.08717f
C18737 a_4516_22020# a_4964_22020# 0.01328f
C18738 a_66116_17316# a_65756_17272# 0.0869f
C18739 a_33776_29123# _362_.B 0.22706f
C18740 _346_.A2 a_22636_25112# 0.00111f
C18741 a_64860_8999# a_65308_8999# 0.0131f
C18742 _371_.ZN _371_.A2 0.30042f
C18743 _218_.ZN _281_.A1 0.01827f
C18744 a_65756_7431# a_66204_7431# 0.0131f
C18745 a_30724_1256# a_31396_1256# 0.00347f
C18746 a_21964_23544# a_22548_23588# 0.01675f
C18747 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN 0.00102f
C18748 a_66652_5863# a_67100_5863# 0.0131f
C18749 a_45820_13703# a_46180_13800# 0.08717f
C18750 a_50300_14136# a_50212_12612# 0.00151f
C18751 a_59820_13703# a_60268_13703# 0.01288f
C18752 a_9980_2727# a_10428_2727# 0.0131f
C18753 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.02459f
C18754 a_53796_20452# a_53884_20408# 0.28563f
C18755 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_64212_23588# 0.00887f
C18756 a_67348_18504# a_67460_17316# 0.02666f
C18757 a_61860_26344# a_62308_26344# 0.01328f
C18758 a_32604_16839# a_32964_16936# 0.08717f
C18759 a_2276_10664# a_2276_9476# 0.05841f
C18760 a_47802_26724# _284_.A2 0.0019f
C18761 _395_.A2 a_51048_26680# 0.06668f
C18762 a_28036_1636# VPWR 0.20348f
C18763 a_52964_29480# VPWR 0.00417f
C18764 a_57604_12612# a_57580_12135# 0.00172f
C18765 a_53660_12568# a_53772_12135# 0.02634f
C18766 a_67236_12612# a_67324_12568# 0.28563f
C18767 _304_.B _330_.A1 0.83737f
C18768 a_14004_31048# a_14460_30951# 0.0065f
C18769 _424_.A2 _475_.D 0.14182f
C18770 a_64324_18504# a_64772_18504# 0.01328f
C18771 a_3172_15368# a_3172_14180# 0.05841f
C18772 a_12892_1592# a_12892_1159# 0.05841f
C18773 a_40668_1592# a_41116_1592# 0.01288f
C18774 a_44612_1636# a_44700_1592# 0.28563f
C18775 a_54916_11044# a_55364_11044# 0.01328f
C18776 a_46068_16936# a_46516_16936# 0.01328f
C18777 _362_.B a_36100_26724# 0.06643f
C18778 _279_.Z a_49764_23588# 0.00723f
C18779 a_4940_15271# a_4964_14180# 0.0016f
C18780 _355_.C _351_.A2 0.22719f
C18781 a_15156_26724# a_14796_26680# 0.08674f
C18782 a_48308_23588# VPWR 1.71927f
C18783 _424_.A1 a_53660_21543# 0.01395f
C18784 _397_.A2 _383_.ZN 0.06763f
C18785 a_34084_2824# a_34084_1636# 0.05841f
C18786 _324_.C a_43400_18909# 0.00445f
C18787 vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN 0.01427f
C18788 a_53996_24679# a_54356_24776# 0.0869f
C18789 a_14796_20408# VPWR 0.31538f
C18790 _304_.B a_54432_31128# 0.99911f
C18791 _336_.Z a_29828_26344# 0.11632f
C18792 a_53572_12612# VPWR 0.20595f
C18793 _363_.Z a_33312_28776# 0.00141f
C18794 a_10788_2824# a_11236_2824# 0.01328f
C18795 a_23868_26247# a_24316_26247# 0.012f
C18796 _379_.Z a_18760_29032# 0.03868f
C18797 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN 0.07074f
C18798 a_6723_30644# uio_oe[7] 0.04236f
C18799 a_8636_29383# a_8996_29480# 0.08717f
C18800 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I 0.11229f
C18801 _268_.A2 _276_.A2 0.03145f
C18802 _444_.D a_36544_24419# 0.01723f
C18803 a_46180_10664# VPWR 0.20348f
C18804 a_46940_15271# a_47300_15368# 0.08717f
C18805 a_23980_21976# a_24004_21640# 0.00172f
C18806 a_54356_23588# VPWR 0.18801f
C18807 _351_.A2 a_24636_25641# 0.00386f
C18808 a_47860_21640# VPWR 0.59274f
C18809 a_35616_24776# a_36212_23588# 0.0111f
C18810 _371_.A1 _359_.ZN 0.00713f
C18811 a_61724_15271# VPWR 0.32866f
C18812 a_19035_28409# a_19328_28733# 0.58767f
C18813 a_16500_22020# a_16140_21976# 0.08707f
C18814 a_60828_2727# a_61188_2824# 0.08717f
C18815 a_65308_15704# VPWR 0.33669f
C18816 a_22964_27967# VPWR 0.00246f
C18817 a_45148_30951# a_45508_31048# 0.08717f
C18818 a_64324_15368# a_64996_15368# 0.00347f
C18819 a_57492_18504# a_58164_18504# 0.00347f
C18820 a_16164_1256# VPWR 0.22423f
C18821 a_20620_25112# a_21068_25112# 0.01288f
C18822 a_64324_7908# VPWR 0.22383f
C18823 a_66116_4772# VPWR 0.23643f
C18824 a_57132_13703# a_57044_13800# 0.28563f
C18825 a_6620_29383# VPWR 0.32962f
C18826 a_51576_25896# _412_.ZN 0.0237f
C18827 a_61972_20452# a_61612_20408# 0.08663f
C18828 a_53012_16936# a_52988_15271# 0.00134f
C18829 _336_.Z a_27328_25227# 0.01889f
C18830 a_43916_16839# a_43828_16936# 0.28563f
C18831 a_2364_1159# a_2724_1256# 0.08717f
C18832 a_46940_1592# a_47076_1256# 0.00168f
C18833 a_31620_16936# VPWR 0.20348f
C18834 a_34172_1592# VPWR 0.30352f
C18835 a_46716_12135# a_47164_12135# 0.0131f
C18836 _330_.A1 VPWR 4.43439f
C18837 a_7652_1636# a_7740_1592# 0.28563f
C18838 a_3708_1592# a_4156_1592# 0.01288f
C18839 a_19188_25156# a_19164_24679# 0.00172f
C18840 a_15244_25112# a_15244_24679# 0.05841f
C18841 _355_.C a_26720_30301# 0.00623f
C18842 a_2724_29860# a_2364_29816# 0.08707f
C18843 a_20191_29611# uio_out[6] 0.00277f
C18844 a_42908_30951# VPWR 0.33226f
C18845 a_64884_12232# a_64972_10567# 0.00151f
C18846 vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I a_67212_20408# 0.0014f
C18847 a_47388_1592# a_48060_1592# 0.00544f
C18848 _395_.A2 _381_.A2 0.29893f
C18849 a_46044_15271# a_46180_14180# 0.00154f
C18850 _304_.B _226_.ZN 0.02485f
C18851 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN 0.64529f
C18852 a_36948_29860# uo_out[2] 0.01862f
C18853 a_52316_1159# a_52764_1159# 0.0131f
C18854 a_47164_18407# a_47524_18504# 0.08717f
C18855 a_38788_20072# a_39236_20072# 0.01328f
C18856 a_16500_27912# a_16240_26795# 0.00187f
C18857 a_32848_29123# _335_.ZN 0.00286f
C18858 a_65668_18884# a_65756_18840# 0.28563f
C18859 a_66540_18407# VPWR 0.3163f
C18860 a_5052_25112# VPWR 0.33516f
C18861 a_29268_20452# VPWR 0.21241f
C18862 a_14796_27815# a_14708_27912# 0.28563f
C18863 a_54432_31128# VPWR 0.97717f
C18864 a_67236_12612# VPWR 0.20622f
C18865 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN clk 0.0019f
C18866 a_4604_15704# a_5052_15704# 0.01222f
C18867 _352_.A2 a_30912_27508# 0.00151f
C18868 _447_.Q a_39684_20452# 0.04521f
C18869 a_56260_15368# a_56708_15368# 0.01328f
C18870 VPWR ui_in[0] 0.54647f
C18871 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN a_57156_14180# 0.0011f
C18872 _330_.A2 a_38852_18884# 0.03591f
C18873 _246_.B2 a_60604_27815# 0.00169f
C18874 a_40804_15748# a_40668_15271# 0.00168f
C18875 a_66652_8999# a_67012_9096# 0.08717f
C18876 a_68020_10664# VPWR 0.21538f
C18877 _316_.ZN a_33636_21640# 0.00586f
C18878 a_24988_21543# a_25012_20452# 0.0016f
C18879 a_35628_16839# a_35652_15748# 0.0016f
C18880 _251_.A1 _228_.ZN 0.55049f
C18881 a_39748_29480# VPWR 0.01438f
C18882 a_62196_16936# VPWR 0.20703f
C18883 a_41476_15368# VPWR 0.21356f
C18884 a_22996_22020# a_23444_22020# 0.01328f
C18885 _474_.CLK vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.04551f
C18886 _294_.A2 _287_.A1 0.86912f
C18887 a_44924_15271# VPWR 0.29679f
C18888 a_41004_16839# a_41452_16839# 0.01288f
C18889 a_1468_16839# VPWR 0.29679f
C18890 a_48988_26369# VPWR 0.00541f
C18891 a_38340_1256# VPWR 0.20968f
C18892 a_53124_1256# a_53572_1256# 0.01328f
C18893 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN 0.00218f
C18894 a_53684_13800# a_54132_13800# 0.01328f
C18895 a_32380_2727# a_32828_2727# 0.0131f
C18896 a_67660_13703# a_68020_13800# 0.08717f
C18897 a_51532_13703# a_51556_12612# 0.0016f
C18898 a_36636_17272# a_36524_16839# 0.02634f
C18899 a_58388_17316# a_58836_17316# 0.01328f
C18900 _324_.C _250_.C 0.00183f
C18901 a_54444_16839# a_54804_16936# 0.08663f
C18902 _474_.CLK a_54444_23544# 0.00332f
C18903 a_4516_17316# VPWR 0.20862f
C18904 _294_.A2 a_31932_26247# 0.03077f
C18905 _355_.C a_27884_25641# 0.03443f
C18906 a_47972_1636# VPWR 0.22423f
C18907 a_53460_16936# VPWR 0.20665f
C18908 a_13788_1159# a_13700_1256# 0.28563f
C18909 a_4156_12135# a_4068_12232# 0.28563f
C18910 a_11012_1636# a_10652_1592# 0.08707f
C18911 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN a_65644_23544# 0.0195f
C18912 a_25936_25597# a_25884_24679# 0.00818f
C18913 a_9220_29860# a_9668_29860# 0.01328f
C18914 a_35652_17316# a_35740_17272# 0.28563f
C18915 a_31708_17272# a_32156_17272# 0.01288f
C18916 a_65444_11044# a_65084_11000# 0.08707f
C18917 a_61500_11000# a_61948_11000# 0.01288f
C18918 a_29788_30345# uo_out[7] 0.01407f
C18919 a_54332_1592# a_54780_1592# 0.01288f
C18920 a_63092_26724# a_63180_26680# 0.28563f
C18921 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN a_62732_26680# 0.00379f
C18922 _459_.CLK a_15244_26680# 0.01626f
C18923 a_18404_2824# VPWR 0.20839f
C18924 vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I VPWR 0.75512f
C18925 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I a_63876_20072# 0.00235f
C18926 a_52988_15271# a_53124_14180# 0.00154f
C18927 _226_.ZN VPWR 0.76666f
C18928 a_20060_23111# a_20508_23111# 0.01288f
C18929 _459_.CLK _352_.ZN 0.09834f
C18930 _416_.A2 a_47768_20569# 0.00114f
C18931 a_2364_24679# a_2724_24776# 0.08717f
C18932 _234_.ZN a_40780_27815# 0.03487f
C18933 a_61836_26680# a_61860_26344# 0.00172f
C18934 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN a_64772_18884# 0.00104f
C18935 a_60940_28248# a_60964_27912# 0.00172f
C18936 vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN a_56596_17316# 0.00622f
C18937 a_4516_14180# VPWR 0.20862f
C18938 _330_.A1 a_50068_27508# 0.34297f
C18939 _474_.CLK a_56148_23588# 0.00983f
C18940 hold1.Z a_42168_22504# 0.01556f
C18941 a_36996_15748# a_36636_15704# 0.08707f
C18942 a_3172_29480# VPWR 0.20993f
C18943 _390_.ZN a_51084_28248# 0.018f
C18944 a_54220_12135# VPWR 0.31547f
C18945 _304_.B _274_.A1 0.05061f
C18946 vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I 0.68196f
C18947 a_33188_2824# a_33636_2824# 0.01328f
C18948 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN 0.01509f
C18949 a_16588_24679# VPWR 0.29679f
C18950 _300_.ZN VPWR 0.65517f
C18951 _294_.A2 _293_.A2 0.14738f
C18952 a_42572_16839# a_42596_15748# 0.0016f
C18953 a_23556_21640# a_23668_20452# 0.02666f
C18954 a_36996_15748# VPWR 0.20622f
C18955 a_39860_25156# VPWR 0.01378f
C18956 _260_.ZN a_44270_21790# 0.00195f
C18957 a_3172_9476# a_2812_9432# 0.08717f
C18958 _359_.B a_34084_28776# 0.01387f
C18959 _470_.Q a_47700_28292# 0.01356f
C18960 a_29716_22020# a_30388_22020# 0.00347f
C18961 _303_.ZN a_42460_20452# 0.03828f
C18962 a_54804_20072# a_54692_18884# 0.02666f
C18963 a_44459_18559# VPWR 0.37472f
C18964 a_50212_14180# a_50300_14136# 0.28563f
C18965 a_46268_14136# a_46716_14136# 0.01288f
C18966 _452_.CLK a_45172_17316# 0.00679f
C18967 _229_.I a_61748_26724# 0.00207f
C18968 a_48396_16839# VPWR 0.31556f
C18969 a_27004_30951# uio_out[1] 0.02833f
C18970 a_60740_1256# VPWR 0.20348f
C18971 a_48420_13800# a_48420_12612# 0.05841f
C18972 a_58476_13703# a_58500_12612# 0.0016f
C18973 _460_.Q a_35818_29860# 0.00447f
C18974 _475_.Q a_51414_22504# 0.00487f
C18975 a_35723_20569# VPWR 0.37162f
C18976 a_40040_17675# VPWR 0.69555f
C18977 _237_.A1 _246_.B2 0.70937f
C18978 a_61636_1636# VPWR 0.20847f
C18979 a_63316_10664# a_63292_9432# 0.0016f
C18980 a_24764_1159# a_25124_1256# 0.08717f
C18981 a_932_12232# a_1380_12232# 0.01328f
C18982 a_17508_1636# a_17956_1636# 0.01328f
C18983 a_54668_12135# a_55028_12232# 0.08707f
C18984 _325_.A1 a_43452_18191# 0.04143f
C18985 _355_.ZN a_26548_24372# 0.00153f
C18986 a_15940_29860# a_16612_29860# 0.00347f
C18987 a_52852_24372# clk 0.01639f
C18988 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I a_65108_23588# 0.03128f
C18989 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN 0.00241f
C18990 a_54332_20408# a_54244_18884# 0.00151f
C18991 _336_.A2 a_28820_24072# 0.50373f
C18992 _304_.B a_44302_23588# 0.00132f
C18993 _336_.A1 a_28012_23544# 0.00223f
C18994 a_55140_27912# a_55252_26724# 0.02666f
C18995 a_40804_2824# VPWR 0.2085f
C18996 a_61636_1636# a_61276_1592# 0.08707f
C18997 _294_.ZN a_33483_29535# 0.05929f
C18998 a_19164_23111# a_19076_23208# 0.28563f
C18999 _330_.A1 a_36636_21543# 0.00448f
C19000 a_22748_24679# a_22660_24776# 0.28563f
C19001 a_4852_24776# a_5300_24776# 0.01328f
C19002 _305_.A2 _302_.Z 0.03805f
C19003 a_47524_9476# VPWR 0.20348f
C19004 a_20379_29977# _378_.I 0.00379f
C19005 a_53572_14180# VPWR 0.20348f
C19006 a_4068_18504# a_4852_18504# 0.00276f
C19007 a_35180_18407# a_35540_18504# 0.0869f
C19008 _388_.B _393_.ZN 0.05184f
C19009 _397_.A2 a_49112_29885# 0.0013f
C19010 a_45904_30180# a_46316_29977# 0.00275f
C19011 a_36748_23544# _437_.ZN 0.00482f
C19012 a_43492_15748# a_43940_15748# 0.01328f
C19013 _274_.A1 VPWR 1.18324f
C19014 a_47972_12232# VPWR 0.20348f
C19015 a_39908_15748# a_39996_15704# 0.28563f
C19016 _398_.C _402_.ZN 0.00253f
C19017 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN a_55700_25156# 0.00589f
C19018 a_56516_26344# vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN 0.00762f
C19019 _402_.A1 a_42368_28733# 0.01701f
C19020 _355_.C a_31124_25156# 0.01436f
C19021 a_21316_24776# VPWR 0.20595f
C19022 a_4964_20452# a_4940_19975# 0.00172f
C19023 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN a_58500_21640# 0.00133f
C19024 _411_.A2 _407_.ZN 0.30875f
C19025 _331_.ZN a_40416_18885# 0.13108f
C19026 _250_.ZN a_60852_28292# 0.02f
C19027 a_30948_21640# a_30836_20452# 0.02666f
C19028 a_22636_28248# _454_.D 0.00799f
C19029 a_4828_2727# a_5188_2824# 0.08717f
C19030 a_43132_15704# VPWR 0.30179f
C19031 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_61748_23588# 0.00122f
C19032 a_31708_19975# a_31620_20072# 0.28563f
C19033 _390_.ZN a_52068_29480# 0.0013f
C19034 _250_.A2 a_62503_28293# 0.04853f
C19035 vgaringosc.workerclkbuff_notouch_.I a_49496_30345# 0.01533f
C19036 a_39684_26344# _260_.A2 0.00129f
C19037 a_52415_31220# uio_in[0] 0.06218f
C19038 a_64412_19975# VPWR 0.32034f
C19039 _350_.A1 _362_.ZN 0.0021f
C19040 a_54020_14180# a_53660_14136# 0.08717f
C19041 a_1020_14136# a_1020_13703# 0.05841f
C19042 _452_.CLK _438_.A2 0.00461f
C19043 _300_.ZN a_40452_22504# 0.00108f
C19044 uio_in[0] ui_in[7] 0.06312f
C19045 _350_.A2 uo_out[6] 0.04103f
C19046 _330_.A1 a_44744_26355# 0.00254f
C19047 _452_.CLK a_33724_21543# 0.05929f
C19048 a_65420_13703# a_65444_12612# 0.0016f
C19049 a_54780_2727# a_55228_2727# 0.0131f
C19050 a_55476_13800# a_55364_12612# 0.02666f
C19051 a_3260_12568# a_3708_12568# 0.0131f
C19052 _474_.CLK a_53908_24776# 0.00309f
C19053 a_43908_26841# VPWR 0.00246f
C19054 _416_.A1 a_45484_28248# 0.01676f
C19055 a_30388_25156# _459_.D 0.00822f
C19056 _398_.C a_54444_23544# 0.00127f
C19057 a_36188_26247# VPWR 0.29679f
C19058 a_50972_17272# VPWR 0.31848f
C19059 a_17786_29480# VPWR 0.01552f
C19060 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I VPWR 0.72731f
C19061 _327_.A2 a_43452_18191# 0.00164f
C19062 a_3708_1159# VPWR 0.33167f
C19063 a_36188_1159# a_36100_1256# 0.28563f
C19064 a_65868_12135# a_65780_12232# 0.28563f
C19065 a_1828_7528# a_1828_6340# 0.05841f
C19066 _451_.Q a_38876_19975# 0.0026f
C19067 a_3620_4392# a_3620_3204# 0.05841f
C19068 a_2724_5960# a_2724_4772# 0.05841f
C19069 _474_.CLK a_56596_29861# 0.00112f
C19070 a_31484_21543# VPWR 0.31547f
C19071 a_62560_25112# vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN 0.01708f
C19072 a_44302_23588# VPWR 0.0044f
C19073 a_51332_17316# a_51780_17316# 0.01328f
C19074 _478_.D a_54088_22895# 0.02417f
C19075 a_47748_17316# a_47836_17272# 0.28563f
C19076 a_55564_10567# a_56012_10567# 0.01288f
C19077 a_1916_10567# a_2276_10664# 0.08717f
C19078 a_63740_1592# a_64188_1592# 0.0131f
C19079 a_66340_1636# a_65980_1592# 0.08717f
C19080 a_63204_2824# VPWR 0.20839f
C19081 a_29692_23111# a_30052_23208# 0.08707f
C19082 a_17396_23208# a_17844_23208# 0.01328f
C19083 a_2812_21543# a_2724_21640# 0.28563f
C19084 _459_.CLK _345_.A2 0.09424f
C19085 a_58500_9476# VPWR 0.21691f
C19086 a_24092_21543# a_24540_21543# 0.01288f
C19087 a_61948_14136# VPWR 0.31389f
C19088 a_1828_3204# VPWR 0.20348f
C19089 a_62308_2824# a_62172_1592# 0.00154f
C19090 a_26020_2824# a_26108_1159# 0.0027f
C19091 _324_.C _424_.A2 0.74593f
C19092 _459_.CLK a_26746_26344# 0.00219f
C19093 a_37888_27555# a_37516_27599# 0.10745f
C19094 _281_.A1 a_51877_21236# 0.00498f
C19095 _476_.Q a_52452_21236# 0.00999f
C19096 a_2276_11044# VPWR 0.20634f
C19097 _229_.I a_59572_29076# 0.00266f
C19098 a_55588_2824# a_56036_2824# 0.01328f
C19099 a_62620_19975# a_62980_20072# 0.08717f
C19100 a_47483_20569# VPWR 0.37397f
C19101 a_51332_24072# a_52452_24072# 0.04556f
C19102 _250_.ZN _238_.I 0.11516f
C19103 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN 0.00101f
C19104 a_38616_24328# VPWR 0.30455f
C19105 a_3260_18840# VPWR 0.30487f
C19106 a_52316_27815# _412_.A1 0.00154f
C19107 _424_.A2 _416_.ZN 0.00219f
C19108 a_16252_2727# a_16164_2824# 0.28563f
C19109 _363_.Z a_32476_29167# 0.01615f
C19110 a_53348_9476# a_52988_9432# 0.08717f
C19111 a_54692_9476# a_55140_9476# 0.01328f
C19112 a_65108_23588# VPWR 0.212f
C19113 a_61860_14180# a_62308_14180# 0.01328f
C19114 a_51556_14180# a_51532_13703# 0.00172f
C19115 _397_.A4 _284_.A2 0.02005f
C19116 a_47612_14136# a_47612_13703# 0.05841f
C19117 _399_.A1 _395_.A3 0.13921f
C19118 a_4068_20452# a_4156_20408# 0.28563f
C19119 _304_.A1 a_36148_21976# 0.16735f
C19120 _246_.B2 _242_.Z 0.00475f
C19121 a_5300_13800# a_5388_12135# 0.0027f
C19122 a_50212_12612# a_49852_12568# 0.08707f
C19123 a_62420_13800# a_62308_12612# 0.02666f
C19124 a_16500_24776# a_16500_23588# 0.05841f
C19125 a_26108_1159# VPWR 0.33411f
C19126 a_47164_1159# a_47524_1256# 0.08717f
C19127 a_62420_12232# a_62868_12232# 0.01328f
C19128 a_27588_1636# a_27676_1592# 0.28563f
C19129 a_31172_1636# a_31620_1636# 0.01328f
C19130 a_28708_21640# VPWR 0.20614f
C19131 a_36188_26247# a_36100_26344# 0.28563f
C19132 uio_oe[6] uio_oe[5] 0.06081f
C19133 _319_.A3 a_35088_20893# 0.00267f
C19134 a_52876_10567# a_52788_10664# 0.28563f
C19135 a_48060_1592# a_48060_1159# 0.05841f
C19136 a_52004_1636# a_51868_1159# 0.00168f
C19137 a_12804_2824# a_12804_1636# 0.05841f
C19138 a_8996_2824# a_8860_1592# 0.00154f
C19139 _229_.I _257_.B 0.00775f
C19140 a_46624_19715# VPWR 0.18835f
C19141 a_932_22020# VPWR 0.22176f
C19142 _402_.A1 a_43132_27815# 0.00708f
C19143 _495_.I a_42368_28733# 0.00503f
C19144 a_18380_23544# VPWR 0.3356f
C19145 _373_.A2 _350_.A2 0.02446f
C19146 a_4156_5863# VPWR 0.3269f
C19147 a_2364_8999# VPWR 0.30029f
C19148 a_22748_21543# a_23108_21640# 0.08707f
C19149 a_56012_13703# VPWR 0.31594f
C19150 a_6172_2727# VPWR 0.31143f
C19151 a_33188_25940# VPWR 0.81432f
C19152 _230_.I a_60401_30300# 0.00179f
C19153 a_51196_11000# VPWR 0.31589f
C19154 a_53572_15748# a_53660_15704# 0.28563f
C19155 _474_.CLK _384_.ZN 0.02683f
C19156 a_49628_15704# a_50076_15704# 0.01288f
C19157 _350_.A1 _287_.A2 0.08405f
C19158 a_2364_26680# VPWR 0.30029f
C19159 a_55788_23544# a_56236_23544# 0.0131f
C19160 _281_.ZN _421_.B 0.0078f
C19161 a_19076_26344# VPWR 0.21778f
C19162 _402_.A1 _470_.Q 1.71307f
C19163 _275_.A2 vgaringosc.workerclkbuff_notouch_.I 0.03613f
C19164 _419_.A4 a_47802_26724# 0.02854f
C19165 a_27004_2727# a_27588_2824# 0.01675f
C19166 a_61524_20452# VPWR 0.20697f
C19167 _274_.A2 a_53412_29480# 0.00259f
C19168 _474_.CLK a_52764_17272# 0.00111f
C19169 a_15604_28292# VPWR 0.20703f
C19170 a_1380_23588# a_1468_23544# 0.28563f
C19171 a_1380_6340# a_1468_6296# 0.28563f
C19172 a_61948_26247# a_62308_26344# 0.08663f
C19173 _400_.ZN _284_.B 0.11488f
C19174 a_3172_3204# a_3260_3160# 0.28563f
C19175 a_2276_4772# a_2364_4728# 0.28563f
C19176 a_55004_14136# a_55116_13703# 0.02634f
C19177 a_17932_20408# a_18516_20452# 0.01675f
C19178 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I a_56964_26724# 0.00341f
C19179 a_57044_23588# a_56684_23544# 0.08717f
C19180 a_62532_30736# _229_.I 0.28728f
C19181 a_7652_1636# VPWR 0.2085f
C19182 a_53124_12612# a_53212_12568# 0.28563f
C19183 a_56708_12612# a_57156_12612# 0.01328f
C19184 _459_.CLK a_18292_25156# 0.00251f
C19185 _334_.A1 uo_out[6] 0.52738f
C19186 _398_.C a_53908_24776# 0.00712f
C19187 a_44864_27165# _284_.A2 0.01476f
C19188 _451_.Q a_39684_20452# 0.00142f
C19189 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I 0.0944f
C19190 _393_.A1 VPWR 0.29877f
C19191 a_58588_1159# a_58500_1256# 0.28563f
C19192 a_23556_24776# a_23444_23588# 0.02666f
C19193 a_4852_18504# a_4940_16839# 0.00151f
C19194 a_34080_22461# _316_.A3 0.00163f
C19195 _316_.ZN a_33584_22137# 0.00242f
C19196 _305_.A2 a_43814_21236# 0.00303f
C19197 _371_.A2 _336_.A2 0.01404f
C19198 a_48508_1159# VPWR 0.29679f
C19199 a_38523_27967# uo_out[7] 0.0021f
C19200 a_3620_11044# a_3708_11000# 0.28563f
C19201 a_66116_18884# VPWR 0.2393f
C19202 a_50660_20452# a_50300_20408# 0.08674f
C19203 _452_.CLK a_33376_23659# 0.07458f
C19204 a_40780_27815# a_40692_27912# 0.28563f
C19205 a_36188_25112# a_36172_24463# 0.0019f
C19206 a_49652_10664# a_50100_10664# 0.01328f
C19207 a_18492_1159# a_18940_1159# 0.0131f
C19208 a_63404_10567# a_63764_10664# 0.08707f
C19209 a_34732_18407# a_34756_17316# 0.0016f
C19210 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I 0.72755f
C19211 _275_.A2 a_52068_29480# 0.00725f
C19212 a_57492_23588# vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN 0.0042f
C19213 a_19276_21976# VPWR 0.35698f
C19214 _365_.ZN a_36116_29167# 0.00122f
C19215 _331_.ZN a_41048_17341# 0.00111f
C19216 a_61300_15748# a_60940_15704# 0.08674f
C19217 a_30924_23544# VPWR 0.31389f
C19218 a_21316_21640# a_21764_21640# 0.01328f
C19219 a_28572_2727# VPWR 0.31143f
C19220 a_33724_21543# a_33636_21640# 0.28563f
C19221 a_50100_13800# VPWR 0.21427f
C19222 _264_.B hold2.I 0.24137f
C19223 _398_.C a_46068_25156# 0.0038f
C19224 _384_.A3 _281_.ZN 1.05126f
C19225 _279_.Z _399_.A2 0.65239f
C19226 _397_.A1 _282_.ZN 0.21951f
C19227 a_46580_23588# VPWR 0.00405f
C19228 a_65084_15271# a_65532_15271# 0.01255f
C19229 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I VPWR 1.01326f
C19230 a_5500_29816# VPWR 0.32965f
C19231 a_64996_11044# VPWR 0.2109f
C19232 _304_.B a_53572_27912# 0.01644f
C19233 a_16140_23111# VPWR 0.29679f
C19234 _223_.I a_31844_26344# 0.00191f
C19235 _304_.A1 a_36288_23208# 0.00674f
C19236 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I 0.00671f
C19237 a_1020_15271# a_1468_15271# 0.0131f
C19238 a_16500_27912# VPWR 0.20374f
C19239 _437_.A1 a_36996_26344# 0.0022f
C19240 a_63068_17272# a_62980_15748# 0.00151f
C19241 a_25124_28776# a_26556_28776# 0.01047f
C19242 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN a_65668_23208# 0.00193f
C19243 a_59172_23208# a_59620_23208# 0.01328f
C19244 a_38428_2727# a_38340_2824# 0.28563f
C19245 _355_.C a_24860_27209# 0.01011f
C19246 _334_.A1 uo_out[5] 0.00854f
C19247 a_65668_7908# a_65756_7864# 0.28563f
C19248 a_67460_7908# a_67908_7908# 0.01328f
C19249 a_18740_23588# a_19188_23588# 0.01328f
C19250 a_15156_23588# a_15244_23544# 0.28563f
C19251 a_4964_7908# a_4940_7431# 0.00172f
C19252 a_19300_1256# a_19972_1256# 0.00347f
C19253 a_30724_26020# _358_.A2 0.04413f
C19254 a_65668_9476# a_66116_9476# 0.01328f
C19255 a_63740_9432# a_64412_9432# 0.00544f
C19256 a_64412_6296# a_64860_6296# 0.0131f
C19257 a_66564_6340# a_66652_6296# 0.28563f
C19258 a_55252_20072# vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I 0.00847f
C19259 a_65308_4728# a_65756_4728# 0.0131f
C19260 a_67460_4772# a_67548_4728# 0.28563f
C19261 a_48508_13703# a_49292_13703# 0.00443f
C19262 a_66204_3160# a_66652_3160# 0.0131f
C19263 a_66340_14180# a_66316_13703# 0.00172f
C19264 _459_.Q a_33148_25641# 0.00769f
C19265 a_23668_20452# a_23756_20408# 0.28563f
C19266 a_9980_29383# a_10428_29383# 0.0131f
C19267 a_63964_17272# a_64076_16839# 0.02634f
C19268 a_13004_30951# a_13364_31048# 0.08674f
C19269 _324_.C a_50197_28776# 0.00999f
C19270 a_13788_1592# VPWR 0.29679f
C19271 a_1468_30951# a_1916_30951# 0.0131f
C19272 a_66676_13800# a_66764_12135# 0.00151f
C19273 a_63404_20408# a_63516_19975# 0.02634f
C19274 _359_.B a_33776_29123# 0.04979f
C19275 a_48420_31048# vgaringosc.workerclkbuff_notouch_.I 0.0066f
C19276 a_38971_18559# a_39256_18559# 0.00277f
C19277 _244_.Z a_60084_25640# 0.00197f
C19278 a_47972_11044# a_48060_11000# 0.28563f
C19279 a_18088_26841# VPWR 0.00195f
C19280 a_64772_9096# VPWR 0.20727f
C19281 a_51556_11044# a_52004_11044# 0.01328f
C19282 _441_.A3 a_39780_22805# 0.00492f
C19283 a_66564_5960# VPWR 0.20631f
C19284 a_37308_1592# a_37756_1592# 0.01288f
C19285 a_35092_16936# a_35540_16936# 0.01328f
C19286 _452_.CLK a_33152_22091# 0.1008f
C19287 a_64212_23588# a_64300_23544# 0.28563f
C19288 a_34084_28776# a_35710_28776# 0.01107f
C19289 input9.Z _274_.A2 0.00219f
C19290 _424_.A2 _281_.A1 0.14759f
C19291 _459_.CLK a_20956_24679# 0.00239f
C19292 a_39324_19975# a_39772_19975# 0.01255f
C19293 a_61188_20072# vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I 0.00102f
C19294 a_63740_1592# a_63740_1159# 0.05841f
C19295 _383_.ZN _393_.A1 0.18148f
C19296 _330_.A1 _311_.Z 0.35274f
C19297 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN a_58588_21543# 0.00577f
C19298 vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.07007f
C19299 a_30924_21976# VPWR 0.31389f
C19300 a_56404_27208# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.00336f
C19301 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_56516_26344# 0.03736f
C19302 _268_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN 0.02744f
C19303 _304_.B _264_.B 0.00314f
C19304 _287_.A1 a_32580_27912# 0.00269f
C19305 a_46044_30951# a_46716_30951# 0.00544f
C19306 _325_.A1 _325_.A2 2.30175f
C19307 a_4068_12612# VPWR 0.2157f
C19308 _247_.B a_59620_27208# 0.41959f
C19309 _421_.A1 a_46848_20893# 0.0013f
C19310 a_50972_2727# VPWR 0.31444f
C19311 a_2276_26344# a_2724_26344# 0.01328f
C19312 _230_.I vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN 0.27837f
C19313 a_16588_26247# a_16948_26344# 0.08717f
C19314 _250_.ZN VPWR 0.35315f
C19315 a_61724_18407# a_61636_18504# 0.28563f
C19316 a_65332_16936# a_65532_15271# 0.00119f
C19317 a_17596_29816# VPWR 0.31278f
C19318 _301_.A1 _317_.A2 0.12243f
C19319 a_51980_10567# VPWR 0.31389f
C19320 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN 0.73388f
C19321 a_35516_15271# a_35876_15368# 0.08717f
C19322 a_24392_28248# VPWR 0.31522f
C19323 a_54332_20408# a_54780_20408# 0.01255f
C19324 _384_.ZN _398_.C 0.11957f
C19325 a_53572_27912# VPWR 0.21088f
C19326 a_4852_23208# VPWR 0.22733f
C19327 _439_.ZN a_39760_23588# 0.00245f
C19328 a_1828_28292# a_1468_28248# 0.08717f
C19329 a_3620_28292# a_4068_28292# 0.01328f
C19330 a_2276_22020# a_2364_21976# 0.28563f
C19331 _251_.A1 _267_.A2 0.25097f
C19332 a_49404_2727# a_49764_2824# 0.08717f
C19333 a_65668_17316# a_65756_17272# 0.28563f
C19334 _474_.Q _427_.B2 0.10644f
C19335 _437_.A1 a_37532_21543# 0.00222f
C19336 a_4068_16936# a_4068_15748# 0.05841f
C19337 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN a_56596_18504# 0.07124f
C19338 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN a_56932_23208# 0.00274f
C19339 a_45732_18504# a_46180_18504# 0.01328f
C19340 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN _245_.I1 0.0051f
C19341 a_17396_25156# a_17844_25156# 0.01328f
C19342 _284_.ZN _470_.D 0.06256f
C19343 _290_.ZN _362_.ZN 0.0068f
C19344 _324_.C a_44948_28292# 0.00755f
C19345 a_28908_20408# a_29356_20408# 0.0131f
C19346 a_45820_13703# a_45732_13800# 0.28563f
C19347 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_63764_23588# 0.04735f
C19348 a_32604_16839# a_32516_16936# 0.28563f
C19349 a_22100_31048# a_20672_30301# 0.00563f
C19350 input9.Z a_56260_31048# 0.06284f
C19351 a_27588_1636# VPWR 0.20909f
C19352 a_52292_29480# VPWR 0.00665f
C19353 a_63292_12568# a_63740_12568# 0.01288f
C19354 a_67236_12612# a_66876_12568# 0.08707f
C19355 a_5052_23544# a_4940_23111# 0.02634f
C19356 a_53684_12232# a_53772_10567# 0.00151f
C19357 _441_.A3 a_39796_22504# 0.00135f
C19358 a_44612_1636# a_44252_1592# 0.08707f
C19359 _362_.B a_35140_26680# 0.25577f
C19360 _279_.Z a_49316_23588# 0.01237f
C19361 _355_.C a_24900_27912# 0.00401f
C19362 a_61836_26680# a_61948_26247# 0.02634f
C19363 a_38576_22504# _301_.Z 0.45654f
C19364 a_60492_28248# a_60604_27815# 0.02634f
C19365 a_59172_23588# VPWR 0.12519f
C19366 a_14708_26724# a_14796_26680# 0.28563f
C19367 hold2.I a_44786_24120# 0.49079f
C19368 _258_.I _324_.C 0.02839f
C19369 _272_.A2 _255_.I 0.00332f
C19370 a_40892_1159# a_41340_1159# 0.0131f
C19371 _327_.A2 _325_.A2 0.92582f
C19372 _264_.B VPWR 0.52966f
C19373 a_53996_24679# a_53908_24776# 0.28563f
C19374 a_17844_20452# VPWR 0.21258f
C19375 a_15604_27912# a_15692_26247# 0.0027f
C19376 _349_.A4 a_26148_28776# 0.00236f
C19377 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I 0.10089f
C19378 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN 0.02352f
C19379 a_53124_12612# VPWR 0.2267f
C19380 a_65332_16936# a_66004_16936# 0.00347f
C19381 a_6172_30951# uio_oe[7] 0.00469f
C19382 _355_.C _358_.A3 0.00257f
C19383 a_8636_29383# a_8548_29480# 0.28563f
C19384 a_44836_15368# a_45284_15368# 0.01328f
C19385 _444_.D a_35616_24776# 0.26623f
C19386 a_5052_28248# a_4940_27815# 0.02634f
C19387 _424_.B1 a_50464_24908# 0.00157f
C19388 a_45732_10664# VPWR 0.20348f
C19389 a_67100_2727# a_67236_1636# 0.00154f
C19390 a_46940_15271# a_46852_15368# 0.28563f
C19391 _474_.CLK a_54780_18840# 0.00775f
C19392 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I rst_n 0.01432f
C19393 _351_.A2 a_25008_25597# 0.00268f
C19394 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I 0.01135f
C19395 a_48284_15271# a_48732_15271# 0.0131f
C19396 a_61276_15271# VPWR 0.32052f
C19397 _337_.ZN _358_.A2 0.01885f
C19398 _332_.Z VPWR 0.61456f
C19399 _434_.ZN _301_.A1 0.55565f
C19400 _384_.ZN _393_.A3 0.02146f
C19401 _386_.ZN _470_.Q 0.31556f
C19402 a_19636_22020# a_20084_22020# 0.01328f
C19403 a_16052_22020# a_16140_21976# 0.28563f
C19404 a_64860_15704# VPWR 0.3337f
C19405 a_60828_2727# a_60740_2824# 0.28563f
C19406 a_4940_16839# a_5388_16839# 0.01222f
C19407 a_45148_30951# a_45060_31048# 0.28563f
C19408 a_37780_16936# a_37892_15748# 0.02666f
C19409 a_38816_27555# _438_.A2 0.00109f
C19410 a_52415_31220# _274_.ZN 0.00374f
C19411 a_26468_23208# a_26556_21543# 0.00151f
C19412 a_26220_23544# a_26668_23544# 0.01255f
C19413 a_15492_1256# VPWR 0.20968f
C19414 a_5052_7864# VPWR 0.33516f
C19415 _244_.Z vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN 0.00217f
C19416 a_41700_1256# a_42148_1256# 0.01328f
C19417 a_65668_4772# VPWR 0.21209f
C19418 _303_.ZN _450_.D 0.01958f
C19419 a_56460_13703# a_57044_13800# 0.01675f
C19420 a_53660_14136# a_53572_12612# 0.00151f
C19421 a_2724_13800# a_3172_13800# 0.01328f
C19422 a_6172_29383# VPWR 0.3289f
C19423 a_20956_2727# a_21404_2727# 0.0131f
C19424 a_61524_20452# a_61612_20408# 0.28563f
C19425 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN 0.00469f
C19426 _245_.I1 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN 0.06924f
C19427 a_4156_17272# a_4156_16839# 0.05841f
C19428 _330_.A1 a_41099_26841# 0.01174f
C19429 a_43468_16839# a_43828_16936# 0.08707f
C19430 a_58924_10567# a_58948_9476# 0.0016f
C19431 a_33724_1592# VPWR 0.30128f
C19432 a_2364_1159# a_2276_1256# 0.28563f
C19433 a_31172_16936# VPWR 0.20348f
C19434 a_4604_12568# a_4516_11044# 0.0027f
C19435 a_21068_23544# a_20956_23111# 0.02634f
C19436 a_7652_1636# a_7292_1592# 0.08707f
C19437 a_44388_27912# VPWR 0.20529f
C19438 a_2276_29860# a_2364_29816# 0.28563f
C19439 a_5860_29860# a_6308_29860# 0.01328f
C19440 a_3260_17272# a_3708_17272# 0.0131f
C19441 a_51108_1636# a_51556_1636# 0.01328f
C19442 a_36772_23208# _301_.A1 0.00856f
C19443 a_57692_11000# a_58140_11000# 0.01288f
C19444 a_36500_29860# uo_out[2] 0.00289f
C19445 a_47164_18407# a_47076_18504# 0.28563f
C19446 _395_.A2 _427_.B2 0.00354f
C19447 a_48868_18504# a_48844_16839# 0.00131f
C19448 a_19412_27912# a_18096_27165# 0.03574f
C19449 a_65668_18884# a_65308_18840# 0.0869f
C19450 a_66092_18407# VPWR 0.35599f
C19451 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I 0.02602f
C19452 _421_.A1 _417_.A2 0.08966f
C19453 a_4604_25112# VPWR 0.33016f
C19454 a_28820_20452# VPWR 0.20622f
C19455 _324_.C hold1.Z 0.0198f
C19456 _476_.Q a_54244_20452# 0.00148f
C19457 a_66788_12612# VPWR 0.20622f
C19458 a_23644_29816# VPWR 0.34964f
C19459 _447_.Q a_38676_20452# 0.00178f
C19460 a_65756_26247# clk 0.00118f
C19461 _352_.A2 a_30520_27508# 0.00649f
C19462 a_21764_2824# a_22212_2824# 0.01328f
C19463 _230_.I a_60852_28292# 0.00192f
C19464 _381_.Z clkbuf_1_0__f_clk.I 0.00637f
C19465 a_67117_30600# vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN 0.02548f
C19466 _246_.B2 a_60156_27815# 0.05374f
C19467 _378_.ZN a_17844_27912# 0.00275f
C19468 a_55252_24776# a_55700_24776# 0.01328f
C19469 a_67572_10664# VPWR 0.20703f
C19470 a_66652_8999# a_66564_9096# 0.28563f
C19471 a_67548_7431# a_67460_7528# 0.28563f
C19472 a_16052_21640# a_16052_20452# 0.05841f
C19473 a_39300_29480# VPWR 0.01802f
C19474 a_61748_16936# VPWR 0.20944f
C19475 _462_.D uo_out[2] 0.00867f
C19476 a_41028_15368# VPWR 0.2059f
C19477 vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN VPWR 0.73508f
C19478 a_43003_28409# a_43288_28409# 0.00277f
C19479 a_19035_28409# uio_out[7] 0.01249f
C19480 a_3260_14136# a_3708_14136# 0.0131f
C19481 _324_.C a_45396_25156# 0.00132f
C19482 a_44476_15271# VPWR 0.29679f
C19483 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I 0.00401f
C19484 a_29804_23544# a_29716_22020# 0.00151f
C19485 a_48560_26369# VPWR 0.00326f
C19486 a_44724_16936# a_44836_15748# 0.02666f
C19487 a_40916_16936# a_40892_15704# 0.0016f
C19488 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I 0.12732f
C19489 a_1020_16839# VPWR 0.30073f
C19490 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN VPWR 0.84918f
C19491 a_37892_1256# VPWR 0.20348f
C19492 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN a_56236_24679# 0.0012f
C19493 a_66204_3160# a_66204_2727# 0.05841f
C19494 a_67660_13703# a_67572_13800# 0.28563f
C19495 _346_.B a_21287_29076# 0.01021f
C19496 _226_.ZN a_41696_24072# 0.00265f
C19497 a_43750_23544# _305_.A2 0.00924f
C19498 a_4068_17316# VPWR 0.2157f
C19499 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN a_67684_24776# 0.00152f
C19500 a_54444_16839# a_54356_16936# 0.28563f
C19501 _355_.C a_28256_25597# 0.00856f
C19502 a_3708_12135# a_4068_12232# 0.08717f
C19503 a_47388_1592# VPWR 0.35728f
C19504 a_48956_12568# a_48868_11044# 0.0027f
C19505 a_13340_1159# a_13700_1256# 0.08717f
C19506 a_53012_16936# VPWR 0.2061f
C19507 a_57580_12135# a_58028_12135# 0.01288f
C19508 a_10564_1636# a_10652_1592# 0.28563f
C19509 a_14148_1636# a_14596_1636# 0.01328f
C19510 a_6532_29480# a_6980_29480# 0.01328f
C19511 vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I VPWR 0.7144f
C19512 _416_.A1 hold2.Z 0.04129f
C19513 a_35652_17316# a_35292_17272# 0.08707f
C19514 a_64996_11044# a_65084_11000# 0.28563f
C19515 a_30160_30301# uo_out[7] 0.00603f
C19516 a_43716_31048# a_44164_31048# 0.01328f
C19517 a_17956_2824# VPWR 0.2067f
C19518 _459_.CLK a_14796_26680# 0.00135f
C19519 a_63092_26724# a_62732_26680# 0.0869f
C19520 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I a_63428_20072# 0.00242f
C19521 _416_.A1 _416_.A3 0.73052f
C19522 _455_.Q a_20756_26724# 0.00519f
C19523 a_44786_24120# VPWR 0.74023f
C19524 a_2364_24679# a_2276_24776# 0.28563f
C19525 a_20060_24679# a_20508_24679# 0.01288f
C19526 _459_.CLK a_24316_26247# 0.0101f
C19527 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I clk 0.0724f
C19528 _360_.ZN a_33188_25940# 0.60215f
C19529 a_40038_28720# a_40780_27815# 0.00198f
C19530 a_63292_1159# a_63740_1159# 0.0131f
C19531 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_65756_26247# 0.02235f
C19532 a_2812_19975# a_3260_19975# 0.0131f
C19533 a_47972_2824# a_47972_1636# 0.05841f
C19534 a_4068_14180# VPWR 0.2157f
C19535 _474_.CLK a_55700_23588# 0.05032f
C19536 a_1380_4392# a_1828_4392# 0.01328f
C19537 a_4156_18407# a_4940_18407# 0.00443f
C19538 _432_.ZN _304_.A1 0.0324f
C19539 _230_.I _238_.I 0.49567f
C19540 a_61188_20072# vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN 0.00147f
C19541 _260_.A1 a_42982_21730# 0.0057f
C19542 a_2724_29480# VPWR 0.20782f
C19543 a_32604_15704# a_33052_15704# 0.01288f
C19544 a_53772_12135# VPWR 0.31547f
C19545 a_36548_15748# a_36636_15704# 0.28563f
C19546 a_45820_15704# a_45956_15368# 0.00168f
C19547 _438_.A2 _447_.Q 0.24976f
C19548 _397_.A4 _419_.A4 0.3738f
C19549 _334_.A1 _460_.Q 0.23234f
C19550 _474_.CLK vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN 0.13001f
C19551 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I a_58476_20408# 0.01277f
C19552 a_16140_24679# VPWR 0.29679f
C19553 _452_.CLK a_46716_18407# 0.00144f
C19554 a_43296_28733# a_43003_28409# 0.49319f
C19555 a_38852_25156# VPWR 0.00672f
C19556 a_36548_15748# VPWR 0.20622f
C19557 a_47552_19715# a_48084_18884# 0.03552f
C19558 a_48060_18407# a_48508_18407# 0.0131f
C19559 a_2724_9476# a_2812_9432# 0.28563f
C19560 _470_.Q a_47476_28292# 0.01423f
C19561 _228_.ZN _255_.I 0.00604f
C19562 _255_.ZN _324_.C 0.06142f
C19563 a_29716_22020# a_29804_21976# 0.28563f
C19564 a_25772_21976# a_26220_21976# 0.01288f
C19565 a_51756_16839# a_52204_16839# 0.0131f
C19566 a_50212_14180# a_49852_14136# 0.08707f
C19567 _229_.I a_60828_26680# 0.00111f
C19568 a_43452_18191# VPWR 0.39888f
C19569 _300_.ZN a_39780_22805# 0.00955f
C19570 _452_.CLK a_44724_17316# 0.0065f
C19571 a_47948_16839# VPWR 0.31556f
C19572 a_51668_16936# a_51780_15748# 0.02666f
C19573 a_47860_16936# a_47836_15704# 0.0016f
C19574 a_60292_1256# VPWR 0.20348f
C19575 a_26556_30951# uio_out[1] 0.00808f
C19576 a_64100_1256# a_64548_1256# 0.01328f
C19577 a_64212_13800# a_64884_13800# 0.00347f
C19578 _460_.Q a_35156_29860# 0.00226f
C19579 a_43828_29860# a_44632_30206# 0.00304f
C19580 a_43356_2727# a_43804_2727# 0.0131f
C19581 a_36016_20893# VPWR 0.51676f
C19582 _379_.A2 VPWR 1.51592f
C19583 _435_.A3 _441_.B 0.02009f
C19584 a_40132_20452# a_40580_20452# 0.01328f
C19585 a_39236_17316# VPWR 0.20765f
C19586 a_24764_1159# a_24676_1256# 0.28563f
C19587 a_54668_12135# a_54580_12232# 0.28563f
C19588 a_61188_1636# VPWR 0.20348f
C19589 _355_.ZN a_27924_24776# 0.03932f
C19590 _325_.A1 a_43824_18147# 0.01254f
C19591 a_55724_22137# VPWR 0.00246f
C19592 a_11996_29816# a_12444_29816# 0.01288f
C19593 a_15940_29860# a_16028_29816# 0.28563f
C19594 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I a_64660_23588# 0.00409f
C19595 a_2276_26344# a_2276_25156# 0.05841f
C19596 a_51332_24372# clk 0.01535f
C19597 _427_.B1 a_52920_22760# 0.02976f
C19598 _336_.A2 a_28460_23544# 0.00513f
C19599 a_40356_2824# VPWR 0.20815f
C19600 _386_.A4 _470_.Q 0.06918f
C19601 a_37668_1636# a_37532_1159# 0.00168f
C19602 a_33724_1592# a_33724_1159# 0.05841f
C19603 a_57244_1592# a_57692_1592# 0.01288f
C19604 a_61188_1636# a_61276_1592# 0.28563f
C19605 a_4940_10567# a_5388_10567# 0.01222f
C19606 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN 0.00681f
C19607 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN 0.01282f
C19608 a_30588_23111# a_31036_23111# 0.01288f
C19609 a_18716_23111# a_19076_23208# 0.08707f
C19610 a_22300_24679# a_22660_24776# 0.08707f
C19611 _330_.A1 a_35816_21192# 0.0247f
C19612 _390_.ZN a_52676_27912# 0.00429f
C19613 a_47076_9476# VPWR 0.20348f
C19614 a_53124_14180# VPWR 0.22915f
C19615 a_3708_21543# a_4156_21543# 0.0131f
C19616 a_35652_31048# _460_.Q 0.01316f
C19617 _388_.B a_45800_30345# 0.00582f
C19618 a_35180_18407# a_35092_18504# 0.28563f
C19619 a_7540_31048# a_7652_29860# 0.02666f
C19620 a_36300_23544# _437_.ZN 0.00217f
C19621 _248_.B1 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I 0.13872f
C19622 a_47524_12232# VPWR 0.20348f
C19623 a_39908_15748# a_39548_15704# 0.08707f
C19624 _398_.C a_51576_25896# 0.03579f
C19625 a_44164_2824# a_44612_2824# 0.01328f
C19626 a_52764_15704# a_52900_15368# 0.00168f
C19627 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN a_55252_25156# 0.00105f
C19628 _392_.A2 a_49652_29480# 0.03524f
C19629 _427_.A2 _427_.B2 0.02189f
C19630 a_2364_20408# a_2364_19975# 0.05841f
C19631 a_20868_24776# VPWR 0.20595f
C19632 a_54692_15748# a_54556_15271# 0.00168f
C19633 _427_.B2 a_51196_21543# 0.00449f
C19634 a_4828_2727# a_4740_2824# 0.28563f
C19635 _250_.ZN a_60404_28292# 0.00118f
C19636 _246_.B2 a_60516_27912# 0.02029f
C19637 a_31260_19975# a_31620_20072# 0.08717f
C19638 a_42684_15704# VPWR 0.3429f
C19639 a_61948_26247# a_62396_26247# 0.012f
C19640 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I 0.00995f
C19641 _359_.B _393_.ZN 0.00914f
C19642 a_47164_9432# a_47612_9432# 0.0131f
C19643 vgaringosc.workerclkbuff_notouch_.I a_49600_30180# 0.01788f
C19644 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN VPWR 0.88816f
C19645 a_14684_29383# a_14708_28292# 0.0016f
C19646 a_63964_19975# VPWR 0.33016f
C19647 _300_.ZN a_39796_22504# 0.00863f
C19648 _325_.A1 _302_.Z 0.06359f
C19649 a_53572_14180# a_53660_14136# 0.28563f
C19650 a_56708_14180# a_57156_14180# 0.01328f
C19651 _304_.B _395_.A3 0.03911f
C19652 _452_.CLK a_37980_26247# 0.00722f
C19653 a_19724_25112# a_19636_23588# 0.00151f
C19654 _294_.A2 _337_.ZN 0.01765f
C19655 _452_.CLK a_33276_21543# 0.02574f
C19656 _416_.A1 a_45036_28248# 0.02833f
C19657 a_53212_17272# a_53100_16839# 0.02634f
C19658 _474_.CLK a_53460_24776# 0.00252f
C19659 _412_.A1 a_51968_26724# 0.00636f
C19660 _251_.A1 _256_.A2 0.03016f
C19661 a_35740_26247# VPWR 0.31306f
C19662 a_50524_17272# VPWR 0.35503f
C19663 _260_.A1 _304_.A1 0.5752f
C19664 a_3260_1159# VPWR 0.30487f
C19665 a_35740_1159# a_36100_1256# 0.08717f
C19666 _327_.A2 a_43824_18147# 0.00128f
C19667 a_49292_12135# a_49316_11044# 0.0016f
C19668 a_20284_1592# a_20732_1592# 0.01288f
C19669 a_65420_12135# a_65780_12232# 0.08717f
C19670 a_51444_12232# a_51892_12232# 0.01328f
C19671 a_31036_21543# VPWR 0.31547f
C19672 a_61836_25515# vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN 0.00606f
C19673 _279_.Z _399_.ZN 0.18882f
C19674 a_39480_28776# uo_out[7] 0.0016f
C19675 a_47748_17316# a_47388_17272# 0.08707f
C19676 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN VPWR 0.78488f
C19677 a_43850_23588# VPWR 0.00401f
C19678 _478_.D a_54192_22851# 0.24091f
C19679 a_1916_10567# a_1828_10664# 0.28563f
C19680 a_62756_2824# VPWR 0.20815f
C19681 a_65892_1636# a_65980_1592# 0.28563f
C19682 _438_.A2 a_40004_23233# 0.0052f
C19683 _395_.A1 a_50732_23233# 0.00158f
C19684 a_29692_23111# a_29604_23208# 0.28563f
C19685 a_24452_24776# a_24900_24776# 0.01328f
C19686 a_58052_9476# VPWR 0.2284f
C19687 a_2364_21543# a_2724_21640# 0.08717f
C19688 a_1380_3204# VPWR 0.20348f
C19689 a_61500_14136# VPWR 0.31389f
C19690 a_60276_29032# _250_.C 0.00355f
C19691 _324_.C a_46198_27060# 0.02825f
C19692 _476_.Q a_52081_21236# 0.00603f
C19693 _230_.I vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN 0.03048f
C19694 a_46404_15748# a_46852_15748# 0.01328f
C19695 a_9668_29860# a_9532_29383# 0.00168f
C19696 a_1828_11044# VPWR 0.20348f
C19697 a_47776_20893# VPWR 0.51898f
C19698 a_51332_24072# a_51988_24072# 0.01436f
C19699 a_62620_19975# a_62532_20072# 0.28563f
C19700 a_20672_30301# uio_out[6] 0.04269f
C19701 a_65308_18840# a_65308_18407# 0.05841f
C19702 _324_.C clkbuf_1_0__f_clk.I 0.15418f
C19703 a_2812_18840# VPWR 0.30213f
C19704 _424_.A2 a_45696_20072# 0.00533f
C19705 a_15580_2727# a_16164_2824# 0.01675f
C19706 _324_.B a_43380_20452# 0.0028f
C19707 _416_.A1 a_49652_29480# 0.00567f
C19708 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I clk 0.0136f
C19709 _264_.B _260_.ZN 0.03319f
C19710 _363_.Z a_32848_29123# 0.0418f
C19711 _417_.A2 a_49034_21640# 0.01021f
C19712 a_52900_9476# a_52988_9432# 0.28563f
C19713 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN 0.0619f
C19714 _302_.Z _327_.A2 0.00642f
C19715 a_51791_30644# input9.Z 0.0014f
C19716 _397_.A4 a_51048_26680# 0.00114f
C19717 a_64660_23588# VPWR 0.21229f
C19718 a_1468_20408# a_1916_20408# 0.0131f
C19719 a_4068_20452# a_3708_20408# 0.08717f
C19720 a_50524_17272# a_50436_15748# 0.00151f
C19721 _395_.A3 VPWR 0.7916f
C19722 hold2.I a_41564_24679# 0.00637f
C19723 a_49764_12612# a_49852_12568# 0.28563f
C19724 _223_.I a_31920_29480# 0.0032f
C19725 a_45820_12568# a_46268_12568# 0.01288f
C19726 a_65756_2727# a_66204_2727# 0.01255f
C19727 _478_.D _281_.A1 0.06713f
C19728 a_47164_1159# a_47076_1256# 0.28563f
C19729 _459_.Q a_34586_27912# 0.00126f
C19730 a_25660_1159# VPWR 0.33232f
C19731 a_4852_5960# a_4940_4295# 0.00151f
C19732 a_65980_12568# a_65892_11044# 0.00151f
C19733 a_46180_12232# a_46180_11044# 0.05841f
C19734 a_65756_27815# a_65668_27912# 0.28563f
C19735 a_27588_1636# a_27228_1592# 0.08707f
C19736 _452_.Q a_40644_17272# 0.02136f
C19737 a_39324_26247# a_39772_26247# 0.01255f
C19738 a_35740_26247# a_36100_26344# 0.0869f
C19739 a_28260_21640# VPWR 0.20614f
C19740 _258_.I a_59796_29480# 0.01327f
C19741 a_52428_10567# a_52788_10664# 0.08707f
C19742 a_66316_10567# a_66764_10567# 0.0131f
C19743 a_7068_1159# a_7516_1159# 0.0131f
C19744 _290_.ZN a_35008_27533# 0.00629f
C19745 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN 0.07488f
C19746 _230_.I VPWR 2.3009f
C19747 a_28260_23208# a_28708_23208# 0.01328f
C19748 _304_.B a_44038_21236# 0.06258f
C19749 a_30240_24776# a_31120_24463# 0.00306f
C19750 a_1916_8999# VPWR 0.297f
C19751 a_17932_23544# VPWR 0.30035f
C19752 a_22748_21543# a_22660_21640# 0.28563f
C19753 a_3708_5863# VPWR 0.33374f
C19754 _416_.A1 _448_.Q 0.00223f
C19755 a_932_21640# a_1380_21640# 0.01328f
C19756 a_5724_2727# VPWR 0.33105f
C19757 a_55564_13703# VPWR 0.31594f
C19758 a_36996_2824# a_37084_1159# 0.0027f
C19759 a_59172_27912# a_60068_27912# 0.00455f
C19760 a_53572_15748# a_53212_15704# 0.08663f
C19761 a_50748_11000# VPWR 0.32523f
C19762 a_66564_2824# a_67012_2824# 0.01328f
C19763 a_1916_21976# a_1916_21543# 0.05841f
C19764 _350_.A1 a_29716_31048# 0.01868f
C19765 a_1916_26680# VPWR 0.297f
C19766 a_63876_15748# a_64324_15748# 0.01328f
C19767 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I 0.01236f
C19768 _416_.A3 a_47300_17316# 0.0014f
C19769 a_32268_20408# a_32156_19975# 0.02634f
C19770 a_50436_30689# vgaringosc.workerclkbuff_notouch_.I 0.00597f
C19771 a_18628_26344# VPWR 0.23332f
C19772 a_26160_27165# a_27228_26680# 0.00506f
C19773 a_27004_2727# a_26916_2824# 0.28563f
C19774 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN 0.00202f
C19775 a_61076_20452# VPWR 0.15188f
C19776 a_25100_30951# uio_out[3] 0.00333f
C19777 _304_.B a_51084_28248# 0.00664f
C19778 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I clk 0.00118f
C19779 _474_.CLK clkload0.Z 0.00123f
C19780 _474_.CLK a_52316_17272# 0.00111f
C19781 a_58140_9432# a_58588_9432# 0.0131f
C19782 a_59844_9476# a_60516_9476# 0.00347f
C19783 a_61948_26247# a_61860_26344# 0.28563f
C19784 _393_.ZN _386_.ZN 0.00193f
C19785 a_15156_28292# VPWR 0.20703f
C19786 a_1380_23588# a_1020_23544# 0.08717f
C19787 a_3172_23588# a_3620_23588# 0.01328f
C19788 a_2276_7908# a_2724_7908# 0.01328f
C19789 a_7876_1256# a_8548_1256# 0.00347f
C19790 a_31820_21976# a_31732_20452# 0.00151f
C19791 a_3172_6340# a_3620_6340# 0.01328f
C19792 a_2276_4772# a_1916_4728# 0.08717f
C19793 a_4068_4772# a_4516_4772# 0.01328f
C19794 a_1380_6340# a_1020_6296# 0.08717f
C19795 a_65084_14136# a_65532_14136# 0.01288f
C19796 a_3172_3204# a_2812_3160# 0.08717f
C19797 _304_.B a_41564_24679# 0.02422f
C19798 a_56596_23588# a_56684_23544# 0.28563f
C19799 a_61860_30736# _229_.I 0.00233f
C19800 _294_.A2 a_30795_29977# 0.06222f
C19801 a_52540_12568# a_53212_12568# 0.00544f
C19802 a_55476_13800# a_55564_12135# 0.00151f
C19803 a_7204_1636# VPWR 0.2085f
C19804 _459_.CLK a_17844_25156# 0.00249f
C19805 _451_.Q a_38676_20452# 0.00143f
C19806 a_59260_21976# vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I 0.00103f
C19807 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I a_58500_21640# 0.00569f
C19808 _398_.C a_53460_24776# 0.0077f
C19809 _397_.A4 _381_.A2 0.03009f
C19810 a_47525_29480# VPWR 0.52191f
C19811 a_7740_29816# a_7876_29480# 0.00168f
C19812 a_48060_1159# VPWR 0.29679f
C19813 a_37516_27599# uo_out[7] 0.00182f
C19814 _371_.A2 a_28036_26724# 0.00291f
C19815 a_58140_1159# a_58500_1256# 0.08717f
C19816 a_65668_18884# VPWR 0.21801f
C19817 a_34084_1636# a_34532_1636# 0.01328f
C19818 a_1020_11000# a_1468_11000# 0.0131f
C19819 a_3620_11044# a_3260_11000# 0.08717f
C19820 _304_.B _325_.A2 0.03409f
C19821 a_53236_12232# a_53124_11044# 0.02666f
C19822 _459_.Q a_30160_30301# 0.01142f
C19823 _424_.B1 _476_.Q 0.33259f
C19824 a_66092_16839# a_66540_16839# 0.01255f
C19825 a_47483_20569# a_47768_20569# 0.00277f
C19826 a_50212_20452# a_50300_20408# 0.28563f
C19827 a_44028_27815# a_44476_27815# 0.01222f
C19828 _373_.ZN a_28432_29535# 0.00144f
C19829 a_63404_10567# a_63316_10664# 0.28563f
C19830 _275_.A2 a_51050_29480# 0.01277f
C19831 _459_.CLK _352_.A2 0.23604f
C19832 _284_.ZN _459_.CLK 0.51624f
C19833 _337_.A3 _337_.ZN 1.25822f
C19834 a_18828_21976# VPWR 0.3241f
C19835 a_60852_15748# a_60940_15704# 0.28563f
C19836 _260_.A2 _304_.A1 0.02302f
C19837 a_44038_21236# VPWR 0.31199f
C19838 a_33276_21543# a_33636_21640# 0.08663f
C19839 a_31620_18884# a_32068_18884# 0.01328f
C19840 a_30476_23544# VPWR 0.3185f
C19841 a_49652_13800# VPWR 0.21158f
C19842 a_28124_2727# VPWR 0.31143f
C19843 a_1468_26247# a_1916_26247# 0.0131f
C19844 _279_.Z a_48516_24080# 0.00161f
C19845 a_44906_23588# VPWR 0.0043f
C19846 a_5052_29816# VPWR 0.3289f
C19847 a_64548_11044# VPWR 0.21169f
C19848 a_17932_21976# a_17932_21543# 0.05841f
C19849 a_52764_2727# a_52900_1636# 0.00154f
C19850 a_21876_22020# a_21852_21543# 0.00172f
C19851 _304_.B a_53124_27912# 0.02325f
C19852 a_15692_23111# VPWR 0.29679f
C19853 _304_.A1 a_36084_23208# 0.00315f
C19854 a_16052_27912# VPWR 0.20348f
C19855 a_25124_28776# a_26148_28776# 0.00825f
C19856 a_65756_23111# a_65668_23208# 0.28563f
C19857 a_37980_2727# a_38340_2824# 0.08717f
C19858 a_51084_28248# VPWR 0.32968f
C19859 _355_.C a_25232_27165# 0.00818f
C19860 a_30724_26020# a_29828_26344# 0.00172f
C19861 a_15156_23588# a_14796_23544# 0.08707f
C19862 a_2364_7864# a_2364_7431# 0.05841f
C19863 a_1828_25156# a_2276_25156# 0.01328f
C19864 a_65668_7908# a_65308_7864# 0.08717f
C19865 a_4156_4728# a_4156_4295# 0.05841f
C19866 a_67460_4772# a_67100_4728# 0.08717f
C19867 a_54804_20072# vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I 0.00131f
C19868 a_3260_6296# a_3260_5863# 0.05841f
C19869 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN 0.65285f
C19870 a_66564_6340# a_66204_6296# 0.08717f
C19871 a_63428_20072# a_63428_18884# 0.05841f
C19872 a_62564_29032# _250_.C 0.02826f
C19873 _250_.ZN _248_.B1 0.00375f
C19874 a_62396_14136# a_62508_13703# 0.02634f
C19875 a_17732_31048# _379_.Z 0.00198f
C19876 a_25012_20452# a_25460_20452# 0.01328f
C19877 a_23668_20452# a_23308_20408# 0.08717f
C19878 _459_.Q a_33520_25597# 0.00286f
C19879 a_41564_24679# VPWR 0.3494f
C19880 a_13004_30951# a_12916_31048# 0.28563f
C19881 _427_.ZN vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.00817f
C19882 a_67908_17316# a_67884_16839# 0.00172f
C19883 a_4940_10567# a_4964_9476# 0.0016f
C19884 a_13340_1592# VPWR 0.29679f
C19885 a_59484_12568# a_59932_12568# 0.01288f
C19886 _424_.B1 a_50084_24328# 0.01433f
C19887 _397_.A2 _279_.Z 0.12443f
C19888 a_46268_12568# a_46268_12135# 0.05841f
C19889 a_50212_12612# a_50188_12135# 0.00172f
C19890 a_47972_31048# vgaringosc.workerclkbuff_notouch_.I 0.0065f
C19891 _255_.I ui_in[3] 0.00206f
C19892 _359_.B a_33483_29535# 0.01597f
C19893 _438_.A2 _451_.Q 0.02764f
C19894 a_30796_24463# a_31284_23588# 0.01025f
C19895 a_64324_9096# VPWR 0.22383f
C19896 _325_.A2 VPWR 1.47367f
C19897 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN _250_.ZN 0.0051f
C19898 a_66116_5960# VPWR 0.23643f
C19899 a_64212_23588# a_63852_23544# 0.0869f
C19900 a_17140_26841# VPWR 0.00246f
C19901 a_47972_11044# a_47612_11000# 0.08707f
C19902 _437_.A1 a_37444_25156# 0.00551f
C19903 a_36524_18407# VPWR 0.30655f
C19904 a_54432_31128# _274_.A2 0.00821f
C19905 a_34084_28776# a_35516_28776# 0.01047f
C19906 _459_.CLK a_20508_24679# 0.00239f
C19907 a_54780_20408# a_54804_20072# 0.00172f
C19908 _325_.A2 a_44364_17272# 0.01303f
C19909 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.00267f
C19910 a_65892_1636# a_65756_1159# 0.00168f
C19911 a_29468_1159# a_29916_1159# 0.0131f
C19912 a_60180_10664# a_60628_10664# 0.01328f
C19913 a_27588_26344# _355_.ZN 0.00964f
C19914 a_22212_24776# a_22300_23111# 0.0027f
C19915 a_3708_26680# a_3708_26247# 0.05841f
C19916 a_30476_21976# VPWR 0.3185f
C19917 _303_.ZN a_38576_22504# 0.00767f
C19918 a_56404_27208# a_56516_26344# 0.0146f
C19919 _287_.A1 a_32132_27912# 0.00873f
C19920 a_31844_21640# a_32292_21640# 0.01328f
C19921 _421_.A1 a_45920_20523# 0.00898f
C19922 vgaringosc.workerclkbuff_notouch_.I VPWR 1.41471f
C19923 a_50524_2727# VPWR 0.35938f
C19924 a_3620_12612# VPWR 0.22347f
C19925 a_16588_26247# a_16500_26344# 0.28563f
C19926 _436_.B a_40468_25157# 0.02346f
C19927 a_33412_15368# a_33860_15368# 0.01328f
C19928 a_26468_27912# a_26160_27165# 0.0022f
C19929 _435_.A3 _452_.Q 0.01666f
C19930 a_17148_29816# VPWR 0.29679f
C19931 _475_.Q a_50300_20408# 0.0069f
C19932 _301_.A1 a_36148_21976# 0.22573f
C19933 _352_.A2 _371_.A3 0.43866f
C19934 a_51532_10567# VPWR 0.31389f
C19935 a_35516_15271# a_35428_15368# 0.28563f
C19936 a_28820_22020# a_28796_21543# 0.00172f
C19937 a_24876_21976# a_24988_21543# 0.02634f
C19938 a_4068_23208# VPWR 0.22146f
C19939 a_53124_27912# VPWR 0.20818f
C19940 a_36860_15271# a_37308_15271# 0.0131f
C19941 _304_.B _427_.B1 0.99631f
C19942 _439_.ZN a_39536_23588# 0.00446f
C19943 _371_.ZN _359_.B 0.46026f
C19944 _350_.A1 _365_.ZN 0.05489f
C19945 a_1380_28292# a_1468_28248# 0.28563f
C19946 a_2276_22020# a_1916_21976# 0.08717f
C19947 a_4068_22020# a_4516_22020# 0.01328f
C19948 a_49404_2727# a_49316_2824# 0.28563f
C19949 a_65668_17316# a_65308_17272# 0.0869f
C19950 _346_.A2 a_22548_25156# 0.00203f
C19951 a_57020_23111# a_56932_23208# 0.28563f
C19952 a_63092_26724# _245_.I1 0.00147f
C19953 a_65308_7431# a_65756_7431# 0.0131f
C19954 a_21516_23544# a_21964_23544# 0.012f
C19955 a_64412_8999# a_64860_8999# 0.0131f
C19956 a_30276_1256# a_30724_1256# 0.01328f
C19957 a_66204_5863# a_66652_5863# 0.0131f
C19958 a_67100_4295# a_67548_4295# 0.0131f
C19959 a_49852_14136# a_49764_12612# 0.00151f
C19960 a_45372_13703# a_45732_13800# 0.08717f
C19961 a_59372_13703# a_59820_13703# 0.01288f
C19962 a_9532_2727# a_9980_2727# 0.0131f
C19963 _268_.A2 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.09146f
C19964 a_41364_16936# a_41564_15271# 0.00119f
C19965 a_61412_26344# a_61860_26344# 0.01328f
C19966 a_66900_18504# a_67012_17316# 0.02666f
C19967 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_63316_23588# 0.03728f
C19968 a_32156_16839# a_32516_16936# 0.08717f
C19969 a_1828_10664# a_1828_9476# 0.05841f
C19970 a_21652_31048# a_20672_30301# 0.03278f
C19971 a_52068_29480# VPWR 0.01379f
C19972 a_59828_26724# _251_.ZN 0.0019f
C19973 a_27140_1636# VPWR 0.25368f
C19974 a_13452_30951# a_14004_31048# 0.01375f
C19975 a_57156_12612# a_57132_12135# 0.00172f
C19976 a_53212_12568# a_53324_12135# 0.02634f
C19977 a_66788_12612# a_66876_12568# 0.28563f
C19978 _424_.A2 _428_.Z 0.49748f
C19979 _388_.B a_45088_29123# 0.0109f
C19980 a_63876_18504# a_64324_18504# 0.01328f
C19981 a_64860_26247# a_64772_26344# 0.28563f
C19982 a_54468_11044# a_54916_11044# 0.01328f
C19983 _284_.ZN uo_out[7] 0.05675f
C19984 a_2724_15368# a_2724_14180# 0.05841f
C19985 a_45620_16936# a_46068_16936# 0.01328f
C19986 a_12444_1592# a_12444_1159# 0.05841f
C19987 a_40220_1592# a_40668_1592# 0.01288f
C19988 a_44164_1636# a_44252_1592# 0.28563f
C19989 _279_.Z a_48308_23588# 0.8271f
C19990 a_58612_16936# vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN 0.00265f
C19991 _362_.B a_34532_27208# 0.01259f
C19992 a_14708_26724# a_15156_26724# 0.01328f
C19993 hold2.I a_44162_24120# 0.06762f
C19994 a_4940_27815# a_4964_26724# 0.0016f
C19995 _470_.Q a_47600_27912# 0.01065f
C19996 a_33636_2824# a_33636_1636# 0.05841f
C19997 _393_.ZN _386_.A4 0.01727f
C19998 a_53548_24679# a_53908_24776# 0.0869f
C19999 a_17396_20452# VPWR 0.20348f
C20000 a_57132_17272# vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN 0.00409f
C20001 _349_.A4 a_25740_28776# 0.00337f
C20002 _400_.ZN a_44571_26841# 0.00428f
C20003 a_52540_12568# VPWR 0.34385f
C20004 a_23420_26247# a_23868_26247# 0.01222f
C20005 _284_.ZN _480_.Q 0.0417f
C20006 a_10340_2824# a_10788_2824# 0.01328f
C20007 a_5724_30951# uio_oe[7] 0.00238f
C20008 a_7964_29383# a_8548_29480# 0.01675f
C20009 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I 0.05184f
C20010 a_45284_10664# VPWR 0.22176f
C20011 a_46492_15271# a_46852_15368# 0.08717f
C20012 a_23532_21976# a_23556_21640# 0.00172f
C20013 _459_.CLK _223_.ZN 0.02472f
C20014 _416_.ZN a_45732_18884# 0.00277f
C20015 _474_.CLK a_54332_18840# 0.01052f
C20016 a_64324_29860# rst_n 0.01008f
C20017 a_36996_26724# a_37444_26724# 0.01328f
C20018 a_34756_24776# a_34939_23705# 0.00123f
C20019 _427_.B1 VPWR 0.81743f
C20020 _337_.ZN a_29828_26344# 0.03191f
C20021 a_50084_24328# _218_.ZN 0.0018f
C20022 a_40244_18180# VPWR 0.77411f
C20023 a_60380_2727# a_60740_2824# 0.08717f
C20024 a_16052_22020# a_15692_21976# 0.08707f
C20025 a_23920_27555# VPWR 0.50741f
C20026 a_64412_15704# VPWR 0.29986f
C20027 a_44700_30951# a_45060_31048# 0.08717f
C20028 a_63876_15368# a_64324_15368# 0.01328f
C20029 a_15044_1256# VPWR 0.20348f
C20030 a_4604_7864# VPWR 0.33016f
C20031 _475_.Q _421_.B 0.00864f
C20032 _267_.A2 _255_.I 0.25795f
C20033 a_20172_25112# a_20620_25112# 0.01288f
C20034 a_65220_4772# VPWR 0.20921f
C20035 a_33948_18840# a_33948_18407# 0.05841f
C20036 a_5724_29383# VPWR 0.3289f
C20037 a_56460_13703# a_56372_13800# 0.28563f
C20038 a_52564_16936# a_52540_15271# 0.00134f
C20039 _350_.A1 a_29856_29123# 0.21345f
C20040 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I a_64412_29816# 0.04674f
C20041 a_61524_20452# a_61164_20408# 0.08674f
C20042 a_43468_16839# a_43380_16936# 0.28563f
C20043 _330_.A1 a_41392_27165# 0.02378f
C20044 _450_.D _452_.D 0.05282f
C20045 _250_.C _250_.B 0.47003f
C20046 a_33276_1592# VPWR 0.29975f
C20047 a_1916_1159# a_2276_1256# 0.08717f
C20048 a_46492_1592# a_46628_1256# 0.00168f
C20049 a_30724_16936# VPWR 0.22176f
C20050 a_3260_1592# a_3708_1592# 0.01288f
C20051 a_7204_1636# a_7292_1592# 0.28563f
C20052 a_46268_12135# a_46716_12135# 0.0131f
C20053 a_18740_25156# a_18716_24679# 0.00172f
C20054 a_43940_27912# VPWR 0.20595f
C20055 a_14796_25112# a_14796_24679# 0.05841f
C20056 a_2276_29860# a_1916_29816# 0.08707f
C20057 _381_.Z _412_.A1 0.07887f
C20058 _319_.A2 a_37384_19624# 0.00453f
C20059 _459_.CLK a_32592_25227# 0.00325f
C20060 a_64212_12232# a_64300_10567# 0.00151f
C20061 a_23332_1636# a_23196_1159# 0.00168f
C20062 a_19388_1592# a_19388_1159# 0.05841f
C20063 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN VPWR 0.94334f
C20064 _319_.A3 _323_.A3 1.08502f
C20065 _251_.A1 a_56388_25940# 0.00164f
C20066 _274_.A1 _274_.A2 0.05048f
C20067 a_4852_20072# a_4964_18884# 0.02666f
C20068 _304_.B a_44162_24120# 0.0377f
C20069 a_46716_18407# a_47076_18504# 0.08717f
C20070 a_51868_1159# a_52316_1159# 0.0131f
C20071 _470_.Q _424_.A2 0.16214f
C20072 a_17844_27912# a_18096_27165# 0.0031f
C20073 a_65220_18884# a_65308_18840# 0.28563f
C20074 a_65308_18407# VPWR 0.32585f
C20075 a_5388_27815# a_5300_27912# 0.28563f
C20076 a_4156_25112# VPWR 0.30552f
C20077 a_28372_20452# VPWR 0.20622f
C20078 _476_.Q a_53796_20452# 0.06575f
C20079 a_66340_12612# VPWR 0.2154f
C20080 a_4156_15704# a_4604_15704# 0.01222f
C20081 a_23196_29816# VPWR 0.31469f
C20082 _352_.A2 a_30128_27508# 0.00571f
C20083 _447_.Q a_38228_20452# 0.04167f
C20084 _230_.I a_60404_28292# 0.05969f
C20085 a_55812_15368# a_56260_15368# 0.01328f
C20086 a_40356_15748# a_40220_15271# 0.00168f
C20087 a_17472_28363# a_17844_27912# 0.00113f
C20088 a_19328_28733# a_20308_27912# 0.00172f
C20089 _311_.A2 _304_.A1 1.16034f
C20090 a_67124_10664# VPWR 0.20703f
C20091 a_66204_8999# a_66564_9096# 0.08717f
C20092 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I a_60268_14136# 0.00262f
C20093 a_67100_7431# a_67460_7528# 0.08717f
C20094 a_35180_16839# a_35204_15748# 0.0016f
C20095 a_24540_21543# a_24564_20452# 0.0016f
C20096 _324_.C a_44476_27815# 0.07112f
C20097 _384_.A3 _475_.Q 1.77536f
C20098 a_61300_16936# VPWR 0.14647f
C20099 _438_.ZN _301_.Z 0.0153f
C20100 a_36288_31048# uo_out[2] 0.00141f
C20101 a_40580_15368# VPWR 0.20348f
C20102 _474_.CLK a_53616_29480# 0.00284f
C20103 _230_.I a_61689_29860# 0.0035f
C20104 a_22548_22020# a_22996_22020# 0.01328f
C20105 _304_.B _422_.ZN 0.00112f
C20106 a_44028_15271# VPWR 0.29679f
C20107 _435_.A3 a_40357_24776# 0.00553f
C20108 a_40556_16839# a_41004_16839# 0.01288f
C20109 a_57468_16839# vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I 0.0016f
C20110 a_59652_25640# vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I 0.01593f
C20111 a_48292_26369# VPWR 0.00542f
C20112 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN 0.00359f
C20113 a_67996_17272# VPWR 0.33674f
C20114 a_37444_1256# VPWR 0.20348f
C20115 a_52676_1256# a_53124_1256# 0.01328f
C20116 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I a_65220_20072# 0.00201f
C20117 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN a_55788_24679# 0.00206f
C20118 a_53236_13800# a_53684_13800# 0.01328f
C20119 a_67212_13703# a_67572_13800# 0.08717f
C20120 a_51084_13703# a_51108_12612# 0.0016f
C20121 a_31932_2727# a_32380_2727# 0.0131f
C20122 _395_.A3 a_52434_22504# 0.00109f
C20123 a_43126_24119# _305_.A2 0.01555f
C20124 a_36188_17272# a_36076_16839# 0.02634f
C20125 a_57940_17316# a_58388_17316# 0.01328f
C20126 _346_.B a_21103_29076# 0.00328f
C20127 _241_.Z _243_.ZN 0.39979f
C20128 a_53996_16839# a_54356_16936# 0.08674f
C20129 a_3620_17316# VPWR 0.22347f
C20130 a_13340_1159# a_13252_1256# 0.28563f
C20131 a_53436_1592# a_53572_1256# 0.00168f
C20132 a_52564_16936# VPWR 0.2061f
C20133 a_46940_1592# VPWR 0.3289f
C20134 a_10564_1636# a_10204_1592# 0.08707f
C20135 a_3708_12135# a_3620_12232# 0.28563f
C20136 a_28460_23544# a_28348_23111# 0.02634f
C20137 a_8772_29860# a_9220_29860# 0.01328f
C20138 a_65668_26344# VPWR 0.23875f
C20139 a_31260_17272# a_31708_17272# 0.01288f
C20140 a_35204_17316# a_35292_17272# 0.28563f
C20141 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I 0.05291f
C20142 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I 0.03134f
C20143 a_64996_11044# a_64636_11000# 0.08707f
C20144 a_61052_11000# a_61500_11000# 0.01288f
C20145 a_17508_2824# VPWR 0.20402f
C20146 a_53884_1592# a_54332_1592# 0.01288f
C20147 a_62644_26724# a_62732_26680# 0.28563f
C20148 _459_.CLK a_15156_26724# 0.00299f
C20149 a_29232_29931# uo_out[6] 0.00209f
C20150 _436_.B _435_.A3 0.49654f
C20151 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I a_62980_20072# 0.00201f
C20152 hold2.I a_44906_24164# 0.00212f
C20153 _430_.ZN _441_.B 0.54745f
C20154 _455_.Q a_20308_26724# 0.00218f
C20155 _424_.A2 _260_.A2 0.03993f
C20156 a_19612_23111# a_20060_23111# 0.01288f
C20157 a_44162_24120# VPWR 0.57906f
C20158 a_1916_24679# a_2276_24776# 0.08717f
C20159 a_62560_25112# clk 0.00999f
C20160 _459_.CLK a_23868_26247# 0.05356f
C20161 a_60492_28248# a_60516_27912# 0.00172f
C20162 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_64860_26247# 0.00713f
C20163 a_3620_14180# VPWR 0.22347f
C20164 _474_.CLK a_55252_23588# 0.01491f
C20165 _335_.ZN uo_out[6] 0.1867f
C20166 _223_.ZN uo_out[7] 0.24593f
C20167 VPWR uio_oe[7] 0.27904f
C20168 _459_.CLK a_19035_28409# 0.00193f
C20169 _260_.A1 a_42778_21812# 0.00455f
C20170 a_53324_12135# VPWR 0.31547f
C20171 a_2276_29480# VPWR 0.20634f
C20172 a_36548_15748# a_36188_15704# 0.08707f
C20173 a_32740_2824# a_33188_2824# 0.01328f
C20174 a_30388_28776# _371_.A1 0.10154f
C20175 _304_.B _302_.Z 0.0026f
C20176 a_15692_24679# VPWR 0.29679f
C20177 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I a_58028_20408# 0.00152f
C20178 a_58500_21640# a_58476_20408# 0.0016f
C20179 _452_.CLK a_46268_18407# 0.00274f
C20180 a_23108_21640# a_23220_20452# 0.02666f
C20181 _355_.C a_30796_24463# 0.00501f
C20182 a_38628_25156# VPWR 0.01396f
C20183 a_36100_15748# VPWR 0.20622f
C20184 _427_.ZN _419_.Z 0.00116f
C20185 _260_.ZN a_44038_21236# 0.06227f
C20186 a_2724_9476# a_2364_9432# 0.08717f
C20187 a_4516_9476# a_4964_9476# 0.01328f
C20188 a_29716_22020# a_29356_21976# 0.08663f
C20189 _422_.ZN VPWR 0.42381f
C20190 a_49764_14180# a_49852_14136# 0.28563f
C20191 a_45820_14136# a_46268_14136# 0.01288f
C20192 _241_.Z a_58140_26680# 0.00519f
C20193 a_58476_18840# a_58924_18840# 0.01255f
C20194 _452_.CLK a_44276_17316# 0.00647f
C20195 a_43824_18147# VPWR 0.18611f
C20196 _229_.I a_59620_27208# 0.00126f
C20197 _416_.A1 _284_.A2 0.46773f
C20198 a_47500_16839# VPWR 0.31556f
C20199 a_26108_30951# uio_out[1] 0.00522f
C20200 a_59844_1256# VPWR 0.20348f
C20201 a_58028_13703# a_58052_12612# 0.0016f
C20202 a_47972_13800# a_47972_12612# 0.05841f
C20203 a_67772_14136# a_67684_12612# 0.00151f
C20204 _460_.Q a_34708_29860# 0.00109f
C20205 _475_.Q a_47524_22021# 0.01154f
C20206 _267_.A1 _324_.C 0.85199f
C20207 a_34716_20937# VPWR 0.42252f
C20208 _304_.B a_49764_26724# 0.19767f
C20209 a_37980_17272# VPWR 0.34506f
C20210 a_60740_1636# VPWR 0.20348f
C20211 a_62868_10664# a_62844_9432# 0.0016f
C20212 a_24316_1159# a_24676_1256# 0.08717f
C20213 a_54220_12135# a_54580_12232# 0.08707f
C20214 _325_.A1 a_42896_18504# 0.05206f
C20215 a_17060_1636# a_17508_1636# 0.01328f
C20216 a_15940_29860# a_15580_29816# 0.08663f
C20217 a_54768_22137# VPWR 0.00204f
C20218 a_61188_1636# a_60828_1592# 0.08707f
C20219 a_39908_2824# VPWR 0.20812f
C20220 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN 0.00214f
C20221 a_4068_24776# a_4852_24776# 0.00276f
C20222 a_18716_23111# a_18628_23208# 0.28563f
C20223 a_22300_24679# a_22212_24776# 0.28563f
C20224 _390_.ZN a_52228_27912# 0.04939f
C20225 _330_.A1 a_35268_21640# 0.00233f
C20226 a_46628_9476# VPWR 0.20348f
C20227 _430_.ZN _300_.A2 0.00146f
C20228 a_52540_14136# VPWR 0.34385f
C20229 _388_.B a_48104_30219# 0.00318f
C20230 a_3620_18504# a_4068_18504# 0.01328f
C20231 a_34732_18407# a_35092_18504# 0.0869f
C20232 _459_.CLK uio_out[7] 0.29569f
C20233 a_47076_12232# VPWR 0.20348f
C20234 _260_.ZN _325_.A2 0.00328f
C20235 a_39460_15748# a_39548_15704# 0.28563f
C20236 a_43044_15748# a_43492_15748# 0.01328f
C20237 a_31484_2727# a_31620_1636# 0.00154f
C20238 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_58276_25156# 0.00374f
C20239 _302_.Z VPWR 0.98403f
C20240 a_20420_24776# VPWR 0.20595f
C20241 _243_.A1 _243_.B2 0.02397f
C20242 a_62956_23111# vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I 0.00189f
C20243 _473_.Q _475_.D 0.02802f
C20244 _246_.B2 a_60068_27912# 0.0136f
C20245 _373_.A2 a_29232_29931# 0.00192f
C20246 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN VPWR 0.85077f
C20247 a_4156_2727# a_4740_2824# 0.01675f
C20248 a_30500_21640# a_30388_20452# 0.02666f
C20249 a_61836_25515# a_61748_23588# 0.00146f
C20250 a_22548_28292# _454_.D 0.00512f
C20251 _474_.CLK _404_.A1 0.03293f
C20252 a_42236_15704# VPWR 0.30565f
C20253 a_31260_19975# a_31172_20072# 0.28563f
C20254 _290_.ZN _365_.ZN 0.00117f
C20255 _359_.B a_45800_30345# 0.00152f
C20256 a_56516_26344# VPWR 0.60567f
C20257 vgaringosc.workerclkbuff_notouch_.I a_49112_29885# 0.048f
C20258 a_63516_19975# VPWR 0.31578f
C20259 a_53572_14180# a_53212_14136# 0.08717f
C20260 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN 0.01338f
C20261 _452_.CLK a_37532_26247# 0.00706f
C20262 _452_.CLK a_32828_21543# 0.02062f
C20263 a_55028_13800# a_54916_12612# 0.02666f
C20264 a_2812_12568# a_3260_12568# 0.0131f
C20265 a_54332_2727# a_54780_2727# 0.0131f
C20266 a_64972_13703# a_64996_12612# 0.0016f
C20267 a_36660_23588# _304_.A1 0.00341f
C20268 a_30388_25156# a_30476_25112# 0.28563f
C20269 a_49764_26724# VPWR 0.62648f
C20270 a_35292_26247# VPWR 0.32431f
C20271 a_26160_27165# _457_.D 0.00281f
C20272 a_50076_17272# VPWR 0.33981f
C20273 _327_.A2 a_42896_18504# 0.00843f
C20274 _459_.Q _352_.A2 0.39016f
C20275 a_1380_7528# a_1380_6340# 0.05841f
C20276 a_35740_1159# a_35652_1256# 0.28563f
C20277 a_65420_12135# a_65332_12232# 0.28563f
C20278 a_2812_1159# VPWR 0.30213f
C20279 a_2276_5960# a_2276_4772# 0.05841f
C20280 a_3172_4392# a_3172_3204# 0.05841f
C20281 a_23780_1636# a_24452_1636# 0.00347f
C20282 a_30588_21543# VPWR 0.31547f
C20283 a_47300_17316# a_47388_17272# 0.28563f
C20284 a_50884_17316# a_51332_17316# 0.01328f
C20285 _267_.A2 _267_.ZN 0.11895f
C20286 _424_.A1 _427_.ZN 0.26399f
C20287 _478_.D a_53704_23219# 0.27796f
C20288 a_57828_25156# a_58276_25156# 0.01328f
C20289 a_62308_2824# VPWR 0.20815f
C20290 a_1468_10567# a_1828_10664# 0.08717f
C20291 a_55116_10567# a_55564_10567# 0.01288f
C20292 a_65892_1636# a_65532_1592# 0.08717f
C20293 _324_.C _412_.A1 0.08758f
C20294 _395_.A1 a_50420_23233# 0.00692f
C20295 a_16948_23208# a_17396_23208# 0.01328f
C20296 a_29244_23111# a_29604_23208# 0.08707f
C20297 _474_.CLK vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.0265f
C20298 _251_.A1 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN 0.01418f
C20299 a_57604_9476# VPWR 0.21273f
C20300 _267_.A2 _390_.ZN 0.00652f
C20301 a_61052_14136# VPWR 0.31945f
C20302 a_2364_21543# a_2276_21640# 0.28563f
C20303 a_23644_21543# a_24092_21543# 0.01288f
C20304 a_25572_2824# a_25660_1159# 0.0027f
C20305 a_61860_2824# a_61724_1592# 0.00154f
C20306 a_43003_28409# a_43580_27815# 0.0295f
C20307 a_43296_28733# a_44028_27815# 0.00433f
C20308 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN 0.00711f
C20309 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I 0.62976f
C20310 _337_.A3 a_27588_26344# 0.01401f
C20311 _476_.Q a_51877_21236# 0.00774f
C20312 _285_.Z a_38472_30169# 0.03484f
C20313 a_1380_11044# VPWR 0.20348f
C20314 a_38428_2727# a_38564_1636# 0.00154f
C20315 a_55140_2824# a_55588_2824# 0.01328f
C20316 a_46476_20937# VPWR 0.39673f
C20317 a_20379_29977# uio_out[6] 0.04643f
C20318 a_62172_19975# a_62532_20072# 0.08717f
C20319 _378_.ZN a_17904_28409# 0.00167f
C20320 a_40468_25157# _433_.ZN 0.00194f
C20321 a_2364_18840# VPWR 0.30029f
C20322 a_15580_2727# a_15492_2824# 0.28563f
C20323 _230_.I _248_.B1 0.11414f
C20324 _324_.B a_43156_20452# 0.00165f
C20325 _264_.B a_41476_24776# 0.01211f
C20326 _363_.Z a_31920_29480# 0.03883f
C20327 a_54244_9476# a_54692_9476# 0.01328f
C20328 a_52316_9432# a_52988_9432# 0.00544f
C20329 a_47164_14136# a_47164_13703# 0.05841f
C20330 a_64212_23588# VPWR 0.20944f
C20331 a_61412_14180# a_61860_14180# 0.01328f
C20332 a_51108_14180# a_51084_13703# 0.00172f
C20333 a_3620_20452# a_3708_20408# 0.28563f
C20334 a_25643_25273# a_26132_23588# 0.00146f
C20335 _294_.A2 _452_.CLK 0.00638f
C20336 _260_.A1 hold1.Z 0.00474f
C20337 a_49764_12612# a_49404_12568# 0.08707f
C20338 a_4852_13800# a_4940_12135# 0.00151f
C20339 _230_.I vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN 0.14664f
C20340 a_61972_13800# a_61860_12612# 0.02666f
C20341 a_48708_29816# a_49056_29977# 0.00277f
C20342 _301_.A1 a_38340_21327# 0.39055f
C20343 a_16052_24776# a_16052_23588# 0.05841f
C20344 _459_.Q a_30912_27508# 0.00263f
C20345 a_25212_1159# VPWR 0.32891f
C20346 a_61972_12232# a_62420_12232# 0.01328f
C20347 a_46716_1159# a_47076_1256# 0.08717f
C20348 a_27140_1636# a_27228_1592# 0.28563f
C20349 a_30724_1636# a_31172_1636# 0.01328f
C20350 _452_.Q a_39324_17272# 0.02634f
C20351 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I _324_.C 0.0382f
C20352 _256_.A2 _255_.I 0.80098f
C20353 a_35740_26247# a_35652_26344# 0.28563f
C20354 a_27812_21640# VPWR 0.20614f
C20355 a_40220_20408# a_40668_20408# 0.012f
C20356 a_51956_26183# a_52352_26031# 0.00232f
C20357 a_51556_1636# a_51420_1159# 0.00168f
C20358 a_52428_10567# a_52340_10664# 0.28563f
C20359 _427_.A2 a_52452_21236# 0.37894f
C20360 a_12356_2824# a_12356_1636# 0.05841f
C20361 a_43008_26795# hold2.Z 0.00106f
C20362 a_34844_24679# a_34756_24776# 0.28563f
C20363 _402_.A1 a_42236_27815# 0.00548f
C20364 _304_.B a_43814_21236# 0.10555f
C20365 a_1468_8999# VPWR 0.29679f
C20366 a_17484_23544# VPWR 0.29719f
C20367 a_3260_5863# VPWR 0.30487f
C20368 a_5276_2727# VPWR 0.32932f
C20369 a_55116_13703# VPWR 0.31594f
C20370 a_67348_20072# a_67796_20072# 0.01328f
C20371 a_22300_21543# a_22660_21640# 0.08707f
C20372 a_58687_31220# ui_in[4] 0.05628f
C20373 _351_.A2 _457_.D 0.00347f
C20374 a_50300_11000# VPWR 0.34677f
C20375 a_49180_15704# a_49628_15704# 0.01288f
C20376 a_53124_15748# a_53212_15704# 0.28563f
C20377 _437_.A1 VPWR 2.98249f
C20378 _402_.A1 _284_.B 0.0457f
C20379 a_55340_23544# a_55788_23544# 0.0131f
C20380 a_1468_26680# VPWR 0.29679f
C20381 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_65668_27912# 0.03152f
C20382 _454_.Q _351_.A2 0.03028f
C20383 a_17844_26344# VPWR 0.21215f
C20384 a_49852_30951# vgaringosc.workerclkbuff_notouch_.I 0.00613f
C20385 a_26556_2727# a_26916_2824# 0.08717f
C20386 _245_.Z _245_.I1 0.09286f
C20387 a_63092_26724# vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN 0.00277f
C20388 a_24652_30951# uio_out[3] 0.00741f
C20389 a_65644_23544# clk 0.00613f
C20390 _474_.CLK a_48384_26724# 0.43386f
C20391 a_59844_9476# a_59932_9432# 0.28563f
C20392 a_932_23588# a_1020_23544# 0.28563f
C20393 a_14708_28292# VPWR 0.22532f
C20394 a_61500_26247# a_61860_26344# 0.0869f
C20395 a_1828_4772# a_1916_4728# 0.28563f
C20396 a_2724_3204# a_2812_3160# 0.28563f
C20397 a_54556_14136# a_54668_13703# 0.02634f
C20398 a_17484_20408# a_17932_20408# 0.0131f
C20399 a_56596_23588# a_56236_23544# 0.08717f
C20400 a_6756_1636# VPWR 0.2085f
C20401 _294_.A2 a_31088_30301# 0.0387f
C20402 _459_.CLK a_17396_25156# 0.00249f
C20403 a_56260_12612# a_56708_12612# 0.01328f
C20404 ui_in[2] ui_in[0] 0.00146f
C20405 _223_.I uo_out[6] 0.07788f
C20406 _439_.ZN _438_.ZN 0.0589f
C20407 a_23108_24776# a_22996_23588# 0.02666f
C20408 _416_.A2 a_48084_18884# 0.00301f
C20409 a_47612_1159# VPWR 0.32982f
C20410 a_37888_27555# uo_out[7] 0.00165f
C20411 a_58140_1159# a_58052_1256# 0.28563f
C20412 a_3172_11044# a_3260_11000# 0.28563f
C20413 _409_.ZN _395_.A1 0.00136f
C20414 a_65220_18884# VPWR 0.20921f
C20415 _340_.ZN VPWR 0.45274f
C20416 a_49068_20408# a_50300_20408# 0.00117f
C20417 _452_.CLK a_32268_23544# 0.01794f
C20418 _261_.ZN a_40468_25157# 0.12427f
C20419 a_49204_10664# a_49652_10664# 0.01328f
C20420 a_62956_10567# a_63316_10664# 0.08707f
C20421 a_18044_1159# a_18492_1159# 0.0131f
C20422 a_19300_2824# a_19300_1636# 0.05841f
C20423 a_57044_23588# a_57492_23588# 0.01328f
C20424 _282_.ZN clk 0.00161f
C20425 a_18380_21976# VPWR 0.33639f
C20426 a_43814_21236# VPWR 0.59129f
C20427 a_32180_23588# VPWR 0.2086f
C20428 a_33276_21543# a_33188_21640# 0.28563f
C20429 a_20868_21640# a_21316_21640# 0.01328f
C20430 a_27676_2727# VPWR 0.31879f
C20431 a_49204_13800# VPWR 0.23105f
C20432 a_64412_15271# a_65084_15271# 0.00544f
C20433 _397_.A1 _421_.A1 0.65244f
C20434 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN a_56572_29383# 0.00537f
C20435 _417_.A2 _399_.A1 0.0018f
C20436 a_4604_29816# VPWR 0.32824f
C20437 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I 0.03014f
C20438 _345_.A2 a_23834_28292# 0.0262f
C20439 a_41564_26247# _435_.A3 0.00862f
C20440 a_64100_11044# VPWR 0.2061f
C20441 _304_.B a_52676_27912# 0.05392f
C20442 _304_.A1 a_36860_23111# 0.02827f
C20443 a_15244_23111# VPWR 0.29679f
C20444 _272_.B1 _272_.A2 0.02019f
C20445 _330_.A1 _441_.B 0.03441f
C20446 a_15604_27912# VPWR 0.20789f
C20447 a_64748_23111# a_65668_23208# 0.00795f
C20448 a_25124_28776# a_25740_28776# 0.00817f
C20449 a_62620_17272# a_62532_15748# 0.00151f
C20450 _430_.ZN _452_.Q 0.00609f
C20451 a_37980_2727# a_37892_2824# 0.28563f
C20452 _223_.I uo_out[5] 0.00349f
C20453 _379_.A2 _378_.I 0.57479f
C20454 a_65220_9476# a_65668_9476# 0.01328f
C20455 a_14708_23588# a_14796_23544# 0.28563f
C20456 a_18292_23588# a_18740_23588# 0.01328f
C20457 a_66116_6340# a_66204_6296# 0.28563f
C20458 a_65220_7908# a_65308_7864# 0.28563f
C20459 a_67012_7908# a_67460_7908# 0.01328f
C20460 a_18852_1256# a_19300_1256# 0.01328f
C20461 a_54804_20072# a_55252_20072# 0.01328f
C20462 a_67012_4772# a_67100_4728# 0.28563f
C20463 a_64860_4728# a_65308_4728# 0.0131f
C20464 a_5300_16936# a_5388_15271# 0.0027f
C20465 a_65892_14180# a_65868_13703# 0.00172f
C20466 a_23220_20452# a_23308_20408# 0.28563f
C20467 a_67908_3204# a_67996_3160# 0.28563f
C20468 a_65756_3160# a_66204_3160# 0.0131f
C20469 _275_.A2 _267_.A2 0.00699f
C20470 a_48060_13703# a_48508_13703# 0.0131f
C20471 _393_.A3 _404_.A1 0.44014f
C20472 _459_.Q a_32592_25227# 0.08736f
C20473 _461_.D _223_.ZN 0.00368f
C20474 a_9532_29383# a_9980_29383# 0.0131f
C20475 a_12548_31048# a_12916_31048# 0.02601f
C20476 _460_.Q _335_.ZN 1.37081f
C20477 _375_.Z a_19328_28733# 0.00634f
C20478 a_63516_17272# a_63628_16839# 0.02634f
C20479 a_12892_1592# VPWR 0.29679f
C20480 a_66228_13800# a_66316_12135# 0.00151f
C20481 _319_.ZN _448_.D 0.01586f
C20482 a_1020_30951# a_1468_30951# 0.0131f
C20483 a_37964_18191# a_38308_18559# 0.00275f
C20484 a_47524_31048# vgaringosc.workerclkbuff_notouch_.I 0.00664f
C20485 a_30240_24776# a_31732_23588# 0.00103f
C20486 _359_.B a_32476_29167# 0.03158f
C20487 _244_.Z a_60212_25156# 0.25725f
C20488 a_34732_19975# VPWR 0.36755f
C20489 a_5300_9096# VPWR 0.21406f
C20490 a_65668_5960# VPWR 0.21209f
C20491 a_63764_23588# a_63852_23544# 0.28563f
C20492 a_51108_11044# a_51556_11044# 0.01328f
C20493 _288_.ZN uo_out[4] 0.0218f
C20494 a_47524_11044# a_47612_11000# 0.28563f
C20495 a_36076_18407# VPWR 0.32636f
C20496 a_36860_1592# a_37308_1592# 0.01288f
C20497 a_34644_16936# a_35092_16936# 0.01328f
C20498 _452_.CLK a_32268_21976# 0.02313f
C20499 a_34084_28776# a_35108_28776# 0.00825f
C20500 _437_.A1 a_36996_25156# 0.00254f
C20501 _424_.A2 _476_.Q 0.14975f
C20502 a_44961_27912# _470_.D 0.2404f
C20503 _400_.ZN _397_.A4 0.01247f
C20504 _330_.A1 _328_.A2 0.17608f
C20505 a_38876_19975# a_39324_19975# 0.01255f
C20506 _260_.A2 hold1.Z 1.92974f
C20507 a_27588_26344# a_27328_25227# 0.00187f
C20508 _435_.A3 _433_.ZN 0.00295f
C20509 a_32180_22020# VPWR 0.20757f
C20510 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN 0.00195f
C20511 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN 0.06931f
C20512 a_49852_2727# VPWR 0.34788f
C20513 a_37360_19325# _330_.A2 0.00163f
C20514 a_45596_30951# a_46044_30951# 0.0131f
C20515 a_37844_29860# VPWR 0.01469f
C20516 a_3172_12612# VPWR 0.20993f
C20517 a_1828_26344# a_2276_26344# 0.01328f
C20518 a_16140_26247# a_16500_26344# 0.08717f
C20519 a_64884_16936# a_65084_15271# 0.00119f
C20520 a_25796_27912# a_25867_26841# 0.00126f
C20521 _359_.B a_34532_27208# 0.00373f
C20522 _475_.Q a_49856_20936# 0.00198f
C20523 a_16700_29816# VPWR 0.30141f
C20524 a_53884_20408# a_54332_20408# 0.01255f
C20525 _384_.ZN _384_.A3 0.04583f
C20526 a_51084_10567# VPWR 0.31389f
C20527 a_35068_15271# a_35428_15368# 0.08717f
C20528 a_52676_27912# VPWR 0.20816f
C20529 a_3620_23208# VPWR 0.22347f
C20530 _350_.A1 a_35740_30951# 0.01422f
C20531 _439_.ZN a_39332_23588# 0.00121f
C20532 a_3172_28292# a_3620_28292# 0.01328f
C20533 a_1380_28292# a_1020_28248# 0.08717f
C20534 a_48956_2727# a_49316_2824# 0.08717f
C20535 a_1828_22020# a_1916_21976# 0.28563f
C20536 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I 0.0331f
C20537 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I 0.0834f
C20538 a_65220_17316# a_65308_17272# 0.28563f
C20539 _346_.A2 a_21964_25112# 0.00112f
C20540 a_3620_16936# a_3620_15748# 0.05841f
C20541 _267_.ZN vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.01696f
C20542 _304_.B vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN 0.13585f
C20543 a_56572_23111# a_56932_23208# 0.08663f
C20544 a_16948_25156# a_17396_25156# 0.01328f
C20545 _324_.C a_43296_28733# 0.01218f
C20546 _393_.ZN a_46804_28292# 0.00297f
C20547 a_45372_13703# a_45284_13800# 0.28563f
C20548 a_28460_20408# a_28908_20408# 0.0131f
C20549 a_56148_24776# a_56148_23588# 0.05841f
C20550 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_62196_23588# 0.00747f
C20551 _260_.ZN _302_.Z 0.07174f
C20552 input9.Z _268_.A1 0.48812f
C20553 a_21204_31048# a_20672_30301# 0.02391f
C20554 a_32156_16839# a_32068_16936# 0.28563f
C20555 _419_.Z a_51240_20452# 0.4546f
C20556 _390_.ZN vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.21639f
C20557 a_62844_12568# a_63292_12568# 0.01288f
C20558 a_66788_12612# a_66428_12568# 0.08707f
C20559 a_26692_1636# VPWR 0.21618f
C20560 a_51050_29480# VPWR 0.0145f
C20561 _324_.C _473_.Q 0.02381f
C20562 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I 0.09391f
C20563 _272_.A2 VPWR 0.31553f
C20564 _474_.CLK _419_.Z 0.00188f
C20565 _388_.B a_44795_29535# 0.00934f
C20566 a_44164_1636# a_43804_1592# 0.08707f
C20567 a_53236_12232# a_53324_10567# 0.00151f
C20568 _417_.Z a_50212_20452# 0.00663f
C20569 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN VPWR 0.72643f
C20570 _424_.B1 _284_.B 0.00199f
C20571 _362_.B a_34348_27208# 0.00498f
C20572 _441_.B _300_.ZN 0.01157f
C20573 _265_.ZN _435_.A3 0.01976f
C20574 _244_.Z VPWR 0.51503f
C20575 _470_.Q a_47376_27912# 0.00513f
C20576 _251_.A1 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN 0.30901f
C20577 a_40444_1159# a_40892_1159# 0.0131f
C20578 _324_.C a_42996_18840# 0.00181f
C20579 a_53548_24679# a_53460_24776# 0.28563f
C20580 a_16948_20452# VPWR 0.20348f
C20581 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN 0.00108f
C20582 a_34440_25273# VPWR 0.00232f
C20583 _226_.ZN _328_.A2 0.0025f
C20584 a_56684_17272# vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN 0.02616f
C20585 _400_.ZN a_44864_27165# 0.02049f
C20586 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN 0.79633f
C20587 a_64884_16936# a_65332_16936# 0.01328f
C20588 a_52092_12568# VPWR 0.31547f
C20589 _359_.B a_45088_29123# 0.20417f
C20590 _284_.ZN a_43232_29480# 0.00357f
C20591 a_44388_15368# a_44836_15368# 0.01328f
C20592 a_7964_29383# a_7876_29480# 0.28563f
C20593 a_5276_30951# uio_oe[7] 0.00148f
C20594 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN 0.09039f
C20595 _416_.A1 _419_.A4 0.03614f
C20596 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN 0.80656f
C20597 a_5300_10664# VPWR 0.21406f
C20598 a_46492_15271# a_46404_15368# 0.28563f
C20599 a_66652_2727# a_66788_1636# 0.00154f
C20600 _384_.A1 _324_.B 0.0018f
C20601 a_35140_26680# a_35756_27216# 0.00478f
C20602 _260_.A1 a_42252_20936# 0.04298f
C20603 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN 0.00775f
C20604 a_47836_15271# a_48284_15271# 0.0131f
C20605 a_39264_18147# VPWR 0.51496f
C20606 _383_.A2 _381_.Z 0.14548f
C20607 a_50792_26344# _412_.B2 0.31441f
C20608 a_15604_22020# a_15692_21976# 0.28563f
C20609 a_60380_2727# a_60292_2824# 0.28563f
C20610 a_19188_22020# a_19636_22020# 0.01328f
C20611 a_63964_15704# VPWR 0.29679f
C20612 a_23627_27967# VPWR 0.3712f
C20613 a_4156_16839# a_4940_16839# 0.00443f
C20614 a_44700_30951# a_44612_31048# 0.28563f
C20615 a_40332_21543# a_40780_21543# 0.01222f
C20616 _303_.ZN _438_.ZN 0.02728f
C20617 a_37332_16936# a_37444_15748# 0.02666f
C20618 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN VPWR 1.34821f
C20619 a_25796_23208# a_25884_21543# 0.00151f
C20620 a_41252_1256# a_41700_1256# 0.01328f
C20621 _334_.A1 uo_out[2] 0.06327f
C20622 _417_.A2 a_49448_20072# 0.12262f
C20623 a_25772_23544# a_26220_23544# 0.01255f
C20624 a_4156_7864# VPWR 0.30552f
C20625 a_14596_1256# VPWR 0.20348f
C20626 a_64772_4772# VPWR 0.20727f
C20627 _355_.B VPWR 0.47347f
C20628 a_54192_22851# a_54088_22895# 0.10745f
C20629 a_56012_13703# a_56372_13800# 0.08663f
C20630 a_53212_14136# a_53124_12612# 0.00151f
C20631 a_2276_13800# a_2724_13800# 0.01328f
C20632 a_5276_29383# VPWR 0.3289f
C20633 a_20508_2727# a_20956_2727# 0.0131f
C20634 _350_.A1 a_29563_29535# 0.01249f
C20635 _475_.D _416_.ZN 0.00633f
C20636 a_61076_20452# a_61164_20408# 0.28563f
C20637 a_3708_17272# a_3708_16839# 0.05841f
C20638 a_64324_29860# a_64412_29816# 0.28563f
C20639 _435_.A3 _261_.ZN 0.04306f
C20640 _417_.A2 a_52920_22760# 0.00105f
C20641 _330_.A1 a_40092_27209# 0.01024f
C20642 _450_.D a_41776_18504# 0.00121f
C20643 a_43020_16839# a_43380_16936# 0.08707f
C20644 a_58476_10567# a_58500_9476# 0.0016f
C20645 _452_.Q _441_.A3 0.46054f
C20646 a_1916_1159# a_1828_1256# 0.28563f
C20647 a_5300_16936# VPWR 0.21406f
C20648 a_32828_1592# VPWR 0.29679f
C20649 a_43492_27912# VPWR 0.20795f
C20650 a_20620_23544# a_20508_23111# 0.02634f
C20651 a_7204_1636# a_6844_1592# 0.08707f
C20652 a_1828_29860# a_1916_29816# 0.28563f
C20653 a_5412_29860# a_5860_29860# 0.01328f
C20654 _272_.B1 _228_.ZN 0.00582f
C20655 a_2812_17272# a_3260_17272# 0.0131f
C20656 _424_.B1 _474_.D 0.09252f
C20657 a_48104_30219# a_48708_29816# 0.49241f
C20658 a_50660_1636# a_51108_1636# 0.01328f
C20659 a_57244_11000# a_57692_11000# 0.01288f
C20660 a_58612_16936# vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I 0.00501f
C20661 vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I a_67124_20452# 0.00249f
C20662 _327_.Z a_40644_17272# 0.00938f
C20663 _402_.ZN _402_.B 0.20844f
C20664 _304_.B a_43750_23544# 0.06163f
C20665 _438_.A2 _441_.A2 0.00246f
C20666 _251_.A1 vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN 0.00105f
C20667 a_42896_18504# a_43284_18191# 0.00393f
C20668 a_57580_18407# a_58252_18407# 0.00544f
C20669 a_46716_18407# a_46628_18504# 0.28563f
C20670 a_43716_31048# _480_.Q 0.00167f
C20671 a_48420_18504# a_48396_16839# 0.00131f
C20672 a_37384_19624# a_37772_19759# 0.00334f
C20673 _470_.Q a_46198_27060# 0.07125f
C20674 _300_.ZN _300_.A2 0.15797f
C20675 a_65220_18884# a_64860_18840# 0.08717f
C20676 a_64860_18407# VPWR 0.30145f
C20677 a_3708_25112# VPWR 0.33374f
C20678 a_19948_27815# a_20396_27815# 0.012f
C20679 _274_.A3 a_52640_29860# 0.02369f
C20680 a_27924_20452# VPWR 0.20622f
C20681 a_4940_27815# a_5300_27912# 0.08674f
C20682 _424_.A1 a_51240_20452# 0.3552f
C20683 _476_.Q a_52136_20936# 0.00146f
C20684 a_65892_12612# VPWR 0.23512f
C20685 a_64660_23208# vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN 0.03996f
C20686 _352_.A2 a_29736_27508# 0.00751f
C20687 a_21316_2824# a_21764_2824# 0.01328f
C20688 a_45732_18504# a_45620_17316# 0.02666f
C20689 _475_.Q _417_.Z 0.23487f
C20690 _474_.CLK _424_.A1 0.08864f
C20691 a_66204_8999# a_66116_9096# 0.28563f
C20692 a_66676_10664# VPWR 0.20704f
C20693 a_54804_24776# a_55252_24776# 0.01328f
C20694 a_67100_7431# a_67012_7528# 0.28563f
C20695 _355_.B a_28903_24776# 0.09809f
C20696 _412_.B2 _281_.ZN 0.00139f
C20697 a_932_5960# a_932_4772# 0.05841f
C20698 a_15604_21640# a_15604_20452# 0.05841f
C20699 _324_.C a_44028_27815# 0.01853f
C20700 a_40132_15368# VPWR 0.20348f
C20701 a_43580_15271# VPWR 0.29679f
C20702 a_2812_14136# a_3260_14136# 0.0131f
C20703 a_67548_17272# VPWR 0.31547f
C20704 a_44276_16936# a_44388_15748# 0.02666f
C20705 a_40468_16936# a_40444_15704# 0.0016f
C20706 a_36996_1256# VPWR 0.20348f
C20707 _251_.A1 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN 0.00971f
C20708 a_65756_3160# a_65756_2727# 0.05841f
C20709 a_67212_13703# a_67124_13800# 0.28563f
C20710 a_42796_23981# _305_.A2 0.01388f
C20711 a_53996_16839# a_53908_16936# 0.28563f
C20712 _324_.C _381_.Z 0.59692f
C20713 a_3172_17316# VPWR 0.20993f
C20714 a_46492_1592# VPWR 0.32824f
C20715 a_21628_28248# _455_.D 0.00259f
C20716 a_52116_16936# VPWR 0.2061f
C20717 a_12892_1159# a_13252_1256# 0.08717f
C20718 a_6084_29480# a_6532_29480# 0.01328f
C20719 a_3260_12135# a_3620_12232# 0.08717f
C20720 a_10116_1636# a_10204_1592# 0.28563f
C20721 a_13700_1636# a_14148_1636# 0.01328f
C20722 a_57132_12135# a_57580_12135# 0.01288f
C20723 a_24080_25227# a_25884_24679# 0.00456f
C20724 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN VPWR 0.71795f
C20725 a_35204_17316# a_34844_17272# 0.08707f
C20726 a_43268_31048# a_43716_31048# 0.01328f
C20727 a_64548_11044# a_64636_11000# 0.28563f
C20728 _438_.A2 a_39772_19975# 0.0021f
C20729 _416_.ZN a_47252_18884# 0.0018f
C20730 a_17060_2824# VPWR 0.20348f
C20731 a_62644_26724# a_62284_26680# 0.0869f
C20732 _455_.Q a_19860_26724# 0.00107f
C20733 _430_.ZN a_38759_24072# 0.0052f
C20734 a_43750_23544# VPWR 0.74963f
C20735 _398_.C _399_.A2 0.24945f
C20736 _459_.CLK a_23420_26247# 0.01837f
C20737 a_1916_24679# a_1828_24776# 0.28563f
C20738 a_19612_24679# a_20060_24679# 0.01288f
C20739 a_2364_19975# a_2812_19975# 0.0131f
C20740 a_61836_25515# clk 0.01079f
C20741 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN 0.39913f
C20742 a_62844_1159# a_63292_1159# 0.0131f
C20743 a_47524_2824# a_47388_1592# 0.00154f
C20744 uio_oe[5] uio_oe[4] 0.05732f
C20745 a_3172_14180# VPWR 0.20993f
C20746 _474_.CLK a_54804_23588# 0.00539f
C20747 a_25643_25273# VPWR 0.38121f
C20748 a_3708_18407# a_4156_18407# 0.0131f
C20749 _404_.A1 a_45577_27509# 0.0021f
C20750 _459_.CLK a_16588_28248# 0.02549f
C20751 _260_.A1 a_42154_21236# 0.02101f
C20752 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I 0.02069f
C20753 _260_.A2 clkbuf_1_0__f_clk.I 0.02942f
C20754 a_36100_15748# a_36188_15704# 0.28563f
C20755 a_32156_15704# a_32604_15704# 0.01288f
C20756 a_1828_29480# VPWR 0.20348f
C20757 a_52876_12135# VPWR 0.33016f
C20758 a_53460_18504# a_53572_17316# 0.02666f
C20759 _275_.A2 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.00603f
C20760 a_42982_21730# a_43254_21236# 0.0013f
C20761 _228_.ZN VPWR 0.42187f
C20762 a_15244_24679# VPWR 0.29679f
C20763 a_20308_27912# uio_out[7] 0.00132f
C20764 _452_.CLK a_45820_18407# 0.0062f
C20765 a_42368_28733# a_43003_28409# 0.02112f
C20766 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.09632f
C20767 a_35652_15748# VPWR 0.20622f
C20768 a_47259_20127# a_47636_18884# 0.0306f
C20769 _260_.ZN a_43814_21236# 0.05098f
C20770 a_47612_18407# a_48060_18407# 0.0131f
C20771 a_2276_9476# a_2364_9432# 0.28563f
C20772 _470_.Q a_46580_28292# 0.00117f
C20773 a_25324_21976# a_25772_21976# 0.01288f
C20774 a_51108_21640# VPWR 0.14544f
C20775 _228_.ZN a_59332_29816# 0.00312f
C20776 a_29268_22020# a_29356_21976# 0.28563f
C20777 _218_.ZN _474_.D 0.59323f
C20778 _473_.Q _281_.A1 0.00242f
C20779 a_49764_14180# a_49404_14136# 0.08707f
C20780 a_42896_18504# VPWR 1.11538f
C20781 a_51308_16839# a_51756_16839# 0.0131f
C20782 a_18400_28733# a_18028_28777# 0.10745f
C20783 _452_.CLK a_40644_17272# 0.00906f
C20784 a_47412_16936# a_47388_15704# 0.0016f
C20785 _229_.I a_59260_26680# 0.00111f
C20786 a_51220_16936# a_51332_15748# 0.02666f
C20787 a_47052_16839# VPWR 0.31556f
C20788 a_63652_1256# a_64100_1256# 0.01328f
C20789 a_25652_31048# uio_out[1] 0.0031f
C20790 a_59396_1256# VPWR 0.20348f
C20791 a_61412_26344# vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN 0.00132f
C20792 a_42908_2727# a_43356_2727# 0.0131f
C20793 a_55364_21640# a_55228_20408# 0.00154f
C20794 a_63764_13800# a_64212_13800# 0.01328f
C20795 a_35088_20893# VPWR 0.20719f
C20796 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN a_64972_26680# 0.01208f
C20797 _350_.A1 VPWR 1.91405f
C20798 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN 0.0124f
C20799 a_45708_17272# a_45708_16839# 0.05841f
C20800 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I 0.71013f
C20801 a_37532_17272# VPWR 0.31547f
C20802 _237_.A1 a_59948_30352# 0.00119f
C20803 a_38228_20452# _319_.A2 0.05239f
C20804 a_60292_1636# VPWR 0.20348f
C20805 _319_.ZN a_34592_20569# 0.00247f
C20806 a_24316_1159# a_24228_1256# 0.28563f
C20807 a_39684_20452# a_40132_20452# 0.01328f
C20808 a_54220_12135# a_54132_12232# 0.28563f
C20809 _424_.B1 _474_.Q 0.18895f
C20810 a_11548_29816# a_11996_29816# 0.01288f
C20811 a_15492_29860# a_15580_29816# 0.28563f
C20812 a_67996_21976# VPWR 0.35182f
C20813 a_1828_26344# a_1828_25156# 0.05841f
C20814 _258_.ZN a_57244_27815# 0.00123f
C20815 _330_.A1 _452_.Q 0.04143f
C20816 _336_.A2 a_27564_23544# 0.00412f
C20817 a_40644_17272# a_41040_17801# 0.00232f
C20818 a_4156_10567# a_4940_10567# 0.00443f
C20819 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_59820_14136# 0.00255f
C20820 _474_.CLK input9.Z 0.46895f
C20821 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I 0.00529f
C20822 a_39460_2824# VPWR 0.20348f
C20823 a_60740_1636# a_60828_1592# 0.28563f
C20824 a_56796_1592# a_57244_1592# 0.01288f
C20825 a_33276_1592# a_33276_1159# 0.05841f
C20826 a_37220_1636# a_37084_1159# 0.00168f
C20827 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN a_56796_15271# 0.02334f
C20828 _294_.ZN a_31920_29480# 0.03233f
C20829 _459_.CLK _346_.ZN 0.01192f
C20830 a_17932_23111# a_18628_23208# 0.01227f
C20831 a_30140_23111# a_30588_23111# 0.01288f
C20832 _441_.A3 a_40357_24776# 0.06035f
C20833 _330_.A1 a_35044_21640# 0.02019f
C20834 a_21852_24679# a_22212_24776# 0.08707f
C20835 a_41564_24679# a_41476_24776# 0.28563f
C20836 a_46180_9476# VPWR 0.20348f
C20837 a_3260_21543# a_3708_21543# 0.0131f
C20838 a_52092_14136# VPWR 0.31547f
C20839 a_34732_18407# a_34644_18504# 0.28563f
C20840 _388_.B a_45904_30180# 0.00916f
C20841 a_7092_31048# a_7204_29860# 0.02666f
C20842 a_39460_15748# a_39100_15704# 0.08707f
C20843 _384_.A3 a_51576_25896# 0.05681f
C20844 a_46628_12232# VPWR 0.20348f
C20845 _274_.A3 _324_.C 0.00212f
C20846 a_52316_15704# a_52452_15368# 0.00168f
C20847 a_43716_2824# a_44164_2824# 0.01328f
C20848 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I a_57828_25156# 0.05921f
C20849 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN a_58476_13703# 0.00404f
C20850 a_1916_20408# a_1916_19975# 0.05841f
C20851 a_54244_15748# a_54108_15271# 0.00168f
C20852 a_19972_24776# VPWR 0.20631f
C20853 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN 0.62578f
C20854 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I 0.00151f
C20855 a_42392_19243# a_43400_18909# 0.02307f
C20856 a_4156_2727# a_4068_2824# 0.28563f
C20857 a_41788_15704# VPWR 0.3357f
C20858 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I 0.02402f
C20859 a_30812_19975# a_31172_20072# 0.08717f
C20860 a_61500_26247# a_61948_26247# 0.01255f
C20861 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_62944_29101# 0.00171f
C20862 vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN a_57132_18407# 0.00146f
C20863 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN 0.03961f
C20864 a_46716_9432# a_47164_9432# 0.0131f
C20865 a_48420_9476# a_49092_9476# 0.00347f
C20866 a_63068_19975# VPWR 0.31581f
C20867 a_53124_14180# a_53212_14136# 0.28563f
C20868 a_56260_14180# a_56708_14180# 0.01328f
C20869 _452_.CLK a_37084_26247# 0.00706f
C20870 a_19276_25112# a_19188_23588# 0.00151f
C20871 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I a_56596_18504# 0.00467f
C20872 _452_.CLK a_32380_21543# 0.00287f
C20873 a_4964_12612# a_5052_12568# 0.28563f
C20874 a_52764_17272# a_52652_16839# 0.02634f
C20875 a_36212_23588# _304_.A1 0.12875f
C20876 _384_.A3 a_51540_23588# 0.00173f
C20877 a_33396_26344# VPWR 0.00438f
C20878 a_49628_17272# VPWR 0.32012f
C20879 a_35292_1159# a_35652_1256# 0.08717f
C20880 a_2364_1159# VPWR 0.30029f
C20881 a_19836_1592# a_20284_1592# 0.01288f
C20882 a_23780_1636# a_23868_1592# 0.28563f
C20883 a_64972_12135# a_65332_12232# 0.08717f
C20884 a_50996_12232# a_51444_12232# 0.01328f
C20885 _256_.A2 ena 0.01057f
C20886 a_30140_21543# VPWR 0.33016f
C20887 a_19524_26344# a_19636_25156# 0.02666f
C20888 _311_.A2 _301_.A1 0.22423f
C20889 a_43246_23610# VPWR 0.00449f
C20890 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_63316_23208# 0.00117f
C20891 a_47300_17316# a_46940_17272# 0.08707f
C20892 a_1468_10567# a_1380_10664# 0.28563f
C20893 a_65444_1636# a_65532_1592# 0.28563f
C20894 a_61860_2824# VPWR 0.22891f
C20895 _243_.A1 a_58052_26724# 0.00234f
C20896 _395_.A1 a_48321_23208# 0.00161f
C20897 a_47271_21640# _475_.D 0.07669f
C20898 a_29244_23111# a_29156_23208# 0.28563f
C20899 a_24004_24776# a_24452_24776# 0.01328f
C20900 a_57156_9476# VPWR 0.21061f
C20901 _452_.Q _226_.ZN 0.03823f
C20902 a_1916_21543# a_2276_21640# 0.08717f
C20903 hold1.Z a_44500_22020# 0.00365f
C20904 a_67684_14180# VPWR 0.20893f
C20905 a_60276_29032# a_60916_29612# 0.0101f
C20906 _252_.ZN a_60656_29612# 0.00759f
C20907 _398_.C a_54804_23588# 0.00114f
C20908 _304_.B a_43736_25896# 0.09968f
C20909 a_43296_28733# a_43580_27815# 0.00139f
C20910 a_45820_15704# a_46404_15748# 0.01675f
C20911 a_932_11044# VPWR 0.22176f
C20912 _229_.I a_63336_29480# 0.12178f
C20913 a_9220_29860# a_9084_29383# 0.00168f
C20914 a_62172_19975# a_62084_20072# 0.28563f
C20915 a_46848_20893# VPWR 0.18781f
C20916 a_64860_18840# a_64860_18407# 0.05841f
C20917 a_37464_24831# VPWR 0.00204f
C20918 _330_.A2 a_38764_16839# 0.00123f
C20919 _303_.ZN a_40692_21640# 0.00501f
C20920 _276_.A2 _390_.ZN 0.00211f
C20921 a_1916_18840# VPWR 0.297f
C20922 _459_.D a_30672_24831# 0.00242f
C20923 _424_.B1 _395_.A2 0.30161f
C20924 a_15132_2727# a_15492_2824# 0.08717f
C20925 _452_.Q _300_.ZN 0.037f
C20926 a_44744_26355# a_45664_26031# 0.00306f
C20927 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I VPWR 0.7326f
C20928 a_67436_19975# a_67884_19975# 0.012f
C20929 a_16612_29860# uio_oe[0] 0.0058f
C20930 _251_.A1 _231_.ZN 0.26477f
C20931 _264_.B a_40973_24776# 0.00127f
C20932 _474_.Q _218_.ZN 0.6022f
C20933 _302_.Z a_39796_22504# 0.283f
C20934 _402_.ZN a_46352_22021# 0.09202f
C20935 a_63764_23588# VPWR 0.20632f
C20936 a_50076_17272# a_49988_15748# 0.0027f
C20937 a_1020_20408# a_1468_20408# 0.0131f
C20938 a_3620_20452# a_3260_20408# 0.08717f
C20939 _294_.A2 a_35874_27937# 0.0068f
C20940 _336_.Z a_30476_23544# 0.00138f
C20941 _474_.CLK _411_.A2 0.33966f
C20942 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN 0.00179f
C20943 a_65084_2727# a_65756_2727# 0.00544f
C20944 a_45372_12568# a_45820_12568# 0.01288f
C20945 _301_.A1 a_37444_21640# 0.0072f
C20946 a_49316_12612# a_49404_12568# 0.28563f
C20947 _255_.I _238_.ZN 0.0186f
C20948 a_24764_1159# VPWR 0.3289f
C20949 a_67460_9096# a_67460_7908# 0.05841f
C20950 a_46716_1159# a_46628_1256# 0.28563f
C20951 a_45732_12232# a_45732_11044# 0.05841f
C20952 a_33860_20072# a_34644_20072# 0.00276f
C20953 a_65532_12568# a_65444_11044# 0.00151f
C20954 a_27140_1636# a_26780_1592# 0.08707f
C20955 a_5300_4392# a_5276_2727# 0.00144f
C20956 _452_.Q a_40040_17675# 0.37217f
C20957 _256_.A2 a_60401_30300# 0.01293f
C20958 a_27364_21640# VPWR 0.22365f
C20959 a_35292_26247# a_35652_26344# 0.0869f
C20960 _352_.ZN _355_.ZN 0.00672f
C20961 a_53660_17272# vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN 0.0031f
C20962 a_51980_10567# a_52340_10664# 0.08707f
C20963 a_65868_10567# a_66316_10567# 0.0131f
C20964 a_6620_1159# a_7068_1159# 0.0131f
C20965 vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN VPWR 0.72828f
C20966 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN 0.63553f
C20967 a_27812_23208# a_28260_23208# 0.01328f
C20968 a_34396_24679# a_34756_24776# 0.08674f
C20969 _402_.A1 a_41228_27815# 0.00709f
C20970 a_22300_21543# a_22212_21640# 0.28563f
C20971 a_21424_25987# a_21404_24679# 0.00112f
C20972 a_17036_23544# VPWR 0.29679f
C20973 a_1020_8999# VPWR 0.30073f
C20974 a_2812_5863# VPWR 0.30213f
C20975 _459_.CLK _371_.A3 0.05047f
C20976 a_36548_2824# a_36636_1159# 0.0027f
C20977 a_54668_13703# VPWR 0.31594f
C20978 a_4828_2727# VPWR 0.33394f
C20979 a_43736_25896# VPWR 0.67516f
C20980 _304_.B _417_.A2 0.00416f
C20981 _390_.ZN _395_.A1 0.68948f
C20982 _384_.A1 a_49604_22020# 0.01673f
C20983 a_49852_11000# VPWR 0.32357f
C20984 a_53124_15748# a_52764_15704# 0.08707f
C20985 a_1468_21976# a_1468_21543# 0.05841f
C20986 a_66116_2824# a_66564_2824# 0.01328f
C20987 a_1020_26680# VPWR 0.30073f
C20988 a_12548_31048# a_12444_29816# 0.0016f
C20989 _454_.Q a_24900_27912# 0.0665f
C20990 a_31820_20408# a_31708_19975# 0.02634f
C20991 a_63428_15748# a_63876_15748# 0.01328f
C20992 a_25867_26841# a_26112_27209# 0.00232f
C20993 a_17396_26344# VPWR 0.20348f
C20994 a_49404_30951# vgaringosc.workerclkbuff_notouch_.I 0.00613f
C20995 a_26556_2727# a_26468_2824# 0.28563f
C20996 _324_.B _416_.A3 0.79062f
C20997 _245_.Z a_62308_26344# 0.00773f
C20998 _267_.A2 _238_.I 0.39713f
C20999 a_24196_31048# uio_out[3] 0.0965f
C21000 a_65196_23544# clk 0.00613f
C21001 _451_.Q a_41642_25156# 0.0087f
C21002 a_7428_1256# a_7876_1256# 0.01328f
C21003 a_5052_28248# VPWR 0.33516f
C21004 a_1828_7908# a_2276_7908# 0.01328f
C21005 a_2724_23588# a_3172_23588# 0.01328f
C21006 a_59844_9476# a_59484_9432# 0.08717f
C21007 a_57692_9432# a_58140_9432# 0.0131f
C21008 _363_.Z uo_out[6] 0.45292f
C21009 a_10004_31048# a_10452_31048# 0.01328f
C21010 a_61500_26247# a_61412_26344# 0.28563f
C21011 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN 0.89113f
C21012 _436_.B _330_.A1 0.16016f
C21013 a_2724_6340# a_3172_6340# 0.01328f
C21014 a_2724_3204# a_2364_3160# 0.08717f
C21015 a_4516_3204# a_4964_3204# 0.01328f
C21016 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN 0.04756f
C21017 a_1828_4772# a_1468_4728# 0.08717f
C21018 a_3620_4772# a_4068_4772# 0.01328f
C21019 a_64636_14136# a_65084_14136# 0.01288f
C21020 a_31372_21976# a_31284_20452# 0.00151f
C21021 a_36148_21976# _317_.A2 0.17084f
C21022 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN 0.00139f
C21023 a_56148_23588# a_56236_23544# 0.28563f
C21024 _459_.CLK uo_out[7] 1.25465f
C21025 a_6308_1636# VPWR 0.2085f
C21026 a_55028_13800# a_55116_12135# 0.00151f
C21027 _459_.CLK a_16948_25156# 0.00249f
C21028 a_31396_31048# uo_out[6] 0.00872f
C21029 a_43008_26795# _284_.A2 0.01514f
C21030 a_57468_1159# a_58052_1256# 0.01675f
C21031 _416_.A2 a_47636_18884# 0.01558f
C21032 a_7292_29816# a_7428_29480# 0.00168f
C21033 a_47164_1159# VPWR 0.3289f
C21034 a_3172_11044# a_2812_11000# 0.08717f
C21035 a_64772_18884# VPWR 0.20727f
C21036 a_65420_16839# a_66092_16839# 0.00544f
C21037 a_33636_1636# a_34084_1636# 0.01328f
C21038 a_49068_20408# a_49856_20936# 0.00403f
C21039 a_43580_27815# a_44028_27815# 0.01222f
C21040 a_24952_29032# a_25340_29167# 0.00334f
C21041 _452_.CLK a_31820_23544# 0.0036f
C21042 _261_.ZN a_40084_25156# 0.00188f
C21043 a_35740_25112# a_35616_24776# 0.00156f
C21044 a_62956_10567# a_62868_10664# 0.28563f
C21045 _459_.CLK _480_.Q 0.00171f
C21046 a_17932_21976# VPWR 0.30035f
C21047 _395_.A2 _218_.ZN 0.00154f
C21048 a_43666_21812# VPWR 0.00401f
C21049 a_31732_23588# VPWR 0.20368f
C21050 _350_.A1 _370_.B 0.06018f
C21051 a_32828_21543# a_33188_21640# 0.08707f
C21052 a_27004_2727# VPWR 0.37622f
C21053 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN 0.79189f
C21054 a_48420_13800# VPWR 0.20924f
C21055 a_31172_18884# a_31620_18884# 0.01328f
C21056 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN 0.03117f
C21057 a_1020_26247# a_1468_26247# 0.0131f
C21058 a_29184_25597# a_29716_23588# 0.0012f
C21059 _417_.A2 VPWR 2.49204f
C21060 a_4156_29816# VPWR 0.30551f
C21061 a_41116_26247# _435_.A3 0.01771f
C21062 a_21428_22020# a_21404_21543# 0.00172f
C21063 a_63652_11044# VPWR 0.20595f
C21064 a_17484_21976# a_17484_21543# 0.05841f
C21065 a_14796_23111# VPWR 0.30073f
C21066 _284_.B a_46794_25156# 0.00253f
C21067 _243_.ZN a_58656_27912# 0.00156f
C21068 a_52316_2727# a_52452_1636# 0.00154f
C21069 _363_.Z uo_out[5] 0.21849f
C21070 _304_.B a_52228_27912# 0.02062f
C21071 a_45088_29123# a_45396_28292# 0.0022f
C21072 a_61748_23588# vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I 0.00465f
C21073 a_57120_31048# _272_.A2 0.00115f
C21074 _250_.ZN a_61948_27815# 0.00161f
C21075 a_15156_27912# VPWR 0.20348f
C21076 _330_.A1 a_38759_24072# 0.00493f
C21077 a_25124_28776# a_25332_28776# 0.00733f
C21078 a_37532_2727# a_37892_2824# 0.08717f
C21079 a_38616_24328# _452_.Q 0.00167f
C21080 a_65220_7908# a_64860_7864# 0.08717f
C21081 a_1916_7864# a_1916_7431# 0.05841f
C21082 VPWR ui_in[3] 0.49121f
C21083 a_1380_25156# a_1828_25156# 0.01328f
C21084 a_66116_6340# a_65756_6296# 0.08717f
C21085 a_2812_6296# a_2812_5863# 0.05841f
C21086 a_39684_26344# _436_.ZN 0.00131f
C21087 a_5052_14136# a_4964_12612# 0.00151f
C21088 a_61948_14136# a_62060_13703# 0.02634f
C21089 a_3708_4728# a_3708_4295# 0.05841f
C21090 a_67012_4772# a_66652_4728# 0.08717f
C21091 a_67908_3204# a_67548_3160# 0.08663f
C21092 a_62980_20072# a_62980_18884# 0.05841f
C21093 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I VPWR 0.77559f
C21094 a_24564_20452# a_25012_20452# 0.01328f
C21095 a_23220_20452# a_22860_20408# 0.08717f
C21096 a_67460_17316# a_67436_16839# 0.00172f
C21097 a_11548_30951# a_12916_31048# 0.00207f
C21098 a_12548_31048# a_11460_31048# 0.00174f
C21099 _424_.B1 _427_.A2 0.00513f
C21100 _411_.A2 _398_.C 0.11163f
C21101 _218_.ZN a_50196_22805# 0.01551f
C21102 a_12444_1592# VPWR 0.29679f
C21103 _424_.B1 a_51196_21543# 0.01082f
C21104 a_45820_12568# a_45820_12135# 0.05841f
C21105 _319_.ZN a_35716_20072# 0.00199f
C21106 a_59036_12568# a_59484_12568# 0.01288f
C21107 a_49764_12612# a_49740_12135# 0.00172f
C21108 _290_.ZN VPWR 1.16809f
C21109 a_29856_29123# _369_.ZN 0.00941f
C21110 a_59332_29816# ui_in[3] 0.00226f
C21111 a_47076_31048# vgaringosc.workerclkbuff_notouch_.I 0.00645f
C21112 _256_.A2 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN 0.03159f
C21113 _359_.B a_32848_29123# 0.0143f
C21114 a_47524_11044# a_47164_11000# 0.08707f
C21115 a_33948_19975# VPWR 0.34938f
C21116 a_4852_9096# VPWR 0.22733f
C21117 a_65220_5960# VPWR 0.20921f
C21118 a_35628_18407# VPWR 0.32798f
C21119 _452_.CLK a_31820_21976# 0.0021f
C21120 a_63764_23588# a_63404_23544# 0.0869f
C21121 a_34084_28776# a_34700_28776# 0.00817f
C21122 _293_.A2 a_39300_29480# 0.00501f
C21123 _242_.Z a_57168_26724# 0.00399f
C21124 a_59732_10664# a_60180_10664# 0.01328f
C21125 a_29020_1159# a_29468_1159# 0.0131f
C21126 a_21764_24776# a_21852_23111# 0.00151f
C21127 a_932_1636# a_1020_1592# 0.28563f
C21128 _397_.A1 _390_.ZN 0.02775f
C21129 a_3260_26680# a_3260_26247# 0.05841f
C21130 a_31732_22020# VPWR 0.20595f
C21131 _251_.A1 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.009f
C21132 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I 0.00855f
C21133 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I 0.18273f
C21134 _304_.ZN a_44038_21236# 0.00523f
C21135 a_2724_12612# VPWR 0.20782f
C21136 a_31396_21640# a_31844_21640# 0.01328f
C21137 a_49404_2727# VPWR 0.31651f
C21138 a_37396_29860# VPWR 0.01455f
C21139 a_16140_26247# a_16052_26344# 0.28563f
C21140 a_32964_15368# a_33412_15368# 0.01328f
C21141 _427_.ZN a_56180_22137# 0.00248f
C21142 a_17956_29860# VPWR 0.21041f
C21143 _359_.B a_34348_27208# 0.00202f
C21144 a_36772_23208# a_36148_21976# 0.00131f
C21145 _395_.A2 a_51016_25940# 0.00282f
C21146 a_50636_10567# VPWR 0.33727f
C21147 a_35068_15271# a_34980_15368# 0.28563f
C21148 a_24428_21976# a_24540_21543# 0.02634f
C21149 a_52228_27912# VPWR 0.20645f
C21150 a_28372_22020# a_28348_21543# 0.00172f
C21151 _249_.A2 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.00637f
C21152 a_3172_23208# VPWR 0.20993f
C21153 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN a_65308_19975# 0.00128f
C21154 _304_.B _267_.A2 0.0246f
C21155 a_36412_15271# a_36860_15271# 0.0131f
C21156 _350_.A1 a_35292_30951# 0.01418f
C21157 a_932_28292# a_1020_28248# 0.28563f
C21158 a_1828_22020# a_1468_21976# 0.08717f
C21159 a_3620_22020# a_4068_22020# 0.01328f
C21160 a_48956_2727# a_48868_2824# 0.28563f
C21161 a_65220_17316# a_64860_17272# 0.08717f
C21162 a_33483_29535# a_33768_29535# 0.00277f
C21163 a_56572_23111# a_56484_23208# 0.28563f
C21164 a_62196_26724# _245_.I1 0.00196f
C21165 a_29828_1256# a_30276_1256# 0.01328f
C21166 a_21068_23544# a_21516_23544# 0.01288f
C21167 a_64860_7431# a_65308_7431# 0.0131f
C21168 a_65756_5863# a_66204_5863# 0.0131f
C21169 a_66652_4295# a_67100_4295# 0.0131f
C21170 a_9084_2727# a_9532_2727# 0.0131f
C21171 a_58924_13703# a_59372_13703# 0.01288f
C21172 a_49404_14136# a_49316_12612# 0.00151f
C21173 _393_.ZN a_46580_28292# 0.0089f
C21174 a_40916_16936# a_41116_15271# 0.00119f
C21175 a_66452_18504# a_66564_17316# 0.02666f
C21176 a_60964_26344# a_61412_26344# 0.01328f
C21177 _398_.C _399_.ZN 1.82422f
C21178 a_31708_16839# a_32068_16936# 0.08717f
C21179 a_54432_31128# _268_.A1 0.02187f
C21180 _419_.A4 a_47636_23588# 0.00222f
C21181 a_26244_1636# VPWR 0.21372f
C21182 a_1380_10664# a_1380_9476# 0.05841f
C21183 _419_.Z a_50748_20408# 0.00763f
C21184 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN 0.05006f
C21185 a_13004_30951# a_13452_30951# 0.01222f
C21186 _371_.A1 _336_.A1 0.02044f
C21187 a_66340_12612# a_66428_12568# 0.28563f
C21188 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I a_58700_16839# 0.00101f
C21189 a_4156_23544# a_4156_23111# 0.05841f
C21190 _294_.A2 _288_.ZN 0.45226f
C21191 _245_.Z a_61836_26680# 0.00791f
C21192 _388_.B a_43788_29167# 0.00187f
C21193 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN 0.00225f
C21194 a_63428_18504# a_63876_18504# 0.01328f
C21195 a_2276_15368# a_2276_14180# 0.05841f
C21196 a_54020_11044# a_54468_11044# 0.01328f
C21197 a_45172_16936# a_45620_16936# 0.01328f
C21198 a_43716_1636# a_43804_1592# 0.28563f
C21199 _417_.Z a_49068_20408# 0.02434f
C21200 _424_.B1 a_52228_19368# 0.46773f
C21201 _407_.A1 _395_.A2 0.00545f
C21202 a_45820_18840# a_45820_18407# 0.05841f
C21203 hold2.I a_43126_24119# 0.00106f
C21204 _251_.A1 a_58364_25112# 0.02327f
C21205 _272_.A2 a_58116_30344# 0.58611f
C21206 a_43736_25896# a_44744_26355# 0.02307f
C21207 _470_.Q a_47172_27912# 0.00162f
C21208 a_33188_2824# a_33188_1636# 0.05841f
C21209 a_18096_27165# a_19524_26344# 0.00172f
C21210 _258_.ZN vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I 0.70603f
C21211 a_33492_25273# VPWR 0.00258f
C21212 a_16500_20452# VPWR 0.20348f
C21213 _349_.A4 a_25124_28776# 1.31484f
C21214 a_51644_12568# VPWR 0.31547f
C21215 _452_.Q a_42630_21236# 0.00236f
C21216 _359_.B a_44795_29535# 0.02978f
C21217 a_22352_25987# a_23420_26247# 0.00506f
C21218 a_9892_2824# a_10340_2824# 0.01328f
C21219 uo_out[0] uo_out[1] 0.06751f
C21220 a_7516_29383# a_7876_29480# 0.08717f
C21221 a_57020_23111# vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN 0.01053f
C21222 a_4156_28248# a_4156_27815# 0.05841f
C21223 a_4852_10664# VPWR 0.22733f
C21224 a_23084_21976# a_23108_21640# 0.00172f
C21225 a_46044_15271# a_46404_15368# 0.08717f
C21226 a_36548_26724# a_36996_26724# 0.01328f
C21227 _312_.ZN VPWR 0.65591f
C21228 a_35140_26680# a_35552_27216# 0.00705f
C21229 _267_.A2 VPWR 1.24734f
C21230 _260_.A1 a_40668_20408# 0.00142f
C21231 a_16140_28248# a_16588_28248# 0.012f
C21232 a_38971_18559# VPWR 0.36806f
C21233 a_15604_22020# a_15244_21976# 0.08707f
C21234 a_63516_15704# VPWR 0.29679f
C21235 a_59932_2727# a_60292_2824# 0.08717f
C21236 _336_.A1 a_30476_25112# 0.00209f
C21237 a_44252_30951# a_44612_31048# 0.08717f
C21238 a_22620_27599# VPWR 0.39801f
C21239 a_63428_15368# a_63876_15368# 0.01328f
C21240 a_53212_29816# VPWR 0.82049f
C21241 _474_.CLK _397_.A2 1.00619f
C21242 a_53572_27912# _412_.ZN 0.00192f
C21243 _433_.ZN _441_.A3 0.04687f
C21244 a_57044_18504# a_57492_18504# 0.01328f
C21245 _267_.A2 a_59332_29816# 0.16549f
C21246 a_14148_1256# VPWR 0.20348f
C21247 a_19724_25112# a_20172_25112# 0.01288f
C21248 a_3708_7864# VPWR 0.33374f
C21249 a_64324_4772# VPWR 0.22383f
C21250 _448_.Q _324_.B 0.01371f
C21251 a_33500_18840# a_33500_18407# 0.05841f
C21252 a_56012_13703# a_55924_13800# 0.28563f
C21253 _417_.Z a_48776_20204# 0.03745f
C21254 _475_.D a_45696_20072# 0.0028f
C21255 a_52116_16936# a_52092_15271# 0.00134f
C21256 a_4828_29383# VPWR 0.33352f
C21257 _360_.ZN a_33396_26344# 0.01509f
C21258 a_53704_23219# a_54088_22895# 1.16391f
C21259 _351_.A2 a_25796_27912# 0.00653f
C21260 _330_.A1 a_40464_27165# 0.01628f
C21261 _250_.C a_61940_29076# 0.40764f
C21262 a_43020_16839# a_42932_16936# 0.28563f
C21263 _417_.A2 a_51240_23340# 0.24404f
C21264 a_1468_1159# a_1828_1256# 0.08717f
C21265 a_4852_16936# VPWR 0.22733f
C21266 a_32380_1592# VPWR 0.30141f
C21267 a_45820_12135# a_46268_12135# 0.0131f
C21268 a_43044_27912# VPWR 0.2117f
C21269 a_2812_1592# a_3260_1592# 0.01288f
C21270 a_6756_1636# a_6844_1592# 0.28563f
C21271 a_1828_29860# a_1468_29816# 0.08707f
C21272 _424_.B1 a_50196_21640# 0.00361f
C21273 _241_.I0 a_57244_27815# 0.00731f
C21274 _319_.A2 a_36612_20072# 0.00208f
C21275 a_4964_17316# a_5052_17272# 0.28563f
C21276 _459_.CLK a_31820_25112# 0.04795f
C21277 _470_.Q _412_.A1 0.01507f
C21278 vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I a_66676_20452# 0.00197f
C21279 a_22884_1636# a_22748_1159# 0.00168f
C21280 a_18940_1592# a_18940_1159# 0.05841f
C21281 a_63764_12232# a_63852_10567# 0.00151f
C21282 _424_.A2 _284_.B 0.13064f
C21283 _402_.ZN a_46356_24072# 0.05691f
C21284 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I 0.00296f
C21285 a_46268_18407# a_46628_18504# 0.08717f
C21286 a_51420_1159# a_51868_1159# 0.0131f
C21287 _474_.CLK a_55140_27912# 0.00168f
C21288 a_64772_18884# a_64860_18840# 0.28563f
C21289 a_64412_18407# VPWR 0.29986f
C21290 _256_.A2 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I 0.00779f
C21291 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I _249_.A2 0.02493f
C21292 a_3260_25112# VPWR 0.30487f
C21293 a_57492_18504# a_57492_17316# 0.05841f
C21294 a_27476_20452# VPWR 0.21518f
C21295 a_4940_27815# a_4852_27912# 0.28563f
C21296 a_61029_30644# ui_in[3] 0.00145f
C21297 a_65444_12612# VPWR 0.21306f
C21298 a_3708_15704# a_4156_15704# 0.0131f
C21299 a_21292_30951# _379_.A2 0.00766f
C21300 a_55364_15368# a_55812_15368# 0.01328f
C21301 a_39908_15748# a_39772_15271# 0.00168f
C21302 a_19035_28409# a_19860_27912# 0.0017f
C21303 a_19328_28733# a_19412_27912# 0.00101f
C21304 a_66228_10664# VPWR 0.22591f
C21305 _355_.B a_28679_24776# 0.0282f
C21306 a_65756_8999# a_66116_9096# 0.08717f
C21307 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I 0.0091f
C21308 a_66652_7431# a_67012_7528# 0.08717f
C21309 a_34732_16839# a_34756_15748# 0.0016f
C21310 a_24092_21543# a_24116_20452# 0.0016f
C21311 a_39684_15368# VPWR 0.20348f
C21312 _340_.A2 _459_.CLK 0.09546f
C21313 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I 0.0641f
C21314 a_41996_28777# a_42340_28409# 0.00275f
C21315 a_21964_21976# a_22548_22020# 0.01675f
C21316 _268_.A2 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I 0.00279f
C21317 a_4964_14180# a_5052_14136# 0.28563f
C21318 a_40108_16839# a_40556_16839# 0.01288f
C21319 _395_.A1 _399_.A1 0.50802f
C21320 a_43132_15271# VPWR 0.30179f
C21321 _230_.I ui_in[2] 0.05347f
C21322 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN 0.29243f
C21323 a_67100_17272# VPWR 0.31547f
C21324 _359_.B a_34844_24679# 0.00244f
C21325 a_52228_1256# a_52676_1256# 0.01328f
C21326 a_36548_1256# VPWR 0.20348f
C21327 _459_.Q _459_.CLK 0.26253f
C21328 a_52788_13800# a_53236_13800# 0.01328f
C21329 a_31484_2727# a_31932_2727# 0.0131f
C21330 a_66764_13703# a_67124_13800# 0.08717f
C21331 a_50636_13703# a_50660_12612# 0.0016f
C21332 a_35740_17272# a_35628_16839# 0.02634f
C21333 a_57492_17316# a_57940_17316# 0.01328f
C21334 a_41488_24072# _305_.A2 0.3859f
C21335 a_2724_17316# VPWR 0.20782f
C21336 a_53548_16839# a_53908_16936# 0.08674f
C21337 _229_.I _243_.ZN 0.01527f
C21338 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I 0.00163f
C21339 _268_.A1 _274_.A1 0.08462f
C21340 a_3260_12135# a_3172_12232# 0.28563f
C21341 a_46044_1592# VPWR 0.29679f
C21342 _402_.A1 a_47802_26724# 0.0029f
C21343 a_12892_1159# a_12804_1256# 0.28563f
C21344 a_52988_1592# a_53124_1256# 0.00168f
C21345 a_51668_16936# VPWR 0.2061f
C21346 a_28012_23544# a_27900_23111# 0.02634f
C21347 a_10116_1636# a_9756_1592# 0.08707f
C21348 a_8188_29816# a_8772_29860# 0.01675f
C21349 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN 0.02665f
C21350 _251_.A1 _270_.A2 0.0236f
C21351 _424_.A2 _474_.D 0.47527f
C21352 a_34756_17316# a_34844_17272# 0.28563f
C21353 a_30812_17272# a_31260_17272# 0.01288f
C21354 _416_.A1 a_40580_26344# 0.00558f
C21355 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I 0.01518f
C21356 _416_.ZN a_47028_18884# 0.00621f
C21357 a_64548_11044# a_64188_11000# 0.08707f
C21358 a_16612_2824# VPWR 0.20348f
C21359 a_53436_1592# a_53884_1592# 0.01288f
C21360 a_62196_26724# a_62284_26680# 0.28563f
C21361 _448_.D a_36060_19369# 0.21954f
C21362 a_43126_24119# VPWR 0.58785f
C21363 a_19164_23111# a_19612_23111# 0.01288f
C21364 a_1468_24679# a_1828_24776# 0.08717f
C21365 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN 0.00209f
C21366 _459_.CLK a_22352_25987# 0.00706f
C21367 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I a_65756_26247# 0.00201f
C21368 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN a_64188_27815# 0.04158f
C21369 _337_.A3 _352_.ZN 0.01066f
C21370 a_2724_14180# VPWR 0.20782f
C21371 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN a_60180_14180# 0.00189f
C21372 _474_.CLK a_54356_23588# 0.00271f
C21373 _363_.Z _460_.Q 1.0846f
C21374 _250_.B vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.00194f
C21375 a_25936_25597# VPWR 0.51865f
C21376 _459_.CLK a_16140_28248# 0.00177f
C21377 a_20672_30301# a_21540_28292# 0.00142f
C21378 VPWR uio_out[5] 1.31828f
C21379 _264_.B _452_.Q 0.00673f
C21380 _261_.ZN _441_.A3 0.5161f
C21381 _260_.A1 a_40780_21543# 0.0087f
C21382 a_52428_12135# VPWR 0.31389f
C21383 a_1380_29480# VPWR 0.20348f
C21384 a_36100_15748# a_35740_15704# 0.08707f
C21385 _459_.CLK _461_.D 0.01324f
C21386 a_32292_2824# a_32740_2824# 0.01328f
C21387 _251_.A1 clk 0.17643f
C21388 a_19860_27912# uio_out[7] 0.00252f
C21389 a_14796_24679# VPWR 0.30073f
C21390 a_22660_21640# a_22772_20452# 0.02666f
C21391 _452_.CLK a_44752_18147# 0.05698f
C21392 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I 0.14093f
C21393 a_35204_15748# VPWR 0.21603f
C21394 _402_.ZN a_46620_22504# 0.00932f
C21395 _355_.C a_30240_24776# 0.00814f
C21396 a_28112_27912# VPWR 0.0139f
C21397 a_2276_9476# a_1916_9432# 0.08717f
C21398 a_4068_9476# a_4516_9476# 0.01328f
C21399 _228_.ZN a_58116_30344# 0.41223f
C21400 _218_.ZN a_50196_21640# 0.00803f
C21401 a_29268_22020# a_28908_21976# 0.08707f
C21402 a_50644_21640# VPWR 0.00753f
C21403 _474_.CLK _330_.A1 0.09879f
C21404 a_45372_14136# a_45820_14136# 0.01288f
C21405 a_49316_14180# a_49404_14136# 0.28563f
C21406 _452_.Q _332_.Z 0.00403f
C21407 a_58028_18840# a_58476_18840# 0.01255f
C21408 _452_.CLK a_39324_17272# 0.00613f
C21409 a_46604_16839# VPWR 0.31556f
C21410 _397_.A2 _398_.C 0.05917f
C21411 a_58948_1256# VPWR 0.20348f
C21412 a_67324_14136# a_67236_12612# 0.00151f
C21413 a_57580_13703# a_57604_12612# 0.0016f
C21414 a_47524_13800# a_47524_12612# 0.05841f
C21415 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_59708_23111# 0.02694f
C21416 _296_.ZN uo_out[2] 0.01592f
C21417 _237_.A1 a_59744_30352# 0.0014f
C21418 a_62420_10664# a_62396_9432# 0.0016f
C21419 a_37084_17272# VPWR 0.31547f
C21420 a_23868_1159# a_24228_1256# 0.08717f
C21421 a_67660_12135# a_68108_12135# 0.0131f
C21422 a_53772_12135# a_54132_12232# 0.08707f
C21423 a_59844_1636# VPWR 0.20348f
C21424 a_17060_29480# _467_.D 0.01756f
C21425 a_16612_1636# a_17060_1636# 0.01328f
C21426 a_15492_29860# a_15132_29816# 0.08707f
C21427 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN VPWR 0.74635f
C21428 a_40644_17272# a_41432_17801# 0.02112f
C21429 _459_.Q _371_.A3 0.31421f
C21430 _336_.A2 a_27116_23544# 0.00613f
C21431 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_59372_14136# 0.00861f
C21432 _304_.B a_44282_24164# 0.00139f
C21433 a_39012_2824# VPWR 0.22423f
C21434 a_52639_30644# input9.Z 0.21367f
C21435 _474_.CLK a_54432_31128# 0.05511f
C21436 a_60740_1636# a_60380_1592# 0.08707f
C21437 _304_.B vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.04381f
C21438 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.21353f
C21439 _459_.CLK a_20308_27912# 0.00277f
C21440 a_3620_24776# a_4068_24776# 0.01328f
C21441 a_17932_23111# a_17844_23208# 0.28563f
C21442 a_21852_24679# a_21764_24776# 0.28563f
C21443 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN 0.02499f
C21444 _330_.A1 a_34308_21640# 0.0069f
C21445 a_45732_9476# VPWR 0.20348f
C21446 a_45036_28248# _403_.ZN 0.00118f
C21447 a_51644_14136# VPWR 0.31547f
C21448 _316_.A3 _319_.A3 0.03468f
C21449 _334_.A1 uo_out[1] 0.01143f
C21450 _388_.B a_45416_29885# 0.01714f
C21451 a_33948_18407# a_34644_18504# 0.01227f
C21452 a_45012_29816# a_45360_29977# 0.00277f
C21453 _251_.A1 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I 1.26433f
C21454 a_3172_18504# a_3620_18504# 0.01328f
C21455 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN clk 0.02061f
C21456 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I 0.00194f
C21457 a_42596_15748# a_43044_15748# 0.01328f
C21458 a_46180_12232# VPWR 0.20348f
C21459 a_61836_23544# vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN 0.00241f
C21460 a_39012_15748# a_39100_15704# 0.28563f
C21461 _340_.A2 uo_out[7] 0.00618f
C21462 _245_.Z a_62396_26247# 0.0066f
C21463 a_19524_24776# VPWR 0.23492f
C21464 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN a_54892_16839# 0.03994f
C21465 a_30052_21640# a_29940_20452# 0.02666f
C21466 a_3708_2727# a_4068_2824# 0.08717f
C21467 a_30812_19975# a_30724_20072# 0.28563f
C21468 a_41340_15704# VPWR 0.33277f
C21469 _290_.ZN a_35292_30951# 0.0042f
C21470 _459_.Q uo_out[7] 0.04762f
C21471 a_48420_9476# a_48508_9432# 0.28563f
C21472 a_62620_19975# VPWR 0.32666f
C21473 a_52540_14136# a_53212_14136# 0.00544f
C21474 _452_.CLK a_36636_26247# 0.00766f
C21475 _444_.D _304_.A1 0.00587f
C21476 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN a_61724_19975# 0.00196f
C21477 _265_.ZN _330_.A1 0.04345f
C21478 _260_.A2 a_42168_22504# 0.02076f
C21479 a_53660_2727# a_54332_2727# 0.00544f
C21480 a_54580_13800# a_54468_12612# 0.02666f
C21481 a_2364_12568# a_2812_12568# 0.0131f
C21482 a_4964_12612# a_4604_12568# 0.08674f
C21483 a_34939_23705# _304_.A1 0.00484f
C21484 _397_.A2 _393_.A3 0.69138f
C21485 _251_.A1 _241_.Z 0.03327f
C21486 a_59955_30600# a_60909_30600# 0.00337f
C21487 _398_.C a_48308_23588# 0.04334f
C21488 a_49180_17272# VPWR 0.318f
C21489 a_1916_1159# VPWR 0.297f
C21490 a_35292_1159# a_35204_1256# 0.28563f
C21491 a_23780_1636# a_23420_1592# 0.08663f
C21492 a_64972_12135# a_64884_12232# 0.28563f
C21493 a_1828_5960# a_1828_4772# 0.05841f
C21494 a_2724_4392# a_2724_3204# 0.05841f
C21495 a_29692_21543# VPWR 0.31389f
C21496 a_23556_29860# _459_.CLK 0.01814f
C21497 a_46852_17316# a_46940_17272# 0.28563f
C21498 _311_.A2 a_37408_23208# 0.00164f
C21499 _424_.A2 _474_.Q 0.10401f
C21500 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_62868_23208# 0.00192f
C21501 _433_.ZN _226_.ZN 0.59449f
C21502 a_50436_17316# a_50884_17316# 0.01328f
C21503 _460_.D a_33076_24776# 0.00219f
C21504 _478_.D a_53300_23047# 0.02548f
C21505 a_54668_10567# a_55116_10567# 0.01288f
C21506 a_1020_10567# a_1380_10664# 0.08717f
C21507 a_65444_1636# a_65084_1592# 0.08717f
C21508 a_67236_1636# a_67684_1636# 0.01328f
C21509 a_61188_2824# VPWR 0.20968f
C21510 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN VPWR 0.44382f
C21511 _294_.ZN uo_out[6] 0.42417f
C21512 _461_.D uo_out[7] 0.00336f
C21513 a_16500_23208# a_16948_23208# 0.01328f
C21514 a_28796_23111# a_29156_23208# 0.08707f
C21515 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN 0.01444f
C21516 a_56708_9476# VPWR 0.23226f
C21517 a_25124_2824# a_25212_1159# 0.0027f
C21518 a_23196_21543# a_23644_21543# 0.01288f
C21519 a_1916_21543# a_1828_21640# 0.28563f
C21520 a_67236_14180# VPWR 0.20348f
C21521 a_60276_29032# a_60656_29612# 0.00217f
C21522 _398_.C a_54356_23588# 0.0117f
C21523 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I a_56596_17316# 0.00167f
C21524 a_43296_28733# a_43132_27815# 0.00119f
C21525 _230_.I a_61948_27815# 0.00175f
C21526 _337_.A3 a_26746_26344# 0.00103f
C21527 a_68020_12232# VPWR 0.21406f
C21528 _433_.ZN _300_.ZN 0.11587f
C21529 a_45920_20523# VPWR 1.10606f
C21530 a_37980_2727# a_38116_1636# 0.00154f
C21531 a_54692_2824# a_55140_2824# 0.01328f
C21532 a_61724_19975# a_62084_20072# 0.08717f
C21533 _365_.ZN _462_.D 0.92582f
C21534 _255_.ZN ui_in[4] 0.01314f
C21535 a_22548_29480# _454_.D 0.00141f
C21536 _460_.Q a_35660_27508# 0.00521f
C21537 _303_.ZN a_40244_21640# 0.00247f
C21538 a_36516_24831# VPWR 0.00246f
C21539 _302_.Z _304_.ZN 1.77121f
C21540 a_1468_18840# VPWR 0.29679f
C21541 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I 0.00682f
C21542 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I a_63404_20408# 0.01978f
C21543 a_15132_2727# a_15044_2824# 0.28563f
C21544 a_55140_15748# VPWR 0.21152f
C21545 _251_.ZN vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN 0.00914f
C21546 _264_.B a_40357_24776# 0.0238f
C21547 _251_.A1 a_58948_26344# 0.02053f
C21548 a_53796_9476# a_54244_9476# 0.01328f
C21549 a_26916_31048# uio_out[1] 0.01885f
C21550 a_63316_23588# VPWR 0.19301f
C21551 a_65756_23111# clk 0.00228f
C21552 a_50660_14180# a_50636_13703# 0.00172f
C21553 a_46716_14136# a_46716_13703# 0.05841f
C21554 a_3172_20452# a_3260_20408# 0.28563f
C21555 a_60964_14180# a_61412_14180# 0.01328f
C21556 a_30388_28776# a_34084_28776# 0.0245f
C21557 _294_.A2 a_34586_27912# 0.01039f
C21558 _256_.A2 VPWR 0.88648f
C21559 _304_.A1 a_34715_22137# 0.00916f
C21560 _230_.I a_61297_30300# 0.52127f
C21561 a_61524_13800# a_61412_12612# 0.02666f
C21562 a_49316_12612# a_48956_12568# 0.08707f
C21563 _294_.ZN uo_out[5] 0.00146f
C21564 a_15604_24776# a_15604_23588# 0.05841f
C21565 _452_.CLK a_46252_19759# 0.00394f
C21566 a_46044_1159# a_46628_1256# 0.01675f
C21567 a_24316_1159# VPWR 0.32824f
C21568 _452_.Q a_39236_17316# 0.00699f
C21569 a_61524_12232# a_61972_12232# 0.01328f
C21570 a_30276_1636# a_30724_1636# 0.01328f
C21571 a_26692_1636# a_26780_1592# 0.28563f
C21572 a_39772_20408# a_40220_20408# 0.01222f
C21573 _438_.A2 a_39324_26247# 0.00883f
C21574 _436_.B _264_.B 0.14398f
C21575 a_35292_26247# a_35204_26344# 0.28563f
C21576 _256_.A2 a_59332_29816# 0.16728f
C21577 a_26916_21640# VPWR 0.22421f
C21578 a_52848_25987# a_53260_26399# 0.00275f
C21579 _352_.ZN a_27328_25227# 0.00421f
C21580 a_54780_26247# a_54692_26344# 0.28563f
C21581 _416_.A1 _400_.ZN 0.03903f
C21582 a_51980_10567# a_51892_10664# 0.28563f
C21583 _474_.CLK _274_.A1 0.04361f
C21584 a_51108_1636# a_50972_1159# 0.00168f
C21585 _325_.A2 _328_.A2 0.32315f
C21586 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I VPWR 0.91619f
C21587 a_61029_31220# VPWR 0.00437f
C21588 _324_.C a_45696_20072# 0.00173f
C21589 a_65668_23208# VPWR 0.24037f
C21590 a_48060_30951# _397_.A2 0.00156f
C21591 _402_.A1 a_40780_27815# 0.0062f
C21592 a_34396_24679# a_34308_24776# 0.28563f
C21593 a_67548_9432# VPWR 0.32994f
C21594 a_16588_23544# VPWR 0.29679f
C21595 a_66900_20072# a_67348_20072# 0.01328f
C21596 a_21852_21543# a_22212_21640# 0.08707f
C21597 a_4156_2727# VPWR 0.3339f
C21598 _459_.CLK a_27004_27815# 0.02166f
C21599 a_2364_5863# VPWR 0.30029f
C21600 _336_.A2 a_29156_23208# 0.00167f
C21601 a_54220_13703# VPWR 0.31594f
C21602 a_15492_29860# uio_oe[1] 0.00143f
C21603 a_48732_15704# a_49180_15704# 0.01288f
C21604 a_52676_15748# a_52764_15704# 0.28563f
C21605 a_49404_11000# VPWR 0.32097f
C21606 a_45696_20072# _416_.ZN 0.30293f
C21607 a_54892_23544# a_55340_23544# 0.0131f
C21608 a_4964_26724# VPWR 0.21167f
C21609 a_59172_23588# _231_.I 0.00549f
C21610 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I 0.80012f
C21611 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I 0.06734f
C21612 a_48956_30951# vgaringosc.workerclkbuff_notouch_.I 0.00613f
C21613 a_16948_26344# VPWR 0.20348f
C21614 a_26108_2727# a_26468_2824# 0.08717f
C21615 _245_.Z a_61860_26344# 0.05199f
C21616 a_23084_30951# uio_out[3] 0.00996f
C21617 a_64748_23544# clk 0.00613f
C21618 _350_.A2 _362_.ZN 0.02937f
C21619 a_59396_9476# a_59484_9432# 0.28563f
C21620 a_4604_28248# VPWR 0.33016f
C21621 a_39884_27815# _330_.A1 0.00839f
C21622 a_61052_26247# a_61412_26344# 0.0869f
C21623 _272_.A2 _274_.A2 0.38675f
C21624 a_1380_4772# a_1468_4728# 0.28563f
C21625 a_57604_14180# a_57580_13703# 0.00172f
C21626 a_54108_14136# a_54220_13703# 0.02634f
C21627 a_2276_3204# a_2364_3160# 0.28563f
C21628 _300_.A2 _325_.A2 0.00216f
C21629 a_17036_20408# a_17484_20408# 0.0131f
C21630 a_56148_23588# a_55788_23544# 0.08717f
C21631 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I a_61388_15704# 0.00131f
C21632 a_55812_12612# a_56260_12612# 0.01328f
C21633 a_5860_1636# VPWR 0.20884f
C21634 _393_.A3 _330_.A1 0.00952f
C21635 _459_.CLK a_16500_25156# 0.00249f
C21636 a_30778_31048# uo_out[6] 0.00172f
C21637 a_47948_23111# _475_.Q 0.00223f
C21638 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN 0.00152f
C21639 a_22660_24776# a_22548_23588# 0.02666f
C21640 clkbuf_1_0__f_clk.I _397_.Z 0.00178f
C21641 a_46716_1159# VPWR 0.33352f
C21642 a_57468_1159# a_57380_1256# 0.28563f
C21643 a_64324_18884# VPWR 0.20554f
C21644 a_2724_11044# a_2812_11000# 0.28563f
C21645 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _275_.ZN 0.47922f
C21646 _244_.Z a_60740_26724# 0.00995f
C21647 _441_.ZN _325_.A1 0.00237f
C21648 a_46476_20937# a_46820_20569# 0.00275f
C21649 a_49068_20408# a_49652_20936# 0.00629f
C21650 _260_.A1 _434_.ZN 0.00269f
C21651 _261_.ZN _300_.ZN 0.11577f
C21652 _452_.CLK a_31372_23544# 0.00176f
C21653 _284_.B hold1.Z 0.0425f
C21654 _241_.Z a_58020_27508# 0.36509f
C21655 a_62508_10567# a_62868_10664# 0.08707f
C21656 a_48420_10664# a_49204_10664# 0.00276f
C21657 _274_.ZN uio_in[0] 0.04462f
C21658 a_17596_1159# a_18044_1159# 0.0131f
C21659 _459_.CLK a_43232_29480# 0.00279f
C21660 a_18852_2824# a_18852_1636# 0.05841f
C21661 a_56596_23588# a_57044_23588# 0.01328f
C21662 _459_.CLK a_27460_28776# 0.00216f
C21663 a_53572_21640# a_52452_21236# 0.07607f
C21664 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I _241_.I0 0.00371f
C21665 a_17484_21976# VPWR 0.29719f
C21666 a_43214_21812# VPWR 0.00468f
C21667 a_31284_23588# VPWR 0.20417f
C21668 _350_.A1 a_32240_31048# 0.0068f
C21669 a_20420_21640# a_20868_21640# 0.01328f
C21670 a_32828_21543# a_32740_21640# 0.28563f
C21671 a_26556_2727# VPWR 0.31932f
C21672 a_54692_18884# vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN 0.00315f
C21673 a_47972_13800# VPWR 0.20348f
C21674 a_47524_2824# a_47612_1159# 0.0027f
C21675 a_63964_15271# a_64412_15271# 0.0131f
C21676 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I 0.00427f
C21677 a_3708_29816# VPWR 0.33374f
C21678 a_63204_11044# VPWR 0.20595f
C21679 _268_.A1 a_52292_29480# 0.00254f
C21680 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN _274_.A2 0.0386f
C21681 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN clk 0.18748f
C21682 a_5388_23111# VPWR 0.35526f
C21683 _284_.B a_45396_25156# 0.00158f
C21684 a_45088_29123# a_44948_28292# 0.01115f
C21685 hold1.Z a_43245_24373# 0.00352f
C21686 a_14708_27912# VPWR 0.22176f
C21687 _260_.ZN a_43126_24119# 0.07579f
C21688 a_67548_15704# a_67996_15704# 0.01222f
C21689 a_27004_27815# _371_.A3 0.01308f
C21690 a_62172_17272# a_62084_15748# 0.00151f
C21691 _419_.A4 _282_.ZN 0.34718f
C21692 a_64748_23111# a_64660_23208# 0.28563f
C21693 a_37532_2727# a_37444_2824# 0.28563f
C21694 a_64772_9476# a_65220_9476# 0.01328f
C21695 a_64772_7908# a_64860_7864# 0.28563f
C21696 a_66564_7908# a_67012_7908# 0.01328f
C21697 a_17844_23588# a_18292_23588# 0.01328f
C21698 a_18404_1256# a_18852_1256# 0.01328f
C21699 a_64412_4728# a_64860_4728# 0.0131f
C21700 a_66564_4772# a_66652_4728# 0.28563f
C21701 a_4964_6340# a_4940_5863# 0.00172f
C21702 a_67460_6340# a_67908_6340# 0.01328f
C21703 a_65668_6340# a_65756_6296# 0.28563f
C21704 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I a_61388_16839# 0.00631f
C21705 a_47612_13703# a_48060_13703# 0.0131f
C21706 a_65308_3160# a_65756_3160# 0.0131f
C21707 a_67460_3204# a_67548_3160# 0.28563f
C21708 a_65444_14180# a_65420_13703# 0.00172f
C21709 _312_.ZN _311_.Z 0.4731f
C21710 _402_.A1 _397_.A4 0.59986f
C21711 a_4852_16936# a_4940_15271# 0.00151f
C21712 _470_.Q _381_.Z 0.14899f
C21713 a_22772_20452# a_22860_20408# 0.28563f
C21714 _459_.Q a_31820_25112# 0.02166f
C21715 a_59172_22020# VPWR 0.14845f
C21716 a_9084_29383# a_9532_29383# 0.0131f
C21717 _323_.A3 VPWR 0.53719f
C21718 a_11548_30951# a_11460_31048# 0.28563f
C21719 _457_.D a_25436_24679# 0.00525f
C21720 a_54824_22045# vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN 0.00634f
C21721 a_63068_17272# a_63180_16839# 0.02634f
C21722 _424_.B1 a_51332_24072# 0.10202f
C21723 a_11996_1592# VPWR 0.33603f
C21724 a_65780_13800# a_65868_12135# 0.00151f
C21725 a_31708_1592# a_31844_1256# 0.00168f
C21726 _319_.ZN a_35492_20072# 0.00661f
C21727 a_62060_20408# a_62172_19975# 0.02634f
C21728 _304_.A1 _301_.Z 0.00753f
C21729 a_46628_31048# vgaringosc.workerclkbuff_notouch_.I 0.00648f
C21730 _359_.B a_31920_29480# 0.02104f
C21731 a_30240_24776# a_30836_23588# 0.0111f
C21732 a_4068_9096# VPWR 0.22146f
C21733 a_33500_19975# VPWR 0.3346f
C21734 a_64772_5960# VPWR 0.20727f
C21735 _441_.A3 a_40316_23233# 0.01528f
C21736 a_63316_23588# a_63404_23544# 0.28563f
C21737 a_50660_11044# a_51108_11044# 0.01328f
C21738 a_47076_11044# a_47164_11000# 0.28563f
C21739 a_33860_16936# a_34644_16936# 0.00276f
C21740 a_36412_1592# a_36860_1592# 0.01288f
C21741 a_35180_18407# VPWR 0.33205f
C21742 a_34084_28776# a_34292_28776# 0.00733f
C21743 a_60492_28248# a_60940_28248# 0.01222f
C21744 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN 0.7916f
C21745 _330_.A1 _327_.Z 0.25212f
C21746 a_31284_22020# VPWR 0.20595f
C21747 a_45148_30951# a_45596_30951# 0.0131f
C21748 a_37067_19001# a_37312_19369# 0.00232f
C21749 _304_.ZN a_43814_21236# 0.02253f
C21750 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN a_63721_28776# 0.00123f
C21751 _355_.B _336_.Z 0.13104f
C21752 a_36948_29860# VPWR 0.01438f
C21753 a_48956_2727# VPWR 0.31477f
C21754 _474_.D a_49988_21236# 0.42658f
C21755 a_2276_12612# VPWR 0.20634f
C21756 a_1380_26344# a_1828_26344# 0.01328f
C21757 a_15692_26247# a_16052_26344# 0.08717f
C21758 _350_.A2 _287_.A2 0.1205f
C21759 a_17508_29860# VPWR 0.20851f
C21760 a_50188_10567# VPWR 0.32969f
C21761 a_34620_15271# a_34980_15368# 0.08717f
C21762 VPWR uio_oe[5] 0.27806f
C21763 a_34404_31048# uo_out[5] 0.00223f
C21764 a_2724_23208# VPWR 0.20782f
C21765 a_25012_31048# uio_out[3] 0.00296f
C21766 a_2724_28292# a_3172_28292# 0.01328f
C21767 a_1380_22020# a_1468_21976# 0.28563f
C21768 a_48508_2727# a_48868_2824# 0.08717f
C21769 _272_.A2 a_58340_29860# 0.01547f
C21770 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN VPWR 0.75226f
C21771 a_64772_17316# a_64860_17272# 0.28563f
C21772 a_3172_16936# a_3172_15748# 0.05841f
C21773 _474_.CLK _393_.A1 0.01901f
C21774 a_53704_23219# a_54624_22895# 0.00306f
C21775 a_56124_23111# a_56484_23208# 0.08674f
C21776 a_1020_8999# a_932_9096# 0.28563f
C21777 a_16500_25156# a_16948_25156# 0.01328f
C21778 a_5388_13703# a_5300_13800# 0.28563f
C21779 _334_.A1 _362_.ZN 0.00791f
C21780 a_28012_20408# a_28460_20408# 0.0131f
C21781 a_55700_24776# a_55700_23588# 0.05841f
C21782 _419_.A4 a_47412_23588# 0.00103f
C21783 _424_.A2 _427_.A2 0.21543f
C21784 a_31708_16839# a_31620_16936# 0.28563f
C21785 _419_.Z a_50300_20408# 0.00435f
C21786 a_25796_1636# VPWR 0.21193f
C21787 _424_.A2 a_51196_21543# 0.00931f
C21788 _379_.A2 uio_out[6] 0.39916f
C21789 a_62396_12568# a_62844_12568# 0.01288f
C21790 a_66340_12612# a_65980_12568# 0.08707f
C21791 _407_.ZN a_52228_27912# 0.0544f
C21792 _388_.B a_44160_29123# 0.01271f
C21793 a_52788_12232# a_52876_10567# 0.0027f
C21794 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I a_67212_20408# 0.00275f
C21795 a_43716_1636# a_43356_1592# 0.08707f
C21796 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN 0.03097f
C21797 a_39996_1159# a_40444_1159# 0.0131f
C21798 _373_.ZN VPWR 0.42806f
C21799 _258_.ZN a_56484_29480# 0.00361f
C21800 a_56572_29383# vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I 0.03367f
C21801 a_18096_27165# a_19076_26344# 0.00172f
C21802 _421_.A1 _416_.A3 0.27965f
C21803 a_16052_20452# VPWR 0.20348f
C21804 a_43232_29480# _480_.Q 0.30513f
C21805 a_51196_12568# VPWR 0.31547f
C21806 a_64436_16936# a_64884_16936# 0.01328f
C21807 _359_.B a_43788_29167# 0.02889f
C21808 a_7516_29383# a_7428_29480# 0.28563f
C21809 _451_.Q _435_.A3 0.90073f
C21810 _246_.B2 a_60492_28248# 0.01282f
C21811 a_43940_15368# a_44388_15368# 0.01328f
C21812 a_4068_10664# VPWR 0.22146f
C21813 _324_.C _260_.A1 0.0025f
C21814 a_46044_15271# a_45956_15368# 0.28563f
C21815 _316_.ZN a_34396_21543# 0.11028f
C21816 a_33636_23208# VPWR 0.21664f
C21817 a_66204_2727# a_66340_1636# 0.00154f
C21818 a_34308_24776# a_33932_24073# 0.00189f
C21819 a_47388_15271# a_47836_15271# 0.0131f
C21820 _352_.A2 _358_.A2 0.33535f
C21821 _324_.C _428_.Z 0.006f
C21822 _476_.Q a_51912_20452# 0.00319f
C21823 a_37964_18191# VPWR 0.39872f
C21824 a_18740_22020# a_19188_22020# 0.01328f
C21825 a_59932_2727# a_59844_2824# 0.28563f
C21826 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I 0.13732f
C21827 _336_.A1 a_30388_25156# 0.01521f
C21828 a_15156_22020# a_15244_21976# 0.28563f
C21829 a_22992_27555# VPWR 0.18684f
C21830 a_63068_15704# VPWR 0.29679f
C21831 _304_.B _395_.A1 0.5893f
C21832 a_3708_16839# a_4156_16839# 0.0131f
C21833 a_44252_30951# a_44164_31048# 0.28563f
C21834 a_53124_27912# _412_.ZN 0.00167f
C21835 a_36884_16936# a_36996_15748# 0.02666f
C21836 a_25348_23208# a_25436_21543# 0.00151f
C21837 _294_.ZN _460_.Q 0.02096f
C21838 _362_.B uo_out[6] 0.0115f
C21839 a_13700_1256# VPWR 0.20348f
C21840 a_3260_7864# VPWR 0.30487f
C21841 a_25324_23544# a_25772_23544# 0.0131f
C21842 _452_.CLK _330_.A1 3.39929f
C21843 _475_.Q a_48529_22460# 0.59206f
C21844 a_40804_1256# a_41252_1256# 0.01328f
C21845 a_28124_26680# VPWR 0.33273f
C21846 a_5052_4728# VPWR 0.33516f
C21847 _276_.A2 VPWR 0.29986f
C21848 _465_.D VPWR 0.70148f
C21849 a_4156_29383# VPWR 0.3339f
C21850 a_20060_2727# a_20508_2727# 0.0131f
C21851 a_1828_13800# a_2276_13800# 0.01328f
C21852 a_53704_23219# a_54192_22851# 0.8399f
C21853 a_55564_13703# a_55924_13800# 0.08707f
C21854 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN 0.0019f
C21855 a_24900_27912# a_25796_27912# 0.00455f
C21856 a_22188_30951# uio_out[5] 0.00409f
C21857 a_3260_17272# a_3260_16839# 0.05841f
C21858 a_42572_16839# a_42932_16936# 0.08707f
C21859 a_39460_1636# VPWR 0.20968f
C21860 a_58028_10567# a_58052_9476# 0.0016f
C21861 a_4068_16936# VPWR 0.22146f
C21862 a_1468_1159# a_1380_1256# 0.28563f
C21863 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN 0.69671f
C21864 a_6756_1636# a_6396_1592# 0.08707f
C21865 a_42596_27912# VPWR 0.23733f
C21866 a_20172_23544# a_20060_23111# 0.02634f
C21867 a_4964_29860# a_5412_29860# 0.01328f
C21868 a_1380_29860# a_1468_29816# 0.28563f
C21869 a_4964_17316# a_4604_17272# 0.08674f
C21870 _470_.Q a_47173_27208# 0.0096f
C21871 _241_.I0 a_56124_27815# 0.01458f
C21872 a_2364_17272# a_2812_17272# 0.0131f
C21873 _369_.ZN VPWR 0.44034f
C21874 a_56796_11000# a_57244_11000# 0.01288f
C21875 a_50212_1636# a_50660_1636# 0.01328f
C21876 _352_.A2 _355_.ZN 0.38236f
C21877 _441_.B _302_.Z 0.0096f
C21878 a_58164_16936# a_58612_16936# 0.01328f
C21879 _395_.A3 _427_.ZN 0.00145f
C21880 _452_.Q _325_.A2 0.04603f
C21881 a_4068_20072# a_4068_18884# 0.05841f
C21882 _424_.A2 a_52228_19368# 0.37578f
C21883 a_46268_18407# a_46180_18504# 0.28563f
C21884 a_57132_18407# a_57580_18407# 0.012f
C21885 a_47972_18504# a_47948_16839# 0.00131f
C21886 _324_.C _249_.A2 0.07379f
C21887 _421_.B _419_.Z 0.00505f
C21888 _474_.CLK a_53572_27912# 0.0152f
C21889 a_64772_18884# a_64412_18840# 0.08717f
C21890 a_63964_18407# VPWR 0.29679f
C21891 _256_.A2 a_61689_29860# 0.00106f
C21892 a_4156_27815# a_4852_27912# 0.01227f
C21893 a_2812_25112# VPWR 0.30213f
C21894 a_19500_27815# a_19948_27815# 0.01222f
C21895 a_27028_20452# VPWR 0.23583f
C21896 _284_.B clkbuf_1_0__f_clk.I 0.00739f
C21897 _474_.Q a_49988_21236# 0.03684f
C21898 a_64996_12612# VPWR 0.2109f
C21899 a_20868_2824# a_21316_2824# 0.01328f
C21900 _234_.ZN uo_out[1] 0.00334f
C21901 _397_.A4 _424_.B1 0.28005f
C21902 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I VPWR 0.906f
C21903 _350_.A1 _336_.Z 0.024f
C21904 a_54356_24776# a_54804_24776# 0.01328f
C21905 uio_out[3] uio_out[2] 0.07417f
C21906 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN a_56708_15368# 0.00293f
C21907 a_65780_10664# VPWR 0.22548f
C21908 a_65756_8999# a_65668_9096# 0.28563f
C21909 a_66652_7431# a_66564_7528# 0.28563f
C21910 a_47636_25940# _281_.ZN 0.00228f
C21911 a_67548_5863# a_67460_5960# 0.28563f
C21912 a_15156_21640# a_15156_20452# 0.05841f
C21913 _355_.C a_24092_24679# 0.00239f
C21914 a_37576_29535# VPWR 0.00204f
C21915 a_39236_15368# VPWR 0.20348f
C21916 _340_.A2 a_23556_29860# 0.00119f
C21917 _268_.A2 a_56484_29480# 0.00366f
C21918 _371_.ZN _371_.A1 0.54715f
C21919 a_53704_23219# _281_.A1 0.00415f
C21920 a_42684_15271# VPWR 0.34015f
C21921 _395_.A1 VPWR 1.65268f
C21922 a_4964_14180# a_4604_14136# 0.08674f
C21923 a_2364_14136# a_2812_14136# 0.0131f
C21924 a_40020_16936# a_39996_15704# 0.0016f
C21925 a_43828_16936# a_43940_15748# 0.02666f
C21926 a_66652_17272# VPWR 0.31547f
C21927 a_36100_1256# VPWR 0.20348f
C21928 a_66764_13703# a_66676_13800# 0.28563f
C21929 _218_.ZN a_50280_19369# 0.00148f
C21930 _238_.ZN _238_.I 0.59926f
C21931 _351_.ZN a_24316_26247# 0.03014f
C21932 _330_.A2 _330_.ZN 0.43686f
C21933 a_60276_29032# _252_.ZN 0.17785f
C21934 _386_.ZN _397_.A4 0.03374f
C21935 a_41488_24072# a_42084_24072# 0.00736f
C21936 _355_.C VPWR 4.69272f
C21937 _324_.C _470_.Q 0.14202f
C21938 a_53548_16839# a_53460_16936# 0.28563f
C21939 a_2276_17316# VPWR 0.20634f
C21940 a_12444_1159# a_12804_1256# 0.08717f
C21941 a_51220_16936# VPWR 0.2061f
C21942 a_45596_1592# VPWR 0.29679f
C21943 a_56460_12135# a_57132_12135# 0.00544f
C21944 a_5636_29480# a_6084_29480# 0.01328f
C21945 a_13252_1636# a_13700_1636# 0.01328f
C21946 a_9668_1636# a_9756_1592# 0.28563f
C21947 a_2812_12135# a_3172_12232# 0.08717f
C21948 _416_.A1 a_40132_26344# 0.00561f
C21949 a_34756_17316# a_34396_17272# 0.08707f
C21950 _384_.A3 _419_.Z 0.00268f
C21951 a_64100_11044# a_64188_11000# 0.28563f
C21952 a_42820_31048# a_43268_31048# 0.01328f
C21953 a_16164_2824# VPWR 0.22915f
C21954 a_39536_26795# a_40416_27209# 0.00306f
C21955 a_62196_26724# a_61836_26680# 0.0869f
C21956 _282_.ZN _381_.A2 0.09359f
C21957 _324_.C a_50464_24908# 0.00163f
C21958 _442_.ZN VPWR 0.52428f
C21959 a_42796_23981# VPWR 0.34716f
C21960 _448_.D a_36432_19325# 0.01037f
C21961 a_1468_24679# a_1380_24776# 0.28563f
C21962 _264_.B _433_.ZN 0.02732f
C21963 a_19164_24679# a_19612_24679# 0.01288f
C21964 a_62396_1159# a_62844_1159# 0.0131f
C21965 _459_.CLK a_22059_26399# 0.00978f
C21966 a_30724_26020# a_31116_26020# 0.00705f
C21967 a_1916_19975# a_2364_19975# 0.0131f
C21968 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN a_59732_14180# 0.0027f
C21969 a_2276_14180# VPWR 0.20634f
C21970 a_47076_2824# a_46940_1592# 0.00154f
C21971 a_3260_18407# a_3708_18407# 0.0131f
C21972 a_24636_25641# VPWR 0.3975f
C21973 a_20672_30301# a_19328_28733# 0.00137f
C21974 _290_.ZN a_32240_31048# 0.00141f
C21975 _260_.A1 a_40332_21543# 0.00134f
C21976 a_932_29480# VPWR 0.22176f
C21977 a_35652_15748# a_35740_15704# 0.28563f
C21978 a_51980_12135# VPWR 0.31389f
C21979 a_31708_15704# a_32156_15704# 0.01288f
C21980 _311_.A2 _317_.A2 0.00131f
C21981 a_49316_18504# a_49180_17272# 0.00154f
C21982 a_53012_18504# a_53124_17316# 0.02666f
C21983 _350_.A1 uio_out[0] 0.01434f
C21984 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.02226f
C21985 _248_.B1 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN 0.07658f
C21986 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN a_62980_20072# 0.00109f
C21987 a_5388_24679# VPWR 0.35526f
C21988 _304_.B _397_.A1 0.43204f
C21989 a_19412_27912# uio_out[7] 0.00617f
C21990 _452_.CLK a_44459_18559# 0.03443f
C21991 a_42784_25640# VPWR 0.00205f
C21992 a_42368_28733# a_41996_28777# 0.10745f
C21993 a_34756_15748# VPWR 0.23058f
C21994 a_27908_27912# VPWR 0.00669f
C21995 a_1828_9476# a_1916_9432# 0.28563f
C21996 a_28820_22020# a_28908_21976# 0.28563f
C21997 _452_.CLK a_35723_20569# 0.00491f
C21998 a_47164_18407# a_47612_18407# 0.0131f
C21999 a_24876_21976# a_25324_21976# 0.01288f
C22000 _300_.ZN a_40316_23233# 0.00162f
C22001 a_50860_16839# a_51308_16839# 0.0131f
C22002 _452_.Q a_40244_18180# 0.21456f
C22003 a_49316_14180# a_48956_14136# 0.08707f
C22004 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.00181f
C22005 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN 0.01002f
C22006 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I 0.94181f
C22007 _452_.CLK a_40040_17675# 0.01333f
C22008 _313_.ZN _316_.ZN 0.00267f
C22009 a_50772_16936# a_50884_15748# 0.02666f
C22010 a_5052_25112# a_4964_23588# 0.00151f
C22011 a_46964_16936# a_46940_15704# 0.0016f
C22012 a_46156_16839# VPWR 0.33058f
C22013 _324_.C _260_.A2 0.00499f
C22014 a_58500_1256# VPWR 0.21417f
C22015 a_63204_1256# a_63652_1256# 0.01328f
C22016 _384_.A1 a_48321_23208# 0.00118f
C22017 a_42236_2727# a_42908_2727# 0.00544f
C22018 _448_.Q _319_.A3 0.3777f
C22019 a_54916_21640# a_54780_20408# 0.00154f
C22020 _416_.A3 a_48172_18840# 0.00196f
C22021 a_63316_13800# a_63764_13800# 0.01328f
C22022 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_59260_23111# 0.00332f
C22023 a_45260_17272# a_45260_16839# 0.05841f
C22024 _393_.A1 _393_.A3 0.00414f
C22025 _383_.ZN _395_.A1 0.05542f
C22026 a_36636_17272# VPWR 0.31547f
C22027 a_59396_1636# VPWR 0.20348f
C22028 a_23868_1159# a_23780_1256# 0.28563f
C22029 a_16612_29480# _467_.D 0.01667f
C22030 a_53772_12135# a_53684_12232# 0.28563f
C22031 _395_.A1 a_50068_27508# 0.0015f
C22032 _478_.D a_55060_23263# 0.00177f
C22033 a_11100_29816# a_11548_29816# 0.01288f
C22034 a_15044_29860# a_15132_29816# 0.28563f
C22035 _437_.A1 _441_.B 0.07001f
C22036 a_1380_26344# a_1380_25156# 0.05841f
C22037 a_45172_17316# a_45620_17316# 0.01328f
C22038 _301_.A1 a_38316_20408# 0.00147f
C22039 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_58924_14136# 0.01342f
C22040 _336_.A2 a_26668_23544# 0.00594f
C22041 a_52415_31220# input9.Z 0.01588f
C22042 a_36772_1636# a_36636_1159# 0.00168f
C22043 a_32828_1592# a_32828_1159# 0.05841f
C22044 a_56348_1592# a_56796_1592# 0.01288f
C22045 a_60292_1636# a_60380_1592# 0.28563f
C22046 a_3708_10567# a_4156_10567# 0.0131f
C22047 a_38340_2824# VPWR 0.21435f
C22048 _270_.A2 _255_.I 0.00831f
C22049 _275_.ZN _416_.A1 0.70357f
C22050 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN clk 0.01686f
C22051 a_38764_20408# a_38788_20072# 0.00172f
C22052 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN 0.03123f
C22053 vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN 0.00577f
C22054 a_29692_23111# a_30140_23111# 0.01288f
C22055 a_17484_23111# a_17844_23208# 0.08717f
C22056 _459_.CLK a_19860_27912# 0.00269f
C22057 input9.Z ui_in[7] 0.5414f
C22058 a_21404_24679# a_21764_24776# 0.08707f
C22059 a_45284_9476# VPWR 0.22176f
C22060 _316_.A3 a_37532_21543# 0.00153f
C22061 a_2812_21543# a_3260_21543# 0.0131f
C22062 _317_.A2 a_37444_21640# 0.01533f
C22063 a_51196_14136# VPWR 0.31547f
C22064 a_33948_18407# a_33860_18504# 0.28563f
C22065 _304_.A1 _439_.ZN 0.51613f
C22066 _428_.Z _281_.A1 0.0035f
C22067 a_45732_12232# VPWR 0.20348f
C22068 a_39012_15748# a_38652_15704# 0.08707f
C22069 a_51868_15704# a_52004_15368# 0.00168f
C22070 a_43268_2824# a_43716_2824# 0.01328f
C22071 a_19076_24776# VPWR 0.21778f
C22072 a_1468_20408# a_1468_19975# 0.05841f
C22073 _245_.Z a_61948_26247# 0.03698f
C22074 a_53660_15704# a_53660_15271# 0.05841f
C22075 _397_.A1 VPWR 2.53364f
C22076 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN a_54444_16839# 0.00276f
C22077 a_3708_2727# a_3620_2824# 0.28563f
C22078 _311_.A2 _434_.ZN 0.29421f
C22079 a_61052_26247# a_61500_26247# 0.01255f
C22080 a_40892_15704# VPWR 0.33008f
C22081 a_29804_30951# uo_out[7] 0.01254f
C22082 a_48420_9476# a_48060_9432# 0.08717f
C22083 a_46268_9432# a_46716_9432# 0.0131f
C22084 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN _267_.ZN 0.16475f
C22085 _452_.CLK a_36188_26247# 0.00768f
C22086 a_62172_19975# VPWR 0.31547f
C22087 _416_.A3 a_49034_21640# 0.02383f
C22088 _231_.ZN vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN 0.00632f
C22089 a_55812_14180# a_56260_14180# 0.01328f
C22090 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN VPWR 0.69951f
C22091 a_18828_25112# a_18740_23588# 0.00151f
C22092 a_41440_28363# _330_.A1 0.0031f
C22093 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN a_61276_19975# 0.00153f
C22094 _294_.A2 _284_.ZN 0.28796f
C22095 _261_.ZN _264_.B 0.33177f
C22096 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN a_53572_17316# 0.00118f
C22097 a_4516_12612# a_4604_12568# 0.28563f
C22098 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN _390_.ZN 0.0346f
C22099 a_34939_23705# a_35184_24073# 0.00232f
C22100 a_35232_24029# _304_.A1 0.18089f
C22101 a_37108_23588# a_37556_23588# 0.01328f
C22102 _251_.A1 a_57244_27815# 0.0175f
C22103 a_52316_17272# a_52204_16839# 0.02634f
C22104 _419_.A4 _324_.B 0.20643f
C22105 a_59955_30600# a_60285_30600# 0.53809f
C22106 a_48732_17272# VPWR 0.3158f
C22107 a_1468_1159# VPWR 0.29679f
C22108 a_932_1256# a_1380_1256# 0.01328f
C22109 a_34620_1159# a_35204_1256# 0.01675f
C22110 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].I 0.06892f
C22111 a_64300_12135# a_64884_12232# 0.01675f
C22112 a_50548_12232# a_50996_12232# 0.01328f
C22113 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN clk 0.22004f
C22114 _438_.A2 a_39684_20452# 0.0375f
C22115 _324_.C _250_.B 0.00381f
C22116 a_23332_1636# a_23420_1592# 0.28563f
C22117 a_19388_1592# a_19836_1592# 0.01288f
C22118 a_23108_29860# _459_.CLK 0.02333f
C22119 _365_.ZN a_35818_29860# 0.00124f
C22120 a_29244_21543# VPWR 0.31389f
C22121 a_46852_17316# a_46492_17272# 0.08707f
C22122 _311_.A2 a_36772_23208# 0.01076f
C22123 a_19076_26344# a_19188_25156# 0.02666f
C22124 a_60740_2824# VPWR 0.20348f
C22125 a_1020_10567# a_932_10664# 0.28563f
C22126 a_64996_1636# a_65084_1592# 0.28563f
C22127 _435_.ZN VPWR 0.3363f
C22128 a_23556_24776# a_24004_24776# 0.01328f
C22129 a_28796_23111# a_28708_23208# 0.28563f
C22130 _388_.B _392_.A2 0.00781f
C22131 a_56124_9432# VPWR 0.33981f
C22132 a_66788_14180# VPWR 0.20348f
C22133 _474_.Q clkbuf_1_0__f_clk.I 0.07449f
C22134 a_1468_21543# a_1828_21640# 0.08717f
C22135 _386_.A4 _397_.A4 0.00751f
C22136 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN a_54356_26724# 0.00225f
C22137 _325_.A1 a_40880_23588# 0.01356f
C22138 _230_.I a_61500_27815# 0.00103f
C22139 a_8772_29860# a_8636_29383# 0.00168f
C22140 a_67572_12232# VPWR 0.20595f
C22141 a_45372_15704# a_45820_15704# 0.012f
C22142 _370_.B _369_.ZN 0.03078f
C22143 a_43380_20452# VPWR 0.00542f
C22144 _365_.ZN a_36288_31048# 0.00898f
C22145 a_35740_30951# _462_.D 0.00679f
C22146 a_61724_19975# a_61636_20072# 0.28563f
C22147 a_64412_18840# a_64412_18407# 0.05841f
C22148 a_19035_28409# a_19320_28409# 0.00277f
C22149 _256_.A2 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN 0.05364f
C22150 _346_.A2 a_23332_26344# 0.00302f
C22151 _303_.ZN a_42982_21730# 0.03017f
C22152 _427_.B2 a_52660_21640# 0.00547f
C22153 a_1020_18840# VPWR 0.30073f
C22154 _248_.B1 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I 0.00193f
C22155 a_14684_2727# a_15044_2824# 0.08717f
C22156 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I a_62060_20408# 0.00487f
C22157 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN _407_.ZN 0.00806f
C22158 a_54692_15748# VPWR 0.20623f
C22159 a_66988_19975# a_67436_19975# 0.01255f
C22160 _238_.ZN VPWR 0.30695f
C22161 a_26468_31048# uio_out[1] 0.00583f
C22162 a_49628_17272# a_49540_15748# 0.00151f
C22163 _397_.A1 _383_.ZN 0.609f
C22164 a_62196_23588# VPWR 0.20902f
C22165 a_64748_23111# clk 0.00239f
C22166 a_3172_20452# a_2812_20408# 0.08717f
C22167 a_30388_28776# a_33720_28776# 0.00748f
C22168 _474_.CLK a_55724_22137# 0.00136f
C22169 _252_.ZN a_60516_26344# 0.00538f
C22170 _304_.A1 a_35008_22461# 0.01192f
C22171 a_48868_12612# a_48956_12568# 0.28563f
C22172 a_64636_2727# a_65084_2727# 0.0131f
C22173 a_59332_29816# _238_.ZN 0.001f
C22174 _427_.B1 _427_.ZN 0.13271f
C22175 _407_.A1 _397_.A4 0.54894f
C22176 a_45284_12232# a_45284_11044# 0.05841f
C22177 a_23868_1159# VPWR 0.30141f
C22178 a_46044_1159# a_45956_1256# 0.28563f
C22179 a_65084_12568# a_64996_11044# 0.00151f
C22180 a_67012_9096# a_67012_7908# 0.05841f
C22181 _452_.CLK a_46624_19715# 0.00164f
C22182 a_33412_20072# a_33860_20072# 0.01328f
C22183 a_26692_1636# a_26332_1592# 0.08707f
C22184 a_4852_4392# a_4828_2727# 0.00134f
C22185 hold2.Z _305_.A2 0.32928f
C22186 a_26468_21640# VPWR 0.23321f
C22187 a_53212_17272# a_53660_17272# 0.012f
C22188 a_51532_10567# a_51892_10664# 0.08707f
C22189 a_52639_30644# _274_.A1 0.00162f
C22190 a_6172_1159# a_6620_1159# 0.0131f
C22191 a_65420_10567# a_65868_10567# 0.0131f
C22192 _334_.A1 a_35008_27533# 0.37235f
C22193 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN VPWR 0.72072f
C22194 a_51196_21543# a_49988_21236# 0.00445f
C22195 a_27364_23208# a_27812_23208# 0.01328f
C22196 a_33612_24679# a_34308_24776# 0.01227f
C22197 _324_.C a_44276_20072# 0.01073f
C22198 a_67100_9432# VPWR 0.29679f
C22199 a_16140_23544# VPWR 0.29679f
C22200 _460_.Q _362_.B 2.50636f
C22201 a_33724_21543# a_34396_21543# 0.00544f
C22202 a_3708_2727# VPWR 0.33374f
C22203 a_53772_13703# VPWR 0.31594f
C22204 a_1916_5863# VPWR 0.297f
C22205 a_36100_2824# a_36188_1159# 0.0027f
C22206 a_21852_21543# a_21764_21640# 0.28563f
C22207 _296_.ZN uo_out[1] 0.18727f
C22208 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN a_59260_23544# 0.0099f
C22209 a_15044_29860# uio_oe[1] 0.00278f
C22210 _388_.B _416_.A1 0.05924f
C22211 _474_.CLK vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.02854f
C22212 _384_.A1 a_54040_22366# 0.00133f
C22213 a_15580_29816# a_15580_29383# 0.05841f
C22214 a_48956_11000# VPWR 0.33429f
C22215 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN _324_.C 0.0371f
C22216 a_52676_15748# a_52316_15704# 0.08707f
C22217 a_1020_21976# a_1020_21543# 0.05841f
C22218 a_65668_2824# a_66116_2824# 0.01328f
C22219 _223_.I _358_.A3 0.10453f
C22220 a_4516_26724# VPWR 0.20862f
C22221 a_65084_30951# vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I 0.0151f
C22222 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN a_64996_31048# 0.00711f
C22223 _381_.Z a_50084_24328# 0.22946f
C22224 a_33076_20452# a_33052_19975# 0.00172f
C22225 a_31372_20408# a_31260_19975# 0.02634f
C22226 a_62980_15748# a_63428_15748# 0.01328f
C22227 _281_.ZN _475_.Q 0.02056f
C22228 _452_.Q _302_.Z 0.12437f
C22229 a_16500_26344# VPWR 0.20348f
C22230 a_48508_30951# vgaringosc.workerclkbuff_notouch_.I 0.00613f
C22231 a_26108_2727# a_26020_2824# 0.28563f
C22232 _245_.Z a_61412_26344# 0.02272f
C22233 a_22636_30951# uio_out[3] 0.00309f
C22234 a_64300_23544# clk 0.00613f
C22235 _460_.Q a_32628_26725# 0.12567f
C22236 a_57244_9432# a_57692_9432# 0.0131f
C22237 a_59396_9476# a_59036_9432# 0.08717f
C22238 a_2276_23588# a_2724_23588# 0.01328f
C22239 a_4156_28248# VPWR 0.30552f
C22240 a_2276_6340# a_2724_6340# 0.01328f
C22241 a_38816_27555# _330_.A1 0.01418f
C22242 a_61052_26247# a_60964_26344# 0.28563f
C22243 a_6980_1256# a_7428_1256# 0.01328f
C22244 a_1380_7908# a_1828_7908# 0.01328f
C22245 _478_.D _427_.A2 0.29391f
C22246 _393_.ZN _383_.A2 0.09975f
C22247 a_30924_21976# a_30836_20452# 0.00151f
C22248 a_1380_4772# a_1020_4728# 0.08717f
C22249 a_3172_4772# a_3620_4772# 0.01328f
C22250 a_2276_3204# a_1916_3160# 0.08717f
C22251 a_4068_3204# a_4516_3204# 0.01328f
C22252 a_64188_14136# a_64636_14136# 0.01288f
C22253 _441_.ZN VPWR 0.68694f
C22254 _379_.A2 a_17472_28363# 0.00108f
C22255 _352_.A2 _351_.ZN 0.0508f
C22256 a_55700_23588# a_55788_23544# 0.28563f
C22257 a_5412_1636# VPWR 0.2094f
C22258 a_41160_29083# uo_out[1] 0.01001f
C22259 _459_.CLK a_16052_25156# 0.00236f
C22260 a_54580_13800# a_54668_12135# 0.00151f
C22261 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I a_60940_15704# 0.00681f
C22262 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN 0.61231f
C22263 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN 0.00773f
C22264 a_57580_18840# a_57580_18407# 0.05841f
C22265 clkbuf_1_0__f_clk.I a_46984_23588# 0.01643f
C22266 a_6844_29816# a_6980_29480# 0.00168f
C22267 a_46044_1159# VPWR 0.32517f
C22268 a_57020_1159# a_57380_1256# 0.08717f
C22269 a_17732_31048# uio_oe[0] 0.00296f
C22270 a_33188_1636# a_33636_1636# 0.01328f
C22271 a_2724_11044# a_2364_11000# 0.08717f
C22272 a_4516_11044# a_4964_11044# 0.01328f
C22273 a_64972_16839# a_65420_16839# 0.01222f
C22274 a_63876_18884# VPWR 0.20348f
C22275 a_49068_20408# a_49448_20936# 0.00736f
C22276 _294_.A2 _223_.ZN 0.02376f
C22277 a_50212_20452# a_50660_20452# 0.01328f
C22278 a_57244_27815# a_58020_27508# 0.0121f
C22279 a_43132_27815# a_43580_27815# 0.01255f
C22280 _373_.ZN a_28556_29167# 0.21093f
C22281 _304_.A1 _303_.ZN 0.40292f
C22282 a_62508_10567# a_62420_10664# 0.28563f
C22283 _378_.I uio_out[5] 0.03839f
C22284 a_65668_23208# vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I 0.0035f
C22285 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I 0.01801f
C22286 _304_.B _389_.ZN 0.00863f
C22287 _459_.CLK a_23834_28292# 0.00703f
C22288 a_53108_21640# a_52452_21236# 0.01565f
C22289 a_56484_29480# _241_.I0 0.0016f
C22290 a_58500_21640# vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I 0.00318f
C22291 _337_.A3 _352_.A2 0.05754f
C22292 a_17036_21976# VPWR 0.29679f
C22293 _267_.A2 _274_.A2 0.10592f
C22294 a_30836_23588# VPWR 0.20549f
C22295 a_47524_13800# VPWR 0.20348f
C22296 a_30724_18884# a_31172_18884# 0.01328f
C22297 a_32380_21543# a_32740_21640# 0.08707f
C22298 a_26108_2727# VPWR 0.31664f
C22299 a_3260_29816# VPWR 0.30486f
C22300 _275_.A2 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.01191f
C22301 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I 0.04064f
C22302 _268_.A1 a_52068_29480# 0.01695f
C22303 a_53212_29816# _274_.A2 0.04751f
C22304 _230_.I a_59036_26247# 0.00588f
C22305 a_62756_11044# VPWR 0.20595f
C22306 _284_.B a_44948_25156# 0.0013f
C22307 a_51868_2727# a_52004_1636# 0.00154f
C22308 a_20980_22020# a_20956_21543# 0.00172f
C22309 a_17036_21976# a_17036_21543# 0.05841f
C22310 a_4940_23111# VPWR 0.31945f
C22311 a_51576_25896# _412_.B2 0.00837f
C22312 _260_.ZN a_42796_23981# 0.08579f
C22313 a_5300_27912# VPWR 0.21406f
C22314 a_64300_23111# a_64660_23208# 0.08663f
C22315 a_37084_2727# a_37444_2824# 0.08717f
C22316 _384_.ZN a_48529_22460# 0.02553f
C22317 a_932_25156# a_1380_25156# 0.01328f
C22318 a_2364_6296# a_2364_5863# 0.05841f
C22319 a_65668_6340# a_65308_6296# 0.08717f
C22320 a_1468_7864# a_1468_7431# 0.05841f
C22321 a_64772_7908# a_64412_7864# 0.08717f
C22322 a_62532_20072# a_62532_18884# 0.05841f
C22323 _327_.Z _332_.Z 0.01641f
C22324 a_66564_4772# a_66204_4728# 0.08717f
C22325 a_3260_4728# a_3260_4295# 0.05841f
C22326 a_24116_20452# a_24564_20452# 0.01328f
C22327 a_22772_20452# a_22412_20408# 0.08717f
C22328 _312_.ZN a_34980_22895# 0.03006f
C22329 a_4156_3160# a_4156_2727# 0.05841f
C22330 a_67460_3204# a_67100_3160# 0.08717f
C22331 a_4604_14136# a_4516_12612# 0.0027f
C22332 a_61500_14136# a_61612_13703# 0.02634f
C22333 _424_.B1 a_50940_24072# 0.00844f
C22334 _457_.D a_24988_24679# 0.00613f
C22335 a_11091_30644# a_11460_31048# 0.02397f
C22336 a_67012_17316# a_66988_16839# 0.00172f
C22337 _411_.A2 _384_.A3 0.02921f
C22338 a_11548_1592# VPWR 0.37589f
C22339 a_49316_12612# a_49292_12135# 0.00172f
C22340 a_45372_12568# a_45372_12135# 0.05841f
C22341 a_58588_12568# a_59036_12568# 0.01288f
C22342 _319_.ZN a_34644_20072# 0.03902f
C22343 a_67884_19975# a_67908_18884# 0.0016f
C22344 a_45956_31048# vgaringosc.workerclkbuff_notouch_.I 0.00649f
C22345 a_30240_24776# a_30388_23588# 0.00179f
C22346 a_3620_9096# VPWR 0.22347f
C22347 _351_.A2 a_25184_27209# 0.00112f
C22348 a_33052_19975# VPWR 0.31493f
C22349 a_932_1256# VPWR 0.22176f
C22350 a_64324_5960# VPWR 0.22383f
C22351 _427_.ZN _422_.ZN 0.45364f
C22352 a_47076_11044# a_46716_11000# 0.08707f
C22353 a_34732_18407# VPWR 0.36097f
C22354 _399_.ZN _421_.B 0.00138f
C22355 a_17820_30951# uio_oe[0] 0.00333f
C22356 VPWR uio_out[3] 0.08918f
C22357 a_59284_10664# a_59732_10664# 0.01328f
C22358 a_28572_1159# a_29020_1159# 0.0131f
C22359 a_21316_24776# a_21404_23111# 0.00151f
C22360 _389_.ZN VPWR 0.4246f
C22361 _258_.I a_59572_29076# 0.8526f
C22362 a_2812_26680# a_2812_26247# 0.05841f
C22363 a_30836_22020# VPWR 0.20595f
C22364 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN 0.00786f
C22365 _304_.ZN a_43666_21812# 0.00161f
C22366 a_48508_2727# VPWR 0.31143f
C22367 a_1828_12612# VPWR 0.20348f
C22368 a_30948_21640# a_31396_21640# 0.01328f
C22369 a_36500_29860# VPWR 0.01707f
C22370 a_50196_21640# a_49988_21236# 0.02745f
C22371 a_15692_26247# a_15604_26344# 0.28563f
C22372 a_5052_3160# a_4964_1636# 0.0027f
C22373 _231_.ZN a_59260_23111# 0.00497f
C22374 uio_oe[4] uio_oe[3] 0.03708f
C22375 _350_.A2 a_29716_31048# 0.06853f
C22376 a_32516_15368# a_32964_15368# 0.01328f
C22377 a_17060_29860# VPWR 0.20845f
C22378 a_49740_10567# VPWR 0.32073f
C22379 _330_.A1 _447_.Q 0.05414f
C22380 _301_.A1 a_34715_22137# 0.00492f
C22381 a_27924_22020# a_27900_21543# 0.00172f
C22382 a_23980_21976# a_24092_21543# 0.02634f
C22383 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I a_61188_15368# 0.00761f
C22384 a_33956_31048# uo_out[5] 0.01666f
C22385 a_34620_15271# a_34532_15368# 0.28563f
C22386 a_2276_23208# VPWR 0.20634f
C22387 _437_.A1 _452_.Q 0.01253f
C22388 a_35964_15271# a_36412_15271# 0.0131f
C22389 a_24564_31048# uio_out[3] 0.01582f
C22390 a_29804_30951# _459_.Q 0.01816f
C22391 _350_.A1 _287_.A1 0.35586f
C22392 a_63092_26724# vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN 0.00691f
C22393 a_48508_2727# a_48420_2824# 0.28563f
C22394 a_3172_22020# a_3620_22020# 0.01328f
C22395 _230_.I _247_.ZN 0.40781f
C22396 a_1380_22020# a_1020_21976# 0.08717f
C22397 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I 0.87069f
C22398 a_64772_17316# a_64412_17272# 0.08717f
C22399 _241_.I0 a_55956_25940# 0.00234f
C22400 a_32476_29167# a_32820_29535# 0.00275f
C22401 _474_.CLK a_47525_29480# 0.00481f
C22402 a_4940_8999# a_5388_8999# 0.01222f
C22403 a_5300_23208# a_5388_21543# 0.0027f
C22404 a_20620_23544# a_21068_23544# 0.01288f
C22405 a_64412_7431# a_64860_7431# 0.0131f
C22406 a_65308_5863# a_65756_5863# 0.0131f
C22407 a_29380_1256# a_29828_1256# 0.01328f
C22408 a_66204_4295# a_66652_4295# 0.0131f
C22409 _462_.D VPWR 0.41136f
C22410 a_4940_13703# a_5300_13800# 0.08674f
C22411 a_66787_30600# a_67237_30644# 0.00184f
C22412 a_40468_16936# a_40668_15271# 0.00119f
C22413 a_8636_2727# a_9084_2727# 0.0131f
C22414 a_58476_13703# a_58924_13703# 0.01288f
C22415 a_48956_14136# a_48868_12612# 0.0027f
C22416 _437_.ZN VPWR 0.41169f
C22417 a_60516_26344# a_60964_26344# 0.01328f
C22418 a_66004_18504# a_66116_17316# 0.02666f
C22419 _424_.A2 a_51332_24072# 0.14193f
C22420 _251_.A1 a_58063_30644# 0.00922f
C22421 a_31260_16839# a_31620_16936# 0.08717f
C22422 _384_.A3 _399_.ZN 0.35237f
C22423 a_18472_29076# uio_out[7] 0.00122f
C22424 a_25348_1636# VPWR 0.20957f
C22425 a_54780_18840# vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN 0.0014f
C22426 a_65892_12612# a_65980_12568# 0.28563f
C22427 _258_.I _257_.B 0.28073f
C22428 a_3708_23544# a_3708_23111# 0.05841f
C22429 _371_.A1 _336_.A2 0.12111f
C22430 a_12548_31048# a_13004_30951# 0.0065f
C22431 _304_.B a_42148_27912# 0.00598f
C22432 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I 0.13254f
C22433 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_60212_25156# 0.02858f
C22434 _287_.A2 a_31068_28292# 0.00267f
C22435 a_62980_18504# a_63428_18504# 0.01328f
C22436 _402_.A1 a_43564_27209# 0.03607f
C22437 a_1828_15368# a_1828_14180# 0.05841f
C22438 a_55228_20408# a_55340_19975# 0.02634f
C22439 _359_.B uo_out[6] 0.07456f
C22440 a_43268_1636# a_43356_1592# 0.28563f
C22441 a_46852_1636# a_47300_1636# 0.01328f
C22442 a_53572_11044# a_54020_11044# 0.01328f
C22443 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN 0.00457f
C22444 a_44724_16936# a_45172_16936# 0.01328f
C22445 _452_.CLK _264_.B 0.00154f
C22446 _443_.D a_37892_26344# 0.00109f
C22447 _359_.B a_28054_30196# 0.75292f
C22448 a_4604_26680# a_5052_26680# 0.01222f
C22449 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I a_65756_27815# 0.00842f
C22450 a_25962_29480# VPWR 0.01533f
C22451 a_43736_25896# a_44340_26183# 0.49241f
C22452 a_32740_2824# a_32740_1636# 0.05841f
C22453 a_45416_29885# _386_.A4 0.00109f
C22454 a_56572_29383# a_56484_29480# 0.28563f
C22455 _448_.Q _305_.A2 0.44319f
C22456 a_15604_20452# VPWR 0.20348f
C22457 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_63764_23208# 0.00385f
C22458 _384_.A1 _399_.A1 0.42711f
C22459 a_50748_12568# VPWR 0.32481f
C22460 _284_.ZN a_40644_29480# 0.00232f
C22461 _359_.B a_44160_29123# 0.01916f
C22462 a_22059_26399# a_22352_25987# 0.49319f
C22463 a_9444_2824# a_9892_2824# 0.01328f
C22464 a_7068_29383# a_7428_29480# 0.08717f
C22465 _452_.CLK _332_.Z 0.07775f
C22466 _241_.Z vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.03181f
C22467 _383_.ZN _389_.ZN 0.01137f
C22468 a_3708_28248# a_3708_27815# 0.05841f
C22469 a_3620_10664# VPWR 0.22347f
C22470 a_22636_21976# a_22660_21640# 0.00172f
C22471 a_45372_15271# a_45956_15368# 0.01675f
C22472 _316_.ZN a_33724_21543# 0.01469f
C22473 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN _245_.I1 0.0549f
C22474 a_33188_23208# VPWR 0.2051f
C22475 a_36100_26724# a_36548_26724# 0.01328f
C22476 a_34308_24776# a_34304_24029# 0.00375f
C22477 _352_.A2 a_29828_26344# 0.15085f
C22478 _245_.Z vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN 0.00863f
C22479 _476_.Q a_51428_20452# 0.0031f
C22480 a_38336_18147# VPWR 0.18842f
C22481 _324_.C a_50084_24328# 0.06569f
C22482 a_15692_28248# a_16140_28248# 0.01255f
C22483 a_15156_22020# a_14796_21976# 0.08707f
C22484 _447_.Q _226_.ZN 0.03458f
C22485 a_59484_2727# a_59844_2824# 0.08717f
C22486 a_62980_15368# a_63428_15368# 0.01328f
C22487 a_62620_15704# VPWR 0.29679f
C22488 _459_.CLK uo_out[4] 0.00167f
C22489 a_43804_30951# a_44164_31048# 0.08717f
C22490 _358_.A3 a_36636_26680# 0.00221f
C22491 a_52676_27912# _412_.ZN 0.00116f
C22492 a_56596_18504# a_57044_18504# 0.01328f
C22493 _359_.B uo_out[5] 0.00253f
C22494 a_19076_31048# VPWR 0.22145f
C22495 a_28372_23588# a_28460_23544# 0.28563f
C22496 a_2812_7864# VPWR 0.30213f
C22497 a_19276_25112# a_19724_25112# 0.01288f
C22498 a_13252_1256# VPWR 0.20348f
C22499 a_4604_4728# VPWR 0.33016f
C22500 a_52871_31198# VPWR 0.00419f
C22501 a_27676_26680# VPWR 0.29869f
C22502 a_33052_18840# a_33052_18407# 0.05841f
C22503 a_3708_29383# VPWR 0.33374f
C22504 _350_.A1 a_28000_29480# 0.00303f
C22505 a_55564_13703# a_55476_13800# 0.28563f
C22506 a_53300_23047# a_54088_22895# 0.02112f
C22507 a_51668_16936# a_51644_15271# 0.00134f
C22508 a_21740_30951# uio_out[5] 0.00668f
C22509 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN a_57916_25112# 0.0032f
C22510 a_42572_16839# a_42484_16936# 0.28563f
C22511 a_39012_1636# VPWR 0.20348f
C22512 a_45372_12135# a_45820_12135# 0.0131f
C22513 a_1020_1159# a_1380_1256# 0.08717f
C22514 a_3620_16936# VPWR 0.22347f
C22515 a_42148_27912# VPWR 0.2372f
C22516 a_2364_1592# a_2812_1592# 0.01288f
C22517 a_6308_1636# a_6396_1592# 0.28563f
C22518 _476_.Q a_53884_20408# 0.01164f
C22519 _346_.B a_22548_28292# 0.0011f
C22520 a_1380_29860# a_1020_29816# 0.08707f
C22521 a_4516_17316# a_4604_17272# 0.28563f
C22522 _241_.I0 a_55676_27815# 0.0027f
C22523 a_56124_28248# a_56124_27815# 0.05841f
C22524 _447_.Q _300_.ZN 0.69551f
C22525 _268_.A2 uio_in[1] 0.03537f
C22526 a_63316_12232# a_63404_10567# 0.00151f
C22527 a_60292_11044# a_60964_11044# 0.00347f
C22528 _352_.A2 a_27328_25227# 0.03116f
C22529 a_18492_1592# a_18492_1159# 0.05841f
C22530 a_22436_1636# a_22300_1159# 0.00168f
C22531 _474_.CLK vgaringosc.workerclkbuff_notouch_.I 2.11003f
C22532 _330_.A1 a_41432_17801# 0.00583f
C22533 a_36860_23111# a_36772_23208# 0.28563f
C22534 _251_.A1 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I 0.15111f
C22535 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN VPWR 1.48456f
C22536 _304_.B a_39536_26795# 0.00702f
C22537 a_50972_1159# a_51420_1159# 0.0131f
C22538 a_45820_18407# a_46180_18504# 0.08717f
C22539 _474_.CLK a_53124_27912# 0.00539f
C22540 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN 0.66304f
C22541 a_2364_25112# VPWR 0.30029f
C22542 a_63516_18407# VPWR 0.29679f
C22543 a_64324_18884# a_64412_18840# 0.28563f
C22544 a_26580_20452# VPWR 0.2131f
C22545 a_4156_27815# a_4068_27912# 0.28563f
C22546 _256_.A2 a_65072_29860# 0.02416f
C22547 a_57044_18504# a_57044_17316# 0.05841f
C22548 a_19372_30345# VPWR 0.43044f
C22549 a_64548_12612# VPWR 0.21169f
C22550 a_3260_15704# a_3708_15704# 0.0131f
C22551 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I VPWR 0.72735f
C22552 a_40038_28720# uo_out[1] 0.00129f
C22553 _447_.Q a_35723_20569# 0.02761f
C22554 a_37532_15704# a_37668_15368# 0.00168f
C22555 a_54916_15368# a_55364_15368# 0.01328f
C22556 a_55228_15704# VPWR 0.34302f
C22557 _330_.A1 a_45169_27509# 0.00552f
C22558 _371_.ZN _349_.A4 0.0011f
C22559 _311_.A2 a_37556_23588# 0.00885f
C22560 a_65308_8999# a_65668_9096# 0.08717f
C22561 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN clk 0.45884f
C22562 a_65332_10664# VPWR 0.21332f
C22563 a_39460_15748# a_39324_15271# 0.00168f
C22564 _373_.A2 _359_.B 0.40601f
C22565 _371_.A1 a_34532_27208# 0.00122f
C22566 a_66204_7431# a_66564_7528# 0.08717f
C22567 a_32268_21976# a_32292_21640# 0.00172f
C22568 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN 0.8877f
C22569 a_56796_15271# a_56708_15368# 0.28563f
C22570 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I 0.00383f
C22571 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I a_57380_16936# 0.07139f
C22572 a_67100_5863# a_67460_5960# 0.08717f
C22573 a_23644_21543# a_23668_20452# 0.0016f
C22574 _355_.C a_23644_24679# 0.00241f
C22575 _301_.A1 _301_.Z 0.00701f
C22576 a_36628_29535# VPWR 0.00246f
C22577 a_38788_15368# VPWR 0.20348f
C22578 a_56684_18407# vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I 0.00209f
C22579 a_21516_21976# a_21964_21976# 0.012f
C22580 a_42236_15271# VPWR 0.31029f
C22581 a_17803_26841# a_18088_26841# 0.00277f
C22582 a_4516_14180# a_4604_14136# 0.28563f
C22583 a_39660_16839# a_40108_16839# 0.01288f
C22584 a_66204_17272# VPWR 0.33522f
C22585 a_35652_1256# VPWR 0.20348f
C22586 a_33376_23659# _313_.ZN 0.25429f
C22587 a_51780_1256# a_52228_1256# 0.01328f
C22588 _218_.ZN a_50384_19204# 0.00315f
C22589 a_50188_13703# a_50212_12612# 0.0016f
C22590 _351_.ZN a_23868_26247# 0.00125f
C22591 _330_.A2 a_37408_18504# 0.04634f
C22592 a_52340_13800# a_52788_13800# 0.01328f
C22593 a_30812_2727# a_31484_2727# 0.00544f
C22594 a_66316_13703# a_66676_13800# 0.08717f
C22595 a_19164_30951# VPWR 0.35785f
C22596 a_41488_24072# a_41880_24072# 0.00629f
C22597 a_57044_17316# a_57492_17316# 0.01328f
C22598 a_35292_17272# a_35180_16839# 0.02634f
C22599 a_53100_16839# a_53460_16936# 0.08717f
C22600 _419_.Z _417_.Z 0.02301f
C22601 _274_.A2 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.00234f
C22602 a_1828_17316# VPWR 0.20348f
C22603 a_50772_16936# VPWR 0.2156f
C22604 _397_.A2 _421_.B 0.0032f
C22605 a_45148_1592# VPWR 0.29679f
C22606 a_12444_1159# a_12356_1256# 0.28563f
C22607 a_52540_1592# a_52676_1256# 0.00168f
C22608 a_48708_29816# _392_.A2 0.00591f
C22609 _452_.CLK a_44786_24120# 0.00261f
C22610 a_2812_12135# a_2724_12232# 0.28563f
C22611 a_9668_1636# a_9308_1592# 0.08707f
C22612 a_27564_23544# a_27452_23111# 0.02634f
C22613 a_7740_29816# a_8188_29816# 0.012f
C22614 _416_.A1 a_39684_26344# 0.02402f
C22615 a_34308_17316# a_34396_17272# 0.28563f
C22616 a_39536_26795# a_39924_27209# 0.00393f
C22617 vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN VPWR 0.7672f
C22618 a_67236_11044# a_67684_11044# 0.01328f
C22619 a_64100_11044# a_63740_11000# 0.08707f
C22620 a_52988_1592# a_53436_1592# 0.01288f
C22621 a_61748_26724# a_61836_26680# 0.28563f
C22622 a_15492_2824# VPWR 0.20968f
C22623 _395_.A1 _407_.ZN 0.00725f
C22624 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I VPWR 0.74172f
C22625 a_41488_24072# VPWR 0.81484f
C22626 _448_.D a_35504_18955# 0.28404f
C22627 a_39536_26795# VPWR 1.10054f
C22628 a_18716_23111# a_19164_23111# 0.01288f
C22629 _459_.CLK a_21052_26031# 0.0422f
C22630 a_1020_24679# a_1380_24776# 0.08717f
C22631 a_30724_26020# a_30932_26020# 0.00478f
C22632 a_64972_26680# a_64860_26247# 0.02634f
C22633 _437_.A1 _436_.B 0.00277f
C22634 a_1828_14180# VPWR 0.20348f
C22635 a_5052_7864# a_4964_6340# 0.00151f
C22636 a_25008_25597# VPWR 0.18871f
C22637 a_19860_27912# a_20308_27912# 0.01328f
C22638 _474_.CLK _427_.B1 0.0106f
C22639 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN 0.08661f
C22640 _260_.A1 _432_.ZN 0.11386f
C22641 a_35652_15748# a_35292_15704# 0.08707f
C22642 a_51532_12135# VPWR 0.31389f
C22643 a_20003_29611# VPWR 0.49244f
C22644 a_31844_2824# a_32292_2824# 0.01328f
C22645 _311_.A2 a_36148_21976# 0.49323f
C22646 a_4940_24679# VPWR 0.31945f
C22647 ena clk 0.03868f
C22648 _476_.Q _281_.A1 1.15826f
C22649 uo_out[2] uo_out[3] 0.08179f
C22650 a_17844_27912# uio_out[7] 0.00368f
C22651 _452_.CLK a_43452_18191# 0.02286f
C22652 a_22212_21640# a_22324_20452# 0.02666f
C22653 _251_.A1 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I 0.14509f
C22654 a_34308_15748# VPWR 0.21526f
C22655 _355_.C a_28679_24776# 0.00406f
C22656 _252_.ZN _245_.Z 0.22353f
C22657 a_26916_27912# VPWR 0.22859f
C22658 _274_.A1 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.00329f
C22659 a_3620_9476# a_4068_9476# 0.01328f
C22660 a_1828_9476# a_1468_9432# 0.08717f
C22661 a_28820_22020# a_28460_21976# 0.08707f
C22662 _252_.ZN a_60604_26247# 0.00621f
C22663 _452_.Q a_39264_18147# 0.01473f
C22664 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN VPWR 0.74245f
C22665 a_58656_27912# a_58020_27508# 0.02745f
C22666 a_48868_14180# a_48956_14136# 0.28563f
C22667 a_54356_20072# a_54244_18884# 0.02666f
C22668 a_57580_18840# a_58028_18840# 0.01255f
C22669 _300_.ZN a_40004_23233# 0.00196f
C22670 _313_.ZN a_33152_22091# 0.00427f
C22671 _452_.CLK a_39236_17316# 0.00649f
C22672 a_45708_16839# VPWR 0.29679f
C22673 a_22548_31048# uio_out[5] 0.00117f
C22674 a_58052_1256# VPWR 0.24377f
C22675 _384_.A1 a_52920_22760# 0.18999f
C22676 a_47076_13800# a_47076_12612# 0.05841f
C22677 _416_.A3 a_47724_18840# 0.01123f
C22678 a_66876_14136# a_66788_12612# 0.00151f
C22679 _448_.Q a_37532_21543# 0.06439f
C22680 a_57132_13703# a_57156_12612# 0.0016f
C22681 a_64188_27815# vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I 0.00391f
C22682 a_36188_17272# VPWR 0.31547f
C22683 a_63764_10664# a_63652_9476# 0.02666f
C22684 a_61972_10664# a_61948_9432# 0.0016f
C22685 a_58948_1636# VPWR 0.20348f
C22686 a_23196_1159# a_23780_1256# 0.01675f
C22687 a_16028_1592# a_16612_1636# 0.01675f
C22688 a_67212_12135# a_67660_12135# 0.0131f
C22689 a_53324_12135# a_53684_12232# 0.08707f
C22690 a_16612_29480# a_17060_29480# 0.01328f
C22691 a_16164_29480# _467_.D 0.00383f
C22692 a_15044_29860# a_14684_29816# 0.08707f
C22693 _412_.A1 a_52360_26355# 0.00298f
C22694 a_40644_17272# a_41048_17341# 0.41635f
C22695 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN a_54804_16936# 0.00241f
C22696 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_57692_14136# 0.00643f
C22697 a_53124_27912# a_52988_26680# 0.00154f
C22698 a_55700_25156# clk 0.00367f
C22699 a_37892_2824# VPWR 0.20815f
C22700 a_60292_1636# a_59932_1592# 0.08707f
C22701 a_54432_31128# ui_in[7] 0.389f
C22702 _459_.CLK a_19412_27912# 0.00563f
C22703 a_17484_23111# a_17396_23208# 0.28563f
C22704 a_21404_24679# a_21316_24776# 0.28563f
C22705 _252_.ZN _252_.B 0.11369f
C22706 a_3172_24776# a_3620_24776# 0.01328f
C22707 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN VPWR 0.84133f
C22708 a_5052_9432# VPWR 0.33516f
C22709 a_67012_9096# a_67460_9096# 0.01328f
C22710 ui_in[3] ui_in[2] 0.25051f
C22711 _316_.A3 a_37084_21543# 0.00796f
C22712 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN 0.00249f
C22713 a_50748_14136# VPWR 0.32481f
C22714 a_2724_18504# a_3172_18504# 0.01328f
C22715 _400_.ZN _282_.ZN 0.03008f
C22716 a_33500_18407# a_33860_18504# 0.08717f
C22717 _388_.B a_45012_29816# 0.01878f
C22718 _379_.A2 a_21204_31048# 0.14142f
C22719 a_33776_29123# a_34084_28776# 0.00106f
C22720 _399_.A1 clk 0.0015f
C22721 a_38564_15748# a_38652_15704# 0.28563f
C22722 a_42148_15748# a_42596_15748# 0.01328f
C22723 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN 0.00123f
C22724 a_45284_12232# VPWR 0.22176f
C22725 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN 0.00609f
C22726 a_31844_26344# a_31732_25156# 0.02666f
C22727 _384_.ZN _281_.ZN 0.04388f
C22728 _417_.A2 a_52036_22504# 0.0014f
C22729 _245_.Z a_61500_26247# 0.02967f
C22730 a_18628_24776# VPWR 0.23332f
C22731 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN a_53996_16839# 0.00144f
C22732 a_42392_19243# a_42996_18840# 0.49241f
C22733 a_3260_2727# a_3620_2824# 0.08717f
C22734 a_40444_15704# VPWR 0.3289f
C22735 a_5388_19975# a_5300_20072# 0.28563f
C22736 _334_.A1 _365_.ZN 0.13283f
C22737 _290_.ZN _287_.A1 1.99814f
C22738 _402_.A1 _392_.A2 0.16262f
C22739 a_47972_9476# a_48060_9432# 0.28563f
C22740 a_33152_22091# _316_.ZN 0.26168f
C22741 _223_.ZN a_32580_27912# 0.00113f
C22742 a_61724_19975# VPWR 0.31589f
C22743 a_65756_27815# VPWR 0.34369f
C22744 _452_.CLK a_35740_26247# 0.00857f
C22745 _417_.A2 a_48888_19243# 0.02352f
C22746 a_1916_12568# a_2364_12568# 0.0131f
C22747 a_4516_12612# a_4156_12568# 0.08674f
C22748 a_54132_13800# a_54020_12612# 0.02666f
C22749 a_53212_2727# a_53660_2727# 0.0131f
C22750 a_33932_24073# _304_.A1 0.00136f
C22751 _251_.A1 _229_.I 0.71897f
C22752 _419_.A4 a_47860_23208# 0.03829f
C22753 a_48284_17272# VPWR 0.31389f
C22754 a_34620_1159# a_34532_1256# 0.28563f
C22755 a_1020_1159# VPWR 0.30073f
C22756 a_23332_1636# a_22972_1592# 0.08707f
C22757 a_1380_5960# a_1380_4772# 0.05841f
C22758 _324_.C a_63952_29480# 0.00995f
C22759 a_64300_12135# a_64212_12232# 0.28563f
C22760 a_2276_4392# a_2276_3204# 0.05841f
C22761 _330_.A1 _451_.Q 0.08808f
C22762 a_22560_30288# _459_.CLK 0.5617f
C22763 a_23108_29860# a_23556_29860# 0.01328f
C22764 a_28796_21543# VPWR 0.31389f
C22765 _246_.B2 a_59828_26724# 0.00358f
C22766 a_49988_17316# a_50436_17316# 0.01328f
C22767 a_46404_17316# a_46492_17272# 0.28563f
C22768 a_40880_23588# VPWR 0.01366f
C22769 a_54220_10567# a_54668_10567# 0.01288f
C22770 a_60292_2824# VPWR 0.20348f
C22771 a_64996_1636# a_64636_1592# 0.08717f
C22772 a_66788_1636# a_67236_1636# 0.01328f
C22773 _284_.ZN _435_.A3 0.03993f
C22774 _362_.ZN _335_.ZN 0.05963f
C22775 a_28348_23111# a_28708_23208# 0.08707f
C22776 a_16052_23208# a_16500_23208# 0.01328f
C22777 a_55676_9432# VPWR 0.31143f
C22778 a_1468_21543# a_1380_21640# 0.28563f
C22779 a_22748_21543# a_23196_21543# 0.01288f
C22780 a_24676_2824# a_24764_1159# 0.0027f
C22781 a_66340_14180# VPWR 0.21266f
C22782 vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I a_66540_19975# 0.0023f
C22783 _455_.Q _345_.A2 0.3451f
C22784 _398_.C _427_.B1 0.33765f
C22785 a_66787_30600# ena 0.0063f
C22786 _408_.ZN _395_.A2 0.01705f
C22787 a_67124_12232# VPWR 0.20595f
C22788 _324_.C vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN 0.02872f
C22789 _474_.CLK _422_.ZN 0.00103f
C22790 a_37532_2727# a_37668_1636# 0.00154f
C22791 a_54244_2824# a_54692_2824# 0.01328f
C22792 a_43156_20452# VPWR 0.00439f
C22793 a_61276_19975# a_61636_20072# 0.08717f
C22794 _365_.ZN a_35652_31048# 0.02071f
C22795 _303_.ZN a_42778_21812# 0.003f
C22796 a_37472_24419# VPWR 0.51569f
C22797 _355_.C a_20756_26724# 0.00125f
C22798 a_4964_18884# VPWR 0.21167f
C22799 _359_.B _460_.Q 0.76382f
C22800 a_14684_2727# a_14596_2824# 0.28563f
C22801 a_44340_26183# a_44736_26031# 0.00232f
C22802 a_54244_15748# VPWR 0.2274f
C22803 _260_.A2 _432_.ZN 0.17966f
C22804 a_53348_9476# a_53796_9476# 0.01328f
C22805 a_26020_31048# uio_out[1] 0.00325f
C22806 _430_.ZN a_39178_23208# 0.02369f
C22807 a_61748_23588# VPWR 0.228f
C22808 a_60268_14136# a_60964_14180# 0.01227f
C22809 a_64300_23111# clk 0.00239f
C22810 a_46268_14136# a_46268_13703# 0.05841f
C22811 a_50212_14180# a_50188_13703# 0.00172f
C22812 a_30388_28776# a_33312_28776# 0.00951f
C22813 a_2724_20452# a_2812_20408# 0.28563f
C22814 _416_.A1 _402_.A1 0.06696f
C22815 _252_.ZN a_60013_26344# 0.00322f
C22816 _304_.A1 a_33708_22505# 0.00265f
C22817 a_48868_12612# a_48508_12568# 0.08707f
C22818 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN a_58588_26247# 0.0064f
C22819 a_61076_13800# a_60964_12612# 0.02666f
C22820 a_15156_24776# a_15156_23588# 0.05841f
C22821 a_23196_1159# VPWR 0.35728f
C22822 a_45596_1159# a_45956_1256# 0.08717f
C22823 a_61076_12232# a_61524_12232# 0.01328f
C22824 a_26244_1636# a_26332_1592# 0.28563f
C22825 a_29828_1636# a_30276_1636# 0.01328f
C22826 a_25796_21640# VPWR 0.21858f
C22827 a_59260_23111# clk 0.00239f
C22828 a_50660_1636# a_50524_1159# 0.00168f
C22829 a_51532_10567# a_51444_10664# 0.28563f
C22830 _325_.A2 _327_.Z 0.21044f
C22831 _451_.Q _226_.ZN 0.00572f
C22832 _424_.B1 a_51892_23340# 0.00244f
C22833 a_64660_23208# VPWR 0.21234f
C22834 _274_.A1 ui_in[7] 0.00327f
C22835 a_60405_31198# VPWR 0.00423f
C22836 a_1468_5863# VPWR 0.29679f
C22837 a_66452_20072# a_66900_20072# 0.01328f
C22838 a_21404_21543# a_21764_21640# 0.08707f
C22839 a_66652_9432# VPWR 0.29679f
C22840 a_15692_23544# VPWR 0.29679f
C22841 _251_.A1 rst_n 0.02683f
C22842 _363_.Z _358_.A3 0.00177f
C22843 a_53324_13703# VPWR 0.31598f
C22844 a_3260_2727# VPWR 0.30487f
C22845 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I a_61972_20452# 0.03006f
C22846 _351_.A2 a_25524_26344# 0.00539f
C22847 _412_.A1 _395_.A2 0.45518f
C22848 _433_.ZN _302_.Z 0.03843f
C22849 a_48508_11000# VPWR 0.29679f
C22850 a_52228_15748# a_52316_15704# 0.28563f
C22851 a_48284_15704# a_48732_15704# 0.01288f
C22852 a_31964_28292# VPWR 0.00979f
C22853 a_4068_26724# VPWR 0.2157f
C22854 a_54444_23544# a_54892_23544# 0.0131f
C22855 a_65084_30951# a_64996_31048# 0.28563f
C22856 _223_.I a_31484_26680# 0.03118f
C22857 _399_.ZN _402_.B 0.43226f
C22858 _451_.Q _300_.ZN 0.15143f
C22859 a_16052_26344# VPWR 0.20348f
C22860 a_48060_30951# vgaringosc.workerclkbuff_notouch_.I 0.00613f
C22861 _231_.ZN VPWR 0.47193f
C22862 a_25660_2727# a_26020_2824# 0.08717f
C22863 _245_.Z a_60964_26344# 0.01663f
C22864 a_63852_23544# clk 0.00232f
C22865 a_29716_31048# _370_.ZN 0.00196f
C22866 _287_.A2 a_29232_29931# 0.01715f
C22867 _355_.C _378_.I 0.4032f
C22868 a_3708_28248# VPWR 0.33374f
C22869 a_58948_9476# a_59036_9432# 0.28563f
C22870 a_60604_26247# a_60964_26344# 0.0869f
C22871 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN 0.01625f
C22872 _260_.A2 a_44948_22020# 0.00311f
C22873 a_38523_27967# _330_.A1 0.00702f
C22874 a_1828_3204# a_1916_3160# 0.28563f
C22875 a_57156_14180# a_57132_13703# 0.00172f
C22876 a_53660_14136# a_53772_13703# 0.02634f
C22877 a_67684_14180# a_67772_14136# 0.28563f
C22878 a_16588_20408# a_17036_20408# 0.0131f
C22879 _359_.B _416_.A1 0.14917f
C22880 a_50084_24328# a_50724_24908# 0.0101f
C22881 a_55700_23588# a_55340_23544# 0.08717f
C22882 a_4964_1636# VPWR 0.20815f
C22883 _287_.A2 _335_.ZN 0.01262f
C22884 a_55364_12612# a_55812_12612# 0.01328f
C22885 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _407_.A1 0.00141f
C22886 _439_.ZN _301_.A1 0.00109f
C22887 _441_.ZN a_39780_22805# 0.48433f
C22888 a_57020_1159# a_56932_1256# 0.28563f
C22889 a_45596_1159# VPWR 0.29679f
C22890 _451_.Q a_40040_17675# 0.00939f
C22891 a_17284_31048# uio_oe[0] 0.01582f
C22892 a_2276_11044# a_2364_11000# 0.28563f
C22893 a_63428_18884# VPWR 0.20348f
C22894 _395_.A2 a_51968_26724# 0.00927f
C22895 _268_.A2 _275_.ZN 0.02625f
C22896 _373_.ZN a_28928_29123# 0.00739f
C22897 _467_.D a_17484_27815# 0.00304f
C22898 a_47972_10664# a_48420_10664# 0.01328f
C22899 a_57604_1636# a_57468_1159# 0.00168f
C22900 a_17148_1159# a_17596_1159# 0.0131f
C22901 a_4852_18504# a_4964_17316# 0.02666f
C22902 a_62060_10567# a_62420_10664# 0.08707f
C22903 a_18404_2824# a_18404_1636# 0.05841f
C22904 _397_.A2 a_50996_28292# 0.00695f
C22905 a_56148_23588# a_56596_23588# 0.01328f
C22906 a_16588_21976# VPWR 0.29679f
C22907 a_52660_21640# a_52452_21236# 0.02745f
C22908 a_30388_23588# VPWR 0.22449f
C22909 a_32380_21543# a_32292_21640# 0.28563f
C22910 a_19972_21640# a_20420_21640# 0.01328f
C22911 a_25660_2727# VPWR 0.31485f
C22912 _260_.A1 _260_.A2 0.47414f
C22913 a_47076_2824# a_47164_1159# 0.0027f
C22914 a_47076_13800# VPWR 0.20348f
C22915 a_63516_15271# a_63964_15271# 0.0131f
C22916 a_61297_30300# ui_in[3] 0.03393f
C22917 a_2812_29816# VPWR 0.30213f
C22918 a_62308_11044# VPWR 0.20595f
C22919 _459_.CLK _358_.A2 0.00214f
C22920 _431_.A3 a_39684_26344# 0.00509f
C22921 a_4156_23111# VPWR 0.3269f
C22922 a_59260_23544# a_59260_23111# 0.05841f
C22923 _268_.A1 _272_.A2 0.00394f
C22924 _276_.A2 _274_.A2 0.08976f
C22925 a_26556_27815# a_27004_27815# 0.01222f
C22926 a_67100_15704# a_67548_15704# 0.01222f
C22927 a_50120_26476# _412_.B2 0.03745f
C22928 a_4852_27912# VPWR 0.22733f
C22929 a_64300_23111# a_64212_23208# 0.28563f
C22930 a_37084_2727# a_36996_2824# 0.28563f
C22931 _419_.A4 _421_.A1 0.70418f
C22932 a_44632_30206# a_44795_29535# 0.00103f
C22933 _411_.A2 a_51436_27208# 0.00144f
C22934 a_52228_19368# a_53436_18840# 0.00445f
C22935 vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN a_58028_20408# 0.0067f
C22936 a_66116_7908# a_66564_7908# 0.01328f
C22937 a_64324_7908# a_64412_7864# 0.28563f
C22938 a_17396_23588# a_17844_23588# 0.01328f
C22939 a_64324_9476# a_64772_9476# 0.01328f
C22940 a_17956_1256# a_18404_1256# 0.01328f
C22941 a_65220_6340# a_65308_6296# 0.28563f
C22942 a_67012_6340# a_67460_6340# 0.01328f
C22943 vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I 0.00102f
C22944 _312_.ZN a_34586_23208# 0.02581f
C22945 a_66116_4772# a_66204_4728# 0.28563f
C22946 a_47164_13703# a_47612_13703# 0.0131f
C22947 a_64860_3160# a_65308_3160# 0.0131f
C22948 a_67012_3204# a_67100_3160# 0.28563f
C22949 a_64996_14180# a_64972_13703# 0.00172f
C22950 _327_.Z a_40244_18180# 0.52522f
C22951 a_16164_31048# a_16252_29383# 0.0027f
C22952 a_22324_20452# a_22412_20408# 0.28563f
C22953 _452_.CLK _325_.A2 0.15876f
C22954 a_8636_29383# a_9084_29383# 0.0131f
C22955 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I 0.05743f
C22956 _424_.B1 a_50532_24072# 0.00193f
C22957 a_62620_17272# a_62732_16839# 0.02634f
C22958 a_10540_30951# a_11460_31048# 0.00794f
C22959 _457_.D a_24540_24679# 0.01614f
C22960 a_11091_30644# a_10452_31048# 0.00397f
C22961 _452_.CLK a_36524_18407# 0.02666f
C22962 a_11100_1592# VPWR 0.33743f
C22963 a_31260_1592# a_31396_1256# 0.00168f
C22964 _459_.CLK _355_.ZN 0.01934f
C22965 _319_.ZN a_33860_20072# 0.00141f
C22966 a_65332_13800# a_65420_12135# 0.00151f
C22967 a_61612_20408# a_61724_19975# 0.02634f
C22968 _443_.D a_38506_26724# 0.02369f
C22969 a_45508_31048# vgaringosc.workerclkbuff_notouch_.I 0.00646f
C22970 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_63316_23208# 0.00129f
C22971 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN _251_.ZN 0.00665f
C22972 uio_oe[1] uio_oe[0] 0.07417f
C22973 a_46628_11044# a_46716_11000# 0.28563f
C22974 a_32604_19975# VPWR 0.31436f
C22975 _261_.ZN _302_.Z 0.02414f
C22976 a_67996_1159# VPWR 0.35017f
C22977 a_50212_11044# a_50660_11044# 0.01328f
C22978 a_3172_9096# VPWR 0.20993f
C22979 a_5300_5960# VPWR 0.21406f
C22980 _461_.D uo_out[4] 0.00384f
C22981 a_33948_18407# VPWR 0.32378f
C22982 a_8100_1636# a_7964_1159# 0.00168f
C22983 a_4156_1592# a_4156_1159# 0.05841f
C22984 a_35964_1592# a_36412_1592# 0.01288f
C22985 a_33412_16936# a_33860_16936# 0.01328f
C22986 a_62196_23588# a_62284_23544# 0.28563f
C22987 a_17372_30951# uio_oe[0] 0.00741f
C22988 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I 0.00127f
C22989 _304_.B vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.02461f
C22990 a_45484_28248# VPWR 0.3444f
C22991 _419_.Z _424_.ZN 0.00556f
C22992 a_4964_26724# a_4940_26247# 0.00172f
C22993 a_30388_22020# VPWR 0.2267f
C22994 _268_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN 0.10136f
C22995 a_57916_25112# vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN 0.03444f
C22996 _304_.B _384_.A1 0.04373f
C22997 a_44700_30951# a_45148_30951# 0.0131f
C22998 a_1380_12612# VPWR 0.20348f
C22999 _317_.A2 a_34160_20523# 0.00166f
C23000 a_48060_2727# VPWR 0.31143f
C23001 a_35818_29860# VPWR 0.01473f
C23002 vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN a_59172_23208# 0.00656f
C23003 a_932_26344# a_1380_26344# 0.01328f
C23004 a_15244_26247# a_15604_26344# 0.08717f
C23005 _402_.ZN a_46156_25112# 0.06558f
C23006 a_55312_22340# a_55724_22137# 0.00275f
C23007 a_16612_29860# VPWR 0.22899f
C23008 _256_.A2 a_67741_30600# 0.00617f
C23009 _475_.Q a_50212_20452# 0.06801f
C23010 _301_.A1 a_35008_22461# 0.18186f
C23011 a_49292_10567# VPWR 0.32402f
C23012 a_33948_15271# a_34532_15368# 0.01675f
C23013 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I a_59172_23588# 0.00464f
C23014 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN a_62284_23544# 0.0053f
C23015 a_33508_31048# uo_out[5] 0.01703f
C23016 a_31920_29480# a_32308_29167# 0.00393f
C23017 a_1828_23208# VPWR 0.20348f
C23018 _337_.ZN _355_.B 0.03169f
C23019 _369_.ZN _336_.Z 0.00154f
C23020 a_47259_20127# a_47544_20127# 0.00277f
C23021 a_22996_31048# uio_out[3] 0.00331f
C23022 a_2276_28292# a_2724_28292# 0.01328f
C23023 a_932_22020# a_1020_21976# 0.28563f
C23024 a_48060_2727# a_48420_2824# 0.08717f
C23025 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN a_55252_20072# 0.00673f
C23026 a_55340_19975# vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I 0.055f
C23027 _474_.Q _473_.Q 0.43036f
C23028 a_64324_17316# a_64412_17272# 0.28563f
C23029 a_2724_16936# a_2724_15748# 0.05841f
C23030 _371_.A3 _358_.A2 0.00177f
C23031 a_67548_9432# a_67548_8999# 0.05841f
C23032 _371_.ZN a_25124_28776# 0.02499f
C23033 a_36288_31048# VPWR 0.01407f
C23034 a_16052_25156# a_16500_25156# 0.01328f
C23035 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I clk 0.01764f
C23036 _223_.I _362_.ZN 0.00287f
C23037 a_4940_13703# a_4852_13800# 0.28563f
C23038 _304_.B a_41708_30644# 0.07615f
C23039 a_29268_20452# a_29940_20452# 0.00347f
C23040 a_27564_20408# a_28012_20408# 0.0131f
C23041 a_55252_24776# a_55252_23588# 0.05841f
C23042 _416_.A1 _386_.ZN 0.03167f
C23043 a_31260_16839# a_31172_16936# 0.28563f
C23044 a_19140_29612# uio_out[7] 0.00151f
C23045 a_24900_1636# VPWR 0.2085f
C23046 a_38204_1592# a_38340_1256# 0.00168f
C23047 _281_.ZN a_51540_23588# 0.00533f
C23048 _371_.A1 a_28036_26724# 0.02636f
C23049 a_65892_12612# a_65532_12568# 0.08707f
C23050 a_61948_12568# a_62396_12568# 0.01288f
C23051 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN a_59652_25640# 0.1228f
C23052 _404_.A1 _470_.D 0.49055f
C23053 _402_.A1 a_43936_27165# 0.02048f
C23054 _237_.A1 _250_.ZN 0.00589f
C23055 a_52340_12232# a_52428_10567# 0.00151f
C23056 a_43268_1636# a_42908_1592# 0.08707f
C23057 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN VPWR 0.49895f
C23058 _443_.D a_37444_26344# 0.00124f
C23059 a_39548_1159# a_39996_1159# 0.0131f
C23060 _249_.A2 _250_.B 0.39889f
C23061 a_17803_26841# a_18628_26344# 0.0017f
C23062 _324_.C a_42392_19243# 0.006f
C23063 a_15156_20452# VPWR 0.20348f
C23064 a_64772_26344# vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I 0.0016f
C23065 a_5300_27912# a_5388_26247# 0.0027f
C23066 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_63316_23208# 0.00402f
C23067 _384_.A1 VPWR 1.31971f
C23068 a_63988_16936# a_64436_16936# 0.01328f
C23069 a_50300_12568# VPWR 0.34604f
C23070 _284_.ZN a_40196_29480# 0.0069f
C23071 a_43492_15368# a_43940_15368# 0.01328f
C23072 _355_.C _336_.Z 0.64766f
C23073 a_7068_29383# a_6980_29480# 0.28563f
C23074 a_57244_27815# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.00324f
C23075 _452_.CLK a_40244_18180# 0.02739f
C23076 a_3172_10664# VPWR 0.20993f
C23077 a_45372_15271# a_45284_15368# 0.28563f
C23078 a_65756_2727# a_65892_1636# 0.00154f
C23079 a_32740_23208# VPWR 0.20544f
C23080 _230_.I _251_.ZN 0.00349f
C23081 a_46940_15271# a_47388_15271# 0.0131f
C23082 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I 0.03349f
C23083 a_14708_22020# a_14796_21976# 0.28563f
C23084 a_18292_22020# a_18740_22020# 0.01328f
C23085 _424_.A1 _424_.ZN 0.67032f
C23086 a_62172_15704# VPWR 0.30235f
C23087 a_59484_2727# a_59396_2824# 0.28563f
C23088 a_3260_16839# a_3708_16839# 0.0131f
C23089 a_43804_30951# a_43716_31048# 0.28563f
C23090 a_50524_30345# VPWR 0.00111f
C23091 _358_.A3 a_36188_26680# 0.00468f
C23092 _301_.A1 _303_.ZN 0.01968f
C23093 a_36436_16936# a_36548_15748# 0.02666f
C23094 a_28372_23588# a_28012_23544# 0.08674f
C23095 _332_.Z a_41432_17801# 0.00343f
C23096 a_24876_23544# a_25324_23544# 0.0131f
C23097 a_24900_23208# a_24988_21543# 0.00151f
C23098 a_12804_1256# VPWR 0.20348f
C23099 a_27228_26680# VPWR 0.32706f
C23100 a_2364_7864# VPWR 0.30029f
C23101 _417_.A2 a_48964_20204# 0.00673f
C23102 a_41708_30644# VPWR 0.00703f
C23103 a_4156_4728# VPWR 0.30552f
C23104 a_40356_1256# a_40804_1256# 0.01328f
C23105 a_18628_31048# VPWR 0.20947f
C23106 a_55116_13703# a_55476_13800# 0.08707f
C23107 a_1380_13800# a_1828_13800# 0.01328f
C23108 a_3260_29383# VPWR 0.30487f
C23109 a_19388_2727# a_20060_2727# 0.00544f
C23110 _448_.Q _325_.A1 0.56734f
C23111 a_2812_17272# a_2812_16839# 0.05841f
C23112 a_21292_30951# uio_out[5] 0.03726f
C23113 a_41900_16839# a_42484_16936# 0.01675f
C23114 a_62564_29032# _250_.B 0.02012f
C23115 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN a_55788_25112# 0.00311f
C23116 a_57580_10567# a_57604_9476# 0.0016f
C23117 _284_.A2 a_45128_26031# 0.00864f
C23118 a_38564_1636# VPWR 0.20874f
C23119 a_3172_16936# VPWR 0.20993f
C23120 a_19724_23544# a_19612_23111# 0.02634f
C23121 a_6308_1636# a_5948_1592# 0.08707f
C23122 _460_.Q a_35710_28776# 0.00156f
C23123 a_4516_29860# a_4964_29860# 0.01328f
C23124 _476_.Q a_52997_20936# 0.00918f
C23125 _346_.B a_21628_28248# 0.00548f
C23126 a_932_29860# a_1020_29816# 0.28563f
C23127 _316_.A3 VPWR 0.78212f
C23128 a_1916_17272# a_2364_17272# 0.0131f
C23129 a_4516_17316# a_4156_17272# 0.08674f
C23130 _370_.ZN a_29856_29123# 0.02253f
C23131 _330_.A1 _319_.A2 0.20342f
C23132 a_49764_31048# uio_in[1] 0.00485f
C23133 a_56348_11000# a_56796_11000# 0.01288f
C23134 a_60292_11044# a_60380_11000# 0.28563f
C23135 a_57380_16936# a_58164_16936# 0.00276f
C23136 a_49764_1636# a_50212_1636# 0.01328f
C23137 a_58364_25112# VPWR 0.37092f
C23138 _251_.A1 a_56484_29480# 0.00518f
C23139 a_3620_20072# a_3620_18884# 0.05841f
C23140 _419_.A4 a_48172_18840# 0.00111f
C23141 _424_.B1 a_52564_18504# 0.00307f
C23142 a_56684_18407# a_57132_18407# 0.01222f
C23143 a_45820_18407# a_45732_18504# 0.28563f
C23144 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN 0.02197f
C23145 a_47524_18504# a_47500_16839# 0.00131f
C23146 _474_.CLK a_52676_27912# 0.00141f
C23147 _330_.A1 _325_.B 0.00162f
C23148 a_63068_18407# VPWR 0.29679f
C23149 a_64324_18884# a_63964_18840# 0.08717f
C23150 a_1916_25112# VPWR 0.297f
C23151 a_3708_27815# a_4068_27912# 0.08717f
C23152 a_26132_20452# VPWR 0.23408f
C23153 _256_.A2 ui_in[2] 0.03158f
C23154 _346_.ZN a_21424_25987# 0.00107f
C23155 a_64100_12612# VPWR 0.2061f
C23156 a_19744_30301# VPWR 0.19265f
C23157 _447_.Q a_36016_20893# 0.21466f
C23158 a_54780_15704# VPWR 0.32971f
C23159 _325_.A2 a_43668_19668# 0.60936f
C23160 _355_.C uio_out[0] 0.00133f
C23161 a_20420_2824# a_20868_2824# 0.01328f
C23162 _397_.A4 a_47376_27912# 0.00177f
C23163 _272_.B1 _270_.A2 0.00537f
C23164 _311_.A2 a_37108_23588# 0.01288f
C23165 a_37532_25112# a_37556_23588# 0.0012f
C23166 a_56236_24679# clk 0.01994f
C23167 a_53908_24776# a_54356_24776# 0.01328f
C23168 a_64884_10664# VPWR 0.232f
C23169 _355_.B a_27924_24776# 0.00303f
C23170 _371_.A1 a_34348_27208# 0.00181f
C23171 a_65308_8999# a_65220_9096# 0.28563f
C23172 a_67100_5863# a_67012_5960# 0.28563f
C23173 a_56348_15271# a_56708_15368# 0.08717f
C23174 a_58836_17316# vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN 0.005f
C23175 a_66204_7431# a_66116_7528# 0.28563f
C23176 _287_.A2 _223_.I 0.19693f
C23177 a_932_4392# a_932_3204# 0.05841f
C23178 a_14708_21640# a_14708_20452# 0.05841f
C23179 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I 0.0049f
C23180 _355_.C a_23196_24679# 0.00241f
C23181 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I a_58476_18840# 0.00275f
C23182 a_38340_15368# VPWR 0.22423f
C23183 _294_.A2 _459_.CLK 0.96972f
C23184 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I a_62172_18840# 0.00197f
C23185 _395_.A1 _279_.Z 0.0263f
C23186 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I clk 0.05711f
C23187 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN _249_.A2 0.00121f
C23188 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I 0.00407f
C23189 a_53300_23047# _281_.A1 0.00526f
C23190 _350_.A1 _337_.ZN 0.45145f
C23191 a_1916_14136# a_2364_14136# 0.0131f
C23192 a_4516_14180# a_4156_14136# 0.08674f
C23193 a_41564_15271# VPWR 0.36254f
C23194 a_43380_16936# a_43492_15748# 0.02666f
C23195 a_39572_16936# a_39548_15704# 0.0016f
C23196 a_65756_17272# VPWR 0.34838f
C23197 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN 0.00437f
C23198 _474_.CLK _272_.A2 0.02218f
C23199 _324_.C _284_.B 0.14458f
C23200 a_56596_29861# a_57220_29861# 0.00329f
C23201 a_35204_1256# VPWR 0.23527f
C23202 _448_.Q _327_.A2 0.00376f
C23203 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN 0.00319f
C23204 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I 0.66739f
C23205 _218_.ZN a_49896_18909# 0.00202f
C23206 a_66316_13703# a_66228_13800# 0.28563f
C23207 a_34155_25273# a_34440_25273# 0.00277f
C23208 a_18716_30951# VPWR 0.31879f
C23209 a_41488_24072# a_41696_24072# 0.00403f
C23210 a_1380_17316# VPWR 0.20348f
C23211 a_53100_16839# a_53012_16936# 0.28563f
C23212 a_2364_12135# a_2724_12232# 0.08717f
C23213 a_44700_1592# VPWR 0.29679f
C23214 a_11772_1159# a_12356_1256# 0.01675f
C23215 a_56012_12135# a_56460_12135# 0.012f
C23216 a_50324_16936# VPWR 0.25347f
C23217 a_5188_29480# a_5636_29480# 0.01328f
C23218 a_9220_1636# a_9308_1592# 0.28563f
C23219 a_12804_1636# a_13252_1636# 0.01328f
C23220 _452_.CLK a_44162_24120# 0.00144f
C23221 a_64772_26344# VPWR 0.16091f
C23222 a_34308_17316# a_33948_17272# 0.08707f
C23223 _416_.A1 a_39236_26344# 0.00992f
C23224 a_63652_11044# a_63740_11000# 0.28563f
C23225 a_15044_2824# VPWR 0.20348f
C23226 a_39536_26795# a_41099_26841# 0.41635f
C23227 a_60828_26680# a_61836_26680# 0.00323f
C23228 _421_.A1 _381_.A2 0.19141f
C23229 a_58588_21543# VPWR 0.32585f
C23230 a_18716_24679# a_19164_24679# 0.01288f
C23231 a_1020_24679# a_932_24776# 0.28563f
C23232 _459_.CLK a_21424_25987# 0.02736f
C23233 a_60212_25156# clk 0.00618f
C23234 _424_.A2 a_53012_18504# 0.00306f
C23235 _437_.A1 a_39884_27815# 0.01371f
C23236 a_1468_19975# a_1916_19975# 0.0131f
C23237 a_61948_1159# a_62396_1159# 0.0131f
C23238 a_46628_2824# a_46492_1592# 0.00154f
C23239 a_1380_14180# VPWR 0.20348f
C23240 _255_.I vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I 0.01418f
C23241 _455_.Q a_24316_26247# 0.00264f
C23242 a_2812_18407# a_3260_18407# 0.0131f
C23243 a_24080_25227# VPWR 1.10855f
C23244 _304_.B clk 0.03151f
C23245 _416_.A1 _386_.A4 0.02712f
C23246 a_46068_25156# a_46156_25112# 0.28563f
C23247 a_31260_15704# a_31708_15704# 0.01288f
C23248 a_51084_12135# VPWR 0.31389f
C23249 a_18760_29032# VPWR 0.35559f
C23250 a_35204_15748# a_35292_15704# 0.28563f
C23251 a_48868_18504# a_48732_17272# 0.00154f
C23252 a_23196_2727# a_23332_1636# 0.00154f
C23253 _424_.B1 a_51332_24372# 0.44823f
C23254 a_52564_18504# a_52676_17316# 0.02666f
C23255 _397_.A4 a_46198_27060# 0.03764f
C23256 a_45088_29123# _383_.A2 0.00489f
C23257 _427_.A2 a_54088_22895# 0.00369f
C23258 _474_.CLK vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN 0.20427f
C23259 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I 0.00104f
C23260 a_17396_27912# uio_out[7] 0.00187f
C23261 a_4156_24679# VPWR 0.3269f
C23262 a_61612_23111# vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN 0.00334f
C23263 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I 0.00106f
C23264 _452_.CLK a_43824_18147# 0.01643f
C23265 _251_.A1 a_55956_25940# 0.78824f
C23266 a_33860_15748# VPWR 0.20799f
C23267 _447_.Q a_43850_23588# 0.00139f
C23268 a_26468_27912# VPWR 0.2334f
C23269 _384_.ZN a_47636_25940# 0.02511f
C23270 _397_.A4 clkbuf_1_0__f_clk.I 0.07669f
C23271 a_46716_18407# a_47164_18407# 0.0131f
C23272 a_1380_9476# a_1468_9432# 0.28563f
C23273 a_24428_21976# a_24876_21976# 0.01288f
C23274 _452_.CLK a_34716_20937# 0.02606f
C23275 a_28372_22020# a_28460_21976# 0.28563f
C23276 _303_.ZN a_42252_20936# 0.05398f
C23277 _452_.Q a_38971_18559# 0.00455f
C23278 a_50412_16839# a_50860_16839# 0.0131f
C23279 a_48868_14180# a_48508_14136# 0.08707f
C23280 a_4604_25112# a_4516_23588# 0.0027f
C23281 a_46516_16936# a_46492_15704# 0.0016f
C23282 _350_.A2 a_29563_29535# 0.04508f
C23283 a_45260_16839# VPWR 0.29679f
C23284 a_50324_16936# a_50436_15748# 0.02666f
C23285 a_57380_1256# VPWR 0.21508f
C23286 a_62756_1256# a_63204_1256# 0.01328f
C23287 a_22100_31048# uio_out[5] 0.00495f
C23288 _384_.A1 a_51240_23340# 0.46078f
C23289 a_62868_13800# a_63316_13800# 0.01328f
C23290 a_54468_21640# a_54332_20408# 0.00154f
C23291 a_41788_2727# a_42236_2727# 0.0131f
C23292 _270_.A2 VPWR 0.43057f
C23293 a_44812_17272# a_44812_16839# 0.05841f
C23294 _416_.A2 a_47544_20127# 0.00163f
C23295 a_35740_17272# VPWR 0.31547f
C23296 a_35723_20569# _319_.A2 0.03091f
C23297 a_38228_20452# a_38676_20452# 0.01328f
C23298 a_23196_1159# a_23108_1256# 0.28563f
C23299 a_53324_12135# a_53236_12232# 0.28563f
C23300 a_58500_1636# VPWR 0.21417f
C23301 a_15492_29480# _467_.D 0.00135f
C23302 _416_.A1 _407_.A1 0.0062f
C23303 a_10652_29816# a_11100_29816# 0.01288f
C23304 a_14596_29860# a_14684_29816# 0.28563f
C23305 _437_.A1 a_38575_24072# 0.00291f
C23306 _358_.A3 a_34756_24776# 0.00117f
C23307 a_932_26344# a_932_25156# 0.05841f
C23308 a_44724_17316# a_45172_17316# 0.01328f
C23309 a_37444_2824# VPWR 0.20815f
C23310 a_36324_1636# a_36188_1159# 0.00168f
C23311 a_32380_1592# a_32380_1159# 0.05841f
C23312 a_55900_1592# a_56348_1592# 0.01288f
C23313 a_59844_1636# a_59932_1592# 0.28563f
C23314 a_3260_10567# a_3708_10567# 0.0131f
C23315 a_54420_21976# a_54244_20452# 0.00146f
C23316 a_55252_25156# clk 0.00151f
C23317 _248_.B1 a_65756_27815# 0.00544f
C23318 _270_.A2 a_59332_29816# 0.02302f
C23319 _381_.Z _395_.A2 0.00586f
C23320 _459_.CLK a_17844_27912# 0.01229f
C23321 a_29244_23111# a_29692_23111# 0.01288f
C23322 a_20956_24679# a_21316_24776# 0.08707f
C23323 a_17036_23111# a_17396_23208# 0.08717f
C23324 a_4604_9432# VPWR 0.33016f
C23325 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN 0.77848f
C23326 a_50300_14136# VPWR 0.34604f
C23327 _316_.A3 a_36636_21543# 0.00822f
C23328 _317_.A2 a_36548_21640# 0.00173f
C23329 a_53572_2824# a_53436_1592# 0.00154f
C23330 a_2364_21543# a_2812_21543# 0.0131f
C23331 _452_.CLK _302_.Z 0.00128f
C23332 _388_.B a_43916_29816# 0.05208f
C23333 a_33500_18407# a_33412_18504# 0.28563f
C23334 _304_.A1 a_37196_23544# 0.00178f
C23335 _451_.Q _264_.B 0.03579f
C23336 hold2.Z hold2.I 0.30878f
C23337 VPWR clk 5.15414f
C23338 a_64100_27912# vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN 0.03118f
C23339 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I 0.61121f
C23340 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_65756_27815# 0.05077f
C23341 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN 0.19291f
C23342 a_5300_12232# VPWR 0.21406f
C23343 a_37980_15704# a_38652_15704# 0.00544f
C23344 a_42820_2824# a_43268_2824# 0.01328f
C23345 a_51420_15704# a_51556_15368# 0.00168f
C23346 _294_.A2 uo_out[7] 0.06057f
C23347 _470_.D _435_.A3 0.00417f
C23348 _397_.A1 _279_.Z 0.00142f
C23349 a_49740_29383# a_49652_29480# 0.28563f
C23350 _245_.Z a_61052_26247# 0.01932f
C23351 a_1020_20408# a_1020_19975# 0.05841f
C23352 a_17844_24776# VPWR 0.21215f
C23353 a_3260_2727# a_3172_2824# 0.28563f
C23354 a_60604_26247# a_61052_26247# 0.01255f
C23355 a_4940_19975# a_5300_20072# 0.08674f
C23356 a_39996_15704# VPWR 0.3289f
C23357 _459_.CLK _351_.ZN 0.03254f
C23358 a_44864_27165# a_46198_27060# 0.00639f
C23359 a_45820_9432# a_46268_9432# 0.0131f
C23360 a_47972_9476# a_47612_9432# 0.08717f
C23361 a_61276_19975# VPWR 0.3167f
C23362 a_55364_14180# a_55812_14180# 0.01328f
C23363 _294_.ZN _358_.A3 0.04329f
C23364 _350_.A1 a_30795_29977# 0.00853f
C23365 a_18380_25112# a_18292_23588# 0.0027f
C23366 _452_.CLK a_35292_26247# 0.03732f
C23367 _265_.ZN a_43492_27912# 0.00195f
C23368 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I 0.00117f
C23369 a_4068_12612# a_4156_12568# 0.28563f
C23370 a_36660_23588# a_37108_23588# 0.01328f
C23371 a_51868_17272# a_51756_16839# 0.02634f
C23372 _416_.A1 a_45396_28292# 0.01715f
C23373 _393_.ZN _470_.Q 0.00497f
C23374 a_58687_31220# a_60285_30600# 0.00301f
C23375 a_29604_23208# a_29716_22020# 0.02666f
C23376 a_47836_17272# VPWR 0.31389f
C23377 a_25796_23208# a_25772_21976# 0.0016f
C23378 a_67772_1592# VPWR 0.34859f
C23379 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN a_53796_30344# 0.00284f
C23380 a_34172_1159# a_34532_1256# 0.08717f
C23381 a_18940_1592# a_19388_1592# 0.01288f
C23382 a_22884_1636# a_22972_1592# 0.28563f
C23383 a_63852_12135# a_64212_12232# 0.08663f
C23384 a_50100_12232# a_50548_12232# 0.01328f
C23385 a_8100_29860# uio_oe[6] 0.00495f
C23386 a_28348_21543# VPWR 0.31389f
C23387 _441_.A3 _441_.A2 0.18964f
C23388 a_18628_26344# a_18740_25156# 0.02666f
C23389 a_45708_17272# a_46492_17272# 0.00443f
C23390 _459_.CLK _337_.A3 0.351f
C23391 a_40656_23588# VPWR 0.01384f
C23392 VPWR uo_out[0] 0.74161f
C23393 a_64548_1636# a_64636_1592# 0.28563f
C23394 a_59844_2824# VPWR 0.20348f
C23395 a_4068_2824# a_4068_1636# 0.05841f
C23396 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I VPWR 1.08893f
C23397 a_51791_30644# _276_.A2 0.0438f
C23398 _459_.Q _358_.A2 0.2316f
C23399 a_28348_23111# a_28260_23208# 0.28563f
C23400 a_23108_24776# a_23556_24776# 0.01328f
C23401 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I 0.1264f
C23402 a_55228_9432# VPWR 0.31143f
C23403 _452_.Q a_43126_24119# 0.00182f
C23404 _452_.CLK a_46476_20937# 0.00187f
C23405 a_1020_21543# a_1380_21640# 0.08717f
C23406 a_65892_14180# VPWR 0.23142f
C23407 _304_.B hold2.Z 0.026f
C23408 a_51108_21640# a_51240_20452# 0.00168f
C23409 a_44924_15704# a_45372_15704# 0.01288f
C23410 a_66676_12232# VPWR 0.20595f
C23411 _403_.ZN _400_.ZN 0.13677f
C23412 a_60401_30300# a_60793_29860# 0.00762f
C23413 _346_.ZN a_21044_27508# 0.57116f
C23414 a_42728_20452# VPWR 0.01214f
C23415 _365_.ZN a_35204_31048# 0.00398f
C23416 a_61276_19975# a_61188_20072# 0.28563f
C23417 a_35740_30951# a_35652_31048# 0.28563f
C23418 _256_.A2 a_61297_30300# 0.02144f
C23419 a_63964_18840# a_63964_18407# 0.05841f
C23420 _303_.ZN a_42154_21236# 0.03109f
C23421 a_37179_24831# VPWR 0.37286f
C23422 _355_.C a_20308_26724# 0.00158f
C23423 a_4516_18884# VPWR 0.20862f
C23424 _248_.B1 a_63313_28776# 0.0039f
C23425 a_14236_2727# a_14596_2824# 0.08717f
C23426 a_53660_15704# VPWR 0.32517f
C23427 VPWR uio_oe[3] 0.16827f
C23428 a_66540_19975# a_66988_19975# 0.01255f
C23429 a_59260_23544# VPWR 0.31037f
C23430 _324_.C _474_.Q 0.00105f
C23431 a_49180_17272# a_49092_15748# 0.00151f
C23432 a_4516_20452# a_4964_20452# 0.01328f
C23433 a_2724_20452# a_2364_20408# 0.08717f
C23434 a_30388_28776# a_32904_28776# 0.00951f
C23435 _241_.Z VPWR 0.45155f
C23436 _252_.ZN a_59397_26344# 0.07774f
C23437 _350_.A2 VPWR 3.08281f
C23438 _452_.Q a_40636_18180# 0.00101f
C23439 _304_.A1 a_34080_22461# 0.00447f
C23440 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_63313_28776# 0.00155f
C23441 a_52004_12612# a_52452_12612# 0.01328f
C23442 a_64188_2727# a_64636_2727# 0.0131f
C23443 a_48420_12612# a_48508_12568# 0.28563f
C23444 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN a_63404_20408# 0.00343f
C23445 a_32964_20072# a_33412_20072# 0.01328f
C23446 uo_out[1] uo_out[3] 0.12767f
C23447 a_66564_9096# a_66564_7908# 0.05841f
C23448 a_45596_1159# a_45508_1256# 0.28563f
C23449 a_22748_1159# VPWR 0.3289f
C23450 a_64636_12568# a_64548_11044# 0.0027f
C23451 a_67460_7528# a_67460_6340# 0.05841f
C23452 a_26244_1636# a_25884_1592# 0.08707f
C23453 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.00123f
C23454 _229_.I _255_.I 0.1175f
C23455 a_49112_29885# a_50524_30345# 0.00393f
C23456 a_25348_21640# VPWR 0.20721f
C23457 a_52764_17272# a_53212_17272# 0.01288f
C23458 _460_.Q a_35728_29480# 0.01897f
C23459 _424_.B1 a_52408_19759# 0.04023f
C23460 a_47552_19715# a_47612_18407# 0.00101f
C23461 a_51084_10567# a_51444_10664# 0.08707f
C23462 a_64972_10567# a_65420_10567# 0.0131f
C23463 a_5724_1159# a_6172_1159# 0.0131f
C23464 _325_.A2 a_40668_19975# 0.00839f
C23465 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I 0.66813f
C23466 a_66787_30600# VPWR 0.31557f
C23467 a_64212_23208# VPWR 0.21036f
C23468 a_26916_23208# a_27364_23208# 0.01328f
C23469 _424_.B1 a_51668_23340# 0.00558f
C23470 _437_.A1 _452_.CLK 0.06853f
C23471 a_33612_24679# a_33524_24776# 0.28563f
C23472 a_66204_9432# VPWR 0.31657f
C23473 a_15244_23544# VPWR 0.29679f
C23474 a_21404_21543# a_21316_21640# 0.28563f
C23475 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN 0.00118f
C23476 a_33276_21543# a_33724_21543# 0.012f
C23477 a_2812_2727# VPWR 0.30213f
C23478 a_35652_2824# a_35740_1159# 0.0027f
C23479 a_1020_5863# VPWR 0.30073f
C23480 _459_.CLK a_21044_27508# 0.0278f
C23481 a_52876_13703# VPWR 0.33058f
C23482 hold2.Z VPWR 0.74854f
C23483 _337_.A3 _371_.A3 0.0222f
C23484 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.05101f
C23485 _351_.A2 a_25300_26344# 0.01994f
C23486 _416_.A3 VPWR 0.93106f
C23487 a_15132_29816# a_15132_29383# 0.05841f
C23488 a_52228_15748# a_51868_15704# 0.08707f
C23489 a_48060_11000# VPWR 0.29679f
C23490 _243_.A1 _243_.ZN 0.54909f
C23491 a_64996_2824# a_65668_2824# 0.00347f
C23492 a_31516_28292# VPWR 0.00866f
C23493 a_3620_26724# VPWR 0.22347f
C23494 a_15460_31048# a_15492_29860# 0.02587f
C23495 _223_.I a_31031_27208# 0.00775f
C23496 _281_.A1 _474_.D 0.00209f
C23497 a_63616_31128# a_64996_31048# 0.00977f
C23498 _304_.ZN a_43380_20452# 0.01859f
C23499 a_62532_15748# a_62980_15748# 0.01328f
C23500 _447_.Q _325_.A2 0.01151f
C23501 a_30924_20408# a_30812_19975# 0.02634f
C23502 a_32628_20452# a_32604_19975# 0.00172f
C23503 _399_.ZN a_46356_24072# 0.50217f
C23504 _300_.A2 _323_.A3 0.01672f
C23505 a_47612_30951# vgaringosc.workerclkbuff_notouch_.I 0.00613f
C23506 a_15604_26344# VPWR 0.20348f
C23507 a_58948_26344# VPWR 0.20618f
C23508 a_25660_2727# a_25572_2824# 0.28563f
C23509 _251_.A1 a_64412_29816# 0.0065f
C23510 _245_.Z a_60516_26344# 0.01464f
C23511 a_29716_31048# a_29232_29931# 0.00263f
C23512 a_3260_28248# VPWR 0.30487f
C23513 a_56796_9432# a_57244_9432# 0.0131f
C23514 a_58948_9476# a_58588_9432# 0.08717f
C23515 a_48104_30219# _383_.A2 0.00398f
C23516 a_1828_23588# a_2276_23588# 0.01328f
C23517 a_6532_1256# a_6980_1256# 0.01328f
C23518 a_60604_26247# a_60516_26344# 0.28563f
C23519 _365_.ZN _296_.ZN 0.00429f
C23520 _260_.A2 a_44500_22020# 0.0037f
C23521 a_30476_21976# a_30388_20452# 0.00151f
C23522 a_1828_6340# a_2276_6340# 0.01328f
C23523 a_2724_4772# a_3172_4772# 0.01328f
C23524 a_63740_14136# a_64188_14136# 0.01288f
C23525 a_67684_14180# a_67324_14136# 0.08707f
C23526 a_3620_3204# a_4068_3204# 0.01328f
C23527 a_1828_3204# a_1468_3160# 0.08717f
C23528 a_50084_24328# a_50464_24908# 0.00217f
C23529 a_34715_22137# _317_.A2 0.00102f
C23530 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I 0.00361f
C23531 a_55252_23588# a_55340_23544# 0.28563f
C23532 _237_.A1 _230_.I 0.01207f
C23533 a_4516_1636# VPWR 0.20812f
C23534 a_54132_13800# a_54220_12135# 0.00151f
C23535 vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I VPWR 0.72465f
C23536 a_6396_29816# a_6532_29480# 0.00168f
C23537 _459_.CLK _342_.ZN 0.14242f
C23538 a_45148_1159# VPWR 0.29679f
C23539 a_16164_31048# uio_oe[0] 0.00622f
C23540 a_56572_1159# a_56932_1256# 0.08717f
C23541 a_62980_18884# VPWR 0.20348f
C23542 a_32740_1636# a_33188_1636# 0.01328f
C23543 a_2276_11044# a_1916_11000# 0.08717f
C23544 a_4068_11044# a_4516_11044# 0.01328f
C23545 a_64524_16839# a_64972_16839# 0.01222f
C23546 a_49068_20408# a_50212_20452# 0.00869f
C23547 _452_.CLK a_32180_23588# 0.00382f
C23548 a_42684_27815# a_43132_27815# 0.01255f
C23549 _373_.ZN a_28000_29480# 0.26027f
C23550 _467_.D a_17036_27815# 0.01471f
C23551 a_62060_10567# a_61972_10664# 0.28563f
C23552 _459_.CLK a_40644_29480# 0.00226f
C23553 a_20003_29611# _378_.I 0.01616f
C23554 a_16140_21976# VPWR 0.29679f
C23555 _242_.Z vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.05059f
C23556 _424_.A2 a_51892_23340# 0.00118f
C23557 _252_.B a_60516_26344# 0.00738f
C23558 _324_.C _395_.A2 0.15744f
C23559 _243_.A1 a_58140_26680# 0.00275f
C23560 a_29804_23544# VPWR 0.34412f
C23561 a_31932_21543# a_32292_21640# 0.08707f
C23562 a_25212_2727# VPWR 0.31144f
C23563 a_46628_13800# VPWR 0.20348f
C23564 _330_.A1 a_40416_18885# 0.00722f
C23565 a_2364_29816# VPWR 0.30029f
C23566 a_61860_11044# VPWR 0.20595f
C23567 _431_.A3 a_39236_26344# 0.07477f
C23568 a_20532_22020# a_20508_21543# 0.00172f
C23569 a_16588_21976# a_16588_21543# 0.05841f
C23570 a_51420_2727# a_51556_1636# 0.00154f
C23571 a_3708_23111# VPWR 0.33374f
C23572 a_4068_27912# VPWR 0.22146f
C23573 a_50120_26476# a_50792_26344# 0.00488f
C23574 hold2.I _448_.Q 0.01022f
C23575 a_36636_2727# a_36996_2824# 0.08717f
C23576 a_63852_23111# a_64212_23208# 0.08717f
C23577 uio_out[2] uio_out[1] 0.0708f
C23578 _327_.A2 a_41664_22020# 0.01553f
C23579 _384_.ZN _475_.Q 0.15749f
C23580 _427_.B1 a_53548_24679# 0.0087f
C23581 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN a_53124_27912# 0.00134f
C23582 a_1020_7864# a_1020_7431# 0.05841f
C23583 a_2812_4728# a_2812_4295# 0.05841f
C23584 a_66116_4772# a_65756_4728# 0.08717f
C23585 _327_.Z a_39264_18147# 0.00197f
C23586 a_65220_6340# a_64860_6296# 0.08717f
C23587 a_1916_6296# a_1916_5863# 0.05841f
C23588 a_62084_20072# a_62084_18884# 0.05841f
C23589 _264_.B a_42161_24776# 0.26809f
C23590 a_61052_14136# a_61164_13703# 0.02634f
C23591 a_3708_3160# a_3708_2727# 0.05841f
C23592 a_67012_3204# a_66652_3160# 0.08717f
C23593 a_21740_20408# a_22412_20408# 0.00544f
C23594 a_23668_20452# a_24116_20452# 0.01328f
C23595 a_10540_30951# a_10452_31048# 0.28563f
C23596 _452_.CLK a_34732_19975# 0.00487f
C23597 _452_.CLK a_36076_18407# 0.00971f
C23598 a_66564_17316# a_66540_16839# 0.00172f
C23599 a_58140_12568# a_58588_12568# 0.01288f
C23600 a_10652_1592# VPWR 0.33458f
C23601 _459_.CLK a_27328_25227# 0.11581f
C23602 a_67436_19975# a_67460_18884# 0.0016f
C23603 _334_.A1 VPWR 2.88913f
C23604 a_45060_31048# vgaringosc.workerclkbuff_notouch_.I 0.00649f
C23605 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_62868_23208# 0.00245f
C23606 a_67548_1159# VPWR 0.3289f
C23607 a_67996_1159# a_67908_1256# 0.28563f
C23608 a_2724_9096# VPWR 0.20782f
C23609 a_32156_19975# VPWR 0.31436f
C23610 a_62196_23588# a_61836_23544# 0.08674f
C23611 a_4852_5960# VPWR 0.22733f
C23612 a_39460_1636# a_40132_1636# 0.00347f
C23613 a_46628_11044# a_46268_11000# 0.08707f
C23614 _452_.CLK a_32180_22020# 0.0092f
C23615 a_33500_18407# VPWR 0.30042f
C23616 _268_.A1 _267_.A2 0.2278f
C23617 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I 0.00472f
C23618 a_54332_20408# a_54356_20072# 0.00172f
C23619 a_16916_31048# uio_oe[0] 0.0965f
C23620 a_58836_10664# a_59284_10664# 0.01328f
C23621 _457_.D VPWR 0.43964f
C23622 a_28124_1159# a_28572_1159# 0.0131f
C23623 a_20868_24776# a_20956_23111# 0.00151f
C23624 a_45036_28248# VPWR 0.3147f
C23625 a_29804_21976# VPWR 0.34427f
C23626 a_2364_26680# a_2364_26247# 0.05841f
C23627 _454_.Q VPWR 1.64933f
C23628 _268_.A1 a_53212_29816# 0.12654f
C23629 _311_.Z _316_.A3 0.40082f
C23630 a_30500_21640# a_30948_21640# 0.01328f
C23631 _304_.B a_52660_24072# 0.00114f
C23632 a_35156_29860# VPWR 0.01725f
C23633 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I 0.00286f
C23634 a_47612_2727# VPWR 0.31143f
C23635 a_932_12612# VPWR 0.22176f
C23636 a_15244_26247# a_15156_26344# 0.28563f
C23637 a_4604_3160# a_4516_1636# 0.0027f
C23638 a_32068_15368# a_32516_15368# 0.01328f
C23639 uio_out[5] uio_out[6] 0.55838f
C23640 _441_.A2 _226_.ZN 0.03021f
C23641 _459_.Q _294_.A2 0.28498f
C23642 _402_.ZN a_46068_25156# 0.04814f
C23643 a_16028_29816# VPWR 0.35704f
C23644 _475_.Q a_49068_20408# 0.13171f
C23645 _256_.A2 a_67117_30600# 0.03309f
C23646 a_48508_10567# VPWR 0.31817f
C23647 a_23532_21976# a_23644_21543# 0.02634f
C23648 a_33948_15271# a_33860_15368# 0.28563f
C23649 a_27476_22020# a_27452_21543# 0.00172f
C23650 _474_.Q _281_.A1 0.52332f
C23651 a_1380_23208# VPWR 0.20348f
C23652 a_33060_31048# uo_out[5] 0.01725f
C23653 a_49764_26724# a_50176_26724# 0.00217f
C23654 _268_.A2 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN 0.00567f
C23655 a_35516_15271# a_35964_15271# 0.0131f
C23656 _304_.B _448_.Q 0.46401f
C23657 a_22548_31048# uio_out[3] 0.00127f
C23658 _346_.B a_21740_29383# 0.00542f
C23659 a_62644_26724# a_63092_26724# 0.01328f
C23660 _363_.Z _362_.ZN 1.09589f
C23661 a_2724_22020# a_3172_22020# 0.01328f
C23662 a_48060_2727# a_47972_2824# 0.28563f
C23663 a_33483_29535# a_33776_29123# 0.49241f
C23664 a_64324_17316# a_63964_17272# 0.08717f
C23665 a_55340_19975# a_55252_20072# 0.28563f
C23666 a_53300_23047# a_53696_22895# 0.00232f
C23667 a_53436_18840# a_53460_18504# 0.00172f
C23668 a_4852_23208# a_4940_21543# 0.00151f
C23669 a_20172_23544# a_20620_23544# 0.01288f
C23670 a_28932_1256# a_29380_1256# 0.01328f
C23671 _441_.A2 _300_.ZN 0.101f
C23672 a_4156_8999# a_4940_8999# 0.00443f
C23673 a_35652_31048# VPWR 0.2071f
C23674 _230_.I _242_.Z 0.01677f
C23675 _284_.ZN _330_.A1 0.03158f
C23676 a_65756_4295# a_66204_4295# 0.0131f
C23677 a_64860_5863# a_65308_5863# 0.0131f
C23678 a_41056_30669# a_41708_30644# 0.00587f
C23679 a_15132_29383# uio_oe[1] 0.00134f
C23680 a_4156_13703# a_4852_13800# 0.01227f
C23681 a_58028_13703# a_58476_13703# 0.01288f
C23682 _355_.C a_28000_29480# 0.05269f
C23683 a_7964_2727# a_8636_2727# 0.00544f
C23684 a_29268_20452# a_29356_20408# 0.28563f
C23685 a_40020_16936# a_40220_15271# 0.00119f
C23686 a_30812_16839# a_31172_16936# 0.08717f
C23687 _402_.B a_46580_23588# 0.01771f
C23688 a_18264_29480# uio_out[7] 0.04166f
C23689 a_49652_29480# VPWR 0.22058f
C23690 a_24452_1636# VPWR 0.22925f
C23691 a_65444_12612# a_65532_12568# 0.28563f
C23692 a_11548_30951# a_12548_31048# 0.00223f
C23693 a_3260_23544# a_3260_23111# 0.05841f
C23694 _371_.A1 a_27588_26724# 0.00321f
C23695 _230_.I a_63105_28293# 0.02342f
C23696 _304_.B a_41140_27912# 0.0152f
C23697 a_62532_18504# a_62980_18504# 0.01328f
C23698 _404_.A1 a_44961_27912# 0.0663f
C23699 _402_.A1 a_43008_26795# 0.05282f
C23700 _365_.ZN _335_.ZN 0.04933f
C23701 a_54780_20408# a_54892_19975# 0.02634f
C23702 a_1380_15368# a_1380_14180# 0.05841f
C23703 a_53124_11044# a_53572_11044# 0.01328f
C23704 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I a_67124_20452# 0.03006f
C23705 a_44276_16936# a_44724_16936# 0.01328f
C23706 a_42820_1636# a_42908_1592# 0.28563f
C23707 a_46404_1636# a_46852_1636# 0.01328f
C23708 a_4156_26680# a_4604_26680# 0.01222f
C23709 a_32292_2824# a_32292_1636# 0.05841f
C23710 _249_.A2 a_63952_29480# 0.14972f
C23711 _350_.A2 _370_.B 0.81891f
C23712 _362_.B _358_.A3 0.06563f
C23713 a_14708_20452# VPWR 0.22176f
C23714 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN a_62868_23208# 0.00198f
C23715 a_49852_12568# VPWR 0.32315f
C23716 a_8996_2824# a_9444_2824# 0.01328f
C23717 _284_.ZN a_39748_29480# 0.00433f
C23718 a_6620_29383# a_6980_29480# 0.08717f
C23719 a_56124_27815# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.00507f
C23720 _452_.CLK a_39264_18147# 0.03084f
C23721 a_3260_28248# a_3260_27815# 0.05841f
C23722 _416_.A1 _424_.A2 1.05826f
C23723 a_2724_10664# VPWR 0.20782f
C23724 a_33152_22091# a_33276_21543# 0.00156f
C23725 a_44924_15271# a_45284_15368# 0.08717f
C23726 a_32292_23208# VPWR 0.20622f
C23727 _324_.C _427_.A2 0.31512f
C23728 a_35140_26680# a_36100_26724# 0.06083f
C23729 _384_.A3 _395_.A3 0.07606f
C23730 _448_.Q VPWR 2.59662f
C23731 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I a_58924_17272# 0.00653f
C23732 a_16500_28292# a_16588_28248# 0.28563f
C23733 a_15244_28248# a_15692_28248# 0.01255f
C23734 a_59036_2727# a_59396_2824# 0.08717f
C23735 a_67908_15748# VPWR 0.21197f
C23736 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN _249_.A2 0.29104f
C23737 _459_.Q a_32268_23544# 0.00111f
C23738 a_62532_15368# a_62980_15368# 0.01328f
C23739 a_43356_30951# a_43716_31048# 0.08717f
C23740 _245_.I1 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I 0.02971f
C23741 _358_.A3 a_32628_26725# 0.14158f
C23742 _332_.Z a_41536_17636# 0.00311f
C23743 a_12356_1256# VPWR 0.22423f
C23744 a_1916_7864# VPWR 0.297f
C23745 a_27924_23588# a_28012_23544# 0.28563f
C23746 a_18828_25112# a_19276_25112# 0.01288f
C23747 a_23284_26724# VPWR 0.00667f
C23748 a_18180_31048# VPWR 0.21194f
C23749 a_3708_4728# VPWR 0.33374f
C23750 a_32604_18840# a_32604_18407# 0.05841f
C23751 a_2812_29383# VPWR 0.30213f
C23752 a_53300_23047# a_53704_23219# 0.41635f
C23753 a_55116_13703# a_55028_13800# 0.28563f
C23754 a_51220_16936# a_51196_15271# 0.00134f
C23755 a_20250_31048# uio_out[5] 0.00295f
C23756 _370_.B a_31516_28292# 0.00113f
C23757 a_4964_17316# a_4940_16839# 0.00172f
C23758 a_41900_16839# a_41812_16936# 0.28563f
C23759 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I 0.04967f
C23760 a_55700_25156# a_55788_25112# 0.28563f
C23761 a_2724_16936# VPWR 0.20782f
C23762 a_38116_1636# VPWR 0.2085f
C23763 a_41140_27912# VPWR 0.2124f
C23764 a_1916_1592# a_2364_1592# 0.01288f
C23765 a_5860_1636# a_5948_1592# 0.28563f
C23766 _460_.Q a_35516_28776# 0.00235f
C23767 _395_.A2 _281_.A1 0.01624f
C23768 a_55676_28248# a_55676_27815# 0.05841f
C23769 a_4068_17316# a_4156_17272# 0.28563f
C23770 _370_.ZN a_29563_29535# 0.05282f
C23771 a_49316_31048# uio_in[1] 0.00158f
C23772 a_62868_12232# a_62956_10567# 0.00151f
C23773 a_60292_11044# a_59932_11000# 0.08663f
C23774 a_21988_1636# a_21852_1159# 0.00168f
C23775 a_18044_1592# a_18044_1159# 0.05841f
C23776 a_57916_25112# VPWR 0.32207f
C23777 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I 0.64208f
C23778 a_61388_15704# a_61412_14180# 0.00131f
C23779 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN a_54892_18407# 0.00223f
C23780 a_44752_18147# a_45732_18504# 0.00702f
C23781 a_50524_1159# a_50972_1159# 0.0131f
C23782 _397_.A4 _408_.ZN 0.1062f
C23783 a_63876_18884# a_63964_18840# 0.28563f
C23784 a_62620_18407# VPWR 0.29679f
C23785 _478_.D a_52852_24372# 0.5718f
C23786 a_1468_25112# VPWR 0.29679f
C23787 a_3708_27815# a_3620_27912# 0.28563f
C23788 a_56596_18504# a_56596_17316# 0.05841f
C23789 a_25548_20408# VPWR 0.3429f
C23790 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN a_62564_29032# 0.05207f
C23791 a_18816_29931# VPWR 1.12792f
C23792 _399_.A2 a_48529_22460# 0.0039f
C23793 a_2812_15704# a_3260_15704# 0.0131f
C23794 a_63652_12612# VPWR 0.20595f
C23795 a_37084_15704# a_37220_15368# 0.00168f
C23796 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.30331f
C23797 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I a_66452_20072# 0.00119f
C23798 a_54332_15704# VPWR 0.33433f
C23799 _247_.B VPWR 0.24972f
C23800 a_54468_15368# a_54916_15368# 0.01328f
C23801 a_39012_15748# a_38876_15271# 0.00168f
C23802 a_67772_24679# a_67684_24776# 0.28563f
C23803 _311_.A2 a_36660_23588# 0.01496f
C23804 a_55788_24679# clk 0.01871f
C23805 a_56348_15271# a_56260_15368# 0.28563f
C23806 a_64212_10664# VPWR 0.21386f
C23807 a_31820_21976# a_31844_21640# 0.00172f
C23808 a_64860_8999# a_65220_9096# 0.08717f
C23809 a_65756_7431# a_66116_7528# 0.08717f
C23810 _371_.A1 a_33940_27208# 0.00811f
C23811 a_66652_5863# a_67012_5960# 0.08717f
C23812 a_23196_21543# a_23220_20452# 0.0016f
C23813 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN 0.02711f
C23814 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN 0.62895f
C23815 a_37668_15368# VPWR 0.20968f
C23816 a_21068_21976# a_21516_21976# 0.01288f
C23817 a_41116_15271# VPWR 0.33252f
C23818 a_39212_16839# a_39660_16839# 0.01288f
C23819 hold2.Z _260_.ZN 0.46425f
C23820 a_4068_14180# a_4156_14136# 0.28563f
C23821 a_28460_23544# a_28372_22020# 0.00151f
C23822 a_65308_17272# VPWR 0.32087f
C23823 a_51332_1256# a_51780_1256# 0.01328f
C23824 _435_.ZN _441_.B 0.01703f
C23825 _390_.ZN a_51048_26680# 0.007f
C23826 a_34532_1256# VPWR 0.21829f
C23827 _448_.Q a_40452_22504# 0.00237f
C23828 a_30364_2727# a_30812_2727# 0.0131f
C23829 a_65868_13703# a_66228_13800# 0.08717f
C23830 a_49740_13703# a_49764_12612# 0.0016f
C23831 a_51892_13800# a_52340_13800# 0.01328f
C23832 a_34844_17272# a_34732_16839# 0.02634f
C23833 a_56596_17316# a_57044_17316# 0.01328f
C23834 a_18268_30951# VPWR 0.31633f
C23835 _451_.Q a_41564_24679# 0.00142f
C23836 _241_.Z a_57156_27912# 0.00654f
C23837 a_62532_30736# ui_in[1] 0.56401f
C23838 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I a_55140_28292# 0.04608f
C23839 a_4852_23208# a_4964_22020# 0.02666f
C23840 a_52652_16839# a_53012_16936# 0.08717f
C23841 a_932_17316# VPWR 0.22176f
C23842 a_44252_1592# VPWR 0.29679f
C23843 a_44632_30206# a_45416_29885# 0.02307f
C23844 a_11772_1159# a_11684_1256# 0.28563f
C23845 a_52092_1592# a_52228_1256# 0.00168f
C23846 a_49652_16936# VPWR 0.21819f
C23847 a_55924_10664# a_56036_9476# 0.02666f
C23848 _452_.CLK a_43750_23544# 0.00146f
C23849 a_9220_1636# a_8860_1592# 0.08707f
C23850 a_2364_12135# a_2276_12232# 0.28563f
C23851 a_27116_23544# a_27004_23111# 0.02634f
C23852 _447_.Q _302_.Z 0.79804f
C23853 _411_.A2 _412_.B2 0.31525f
C23854 a_7292_29816# a_7740_29816# 0.01288f
C23855 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I a_67772_21543# 0.02166f
C23856 a_33860_17316# a_33948_17272# 0.28563f
C23857 a_37444_17316# a_37892_17316# 0.01328f
C23858 a_66788_11044# a_67236_11044# 0.01328f
C23859 a_63652_11044# a_63292_11000# 0.08707f
C23860 _330_.A1 a_39772_26247# 0.00163f
C23861 a_14596_2824# VPWR 0.20348f
C23862 _442_.ZN a_40092_27209# 0.21751f
C23863 a_39536_26795# a_41392_27165# 0.02307f
C23864 _250_.ZN a_62503_28293# 0.07669f
C23865 a_52540_1592# a_52988_1592# 0.01288f
C23866 _451_.Q _325_.A2 0.32021f
C23867 _398_.C _417_.A2 0.00221f
C23868 a_37532_26680# VPWR 0.31901f
C23869 a_17932_23111# a_18716_23111# 0.00443f
C23870 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.00704f
C23871 _437_.A1 a_38816_27555# 0.22432f
C23872 _424_.A2 a_52564_18504# 0.00228f
C23873 _459_.CLK a_20496_26344# 0.09805f
C23874 _455_.Q a_23868_26247# 0.00225f
C23875 _300_.A2 a_38784_22504# 0.00265f
C23876 a_4604_7864# a_4516_6340# 0.0027f
C23877 _397_.A4 _412_.A1 0.11922f
C23878 a_932_14180# VPWR 0.22176f
C23879 _474_.CLK _267_.A2 0.07571f
C23880 a_19412_27912# a_19860_27912# 0.01328f
C23881 _459_.CLK a_16500_28292# 0.00434f
C23882 _334_.A1 _370_.B 0.59497f
C23883 a_50636_12135# VPWR 0.33727f
C23884 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I 0.092f
C23885 a_35204_15748# a_34844_15704# 0.08707f
C23886 a_31396_2824# a_31844_2824# 0.01328f
C23887 _427_.A2 a_54192_22851# 0.0035f
C23888 _474_.CLK a_53212_29816# 0.05954f
C23889 a_3708_24679# VPWR 0.33374f
C23890 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_62420_22020# 0.07299f
C23891 _452_.CLK a_42896_18504# 0.08446f
C23892 a_21764_21640# a_21740_20408# 0.0016f
C23893 a_33412_15748# VPWR 0.20644f
C23894 _419_.A4 a_47689_25156# 0.00215f
C23895 _267_.A1 a_52756_29076# 0.00158f
C23896 a_43380_20452# _328_.A2 0.00152f
C23897 a_1380_9476# a_1020_9432# 0.08717f
C23898 a_3172_9476# a_3620_9476# 0.01328f
C23899 a_28372_22020# a_28012_21976# 0.08707f
C23900 _452_.CLK a_35088_20893# 0.04293f
C23901 a_48420_14180# a_48508_14136# 0.28563f
C23902 a_52004_14180# a_52452_14180# 0.01328f
C23903 _452_.CLK a_37532_17272# 0.00613f
C23904 a_44812_16839# VPWR 0.29679f
C23905 _350_.A2 a_28556_29167# 0.00188f
C23906 _248_.B1 clk 0.02967f
C23907 a_21652_31048# uio_out[5] 0.00935f
C23908 a_52848_25987# a_52744_26031# 0.10745f
C23909 _325_.A1 _450_.D 0.25406f
C23910 a_56932_1256# VPWR 0.20704f
C23911 a_52452_24072# a_52920_22760# 0.01248f
C23912 a_46628_13800# a_46628_12612# 0.05841f
C23913 a_66428_14136# a_66340_12612# 0.00151f
C23914 _359_.B uo_out[2] 0.04564f
C23915 a_59143_31198# VPWR 0.00423f
C23916 a_35292_17272# VPWR 0.32253f
C23917 a_36016_20893# _319_.A2 0.02333f
C23918 a_58052_1636# VPWR 0.2247f
C23919 a_22748_1159# a_23108_1256# 0.08717f
C23920 a_61524_10664# a_61500_9432# 0.0016f
C23921 a_63316_10664# a_63204_9476# 0.02666f
C23922 a_16164_29480# a_16612_29480# 0.01328f
C23923 a_66764_12135# a_67212_12135# 0.0131f
C23924 _402_.A1 _282_.ZN 0.00817f
C23925 a_52876_12135# a_53236_12232# 0.08707f
C23926 a_15580_1592# a_16028_1592# 0.012f
C23927 a_25772_23544# a_25796_23208# 0.00172f
C23928 _325_.B a_43452_18191# 0.00739f
C23929 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN clk 0.01941f
C23930 a_63952_29480# _250_.B 0.12839f
C23931 a_14596_29860# a_14236_29816# 0.08707f
C23932 _412_.A1 a_51956_26183# 0.01905f
C23933 a_40040_17675# a_41048_17341# 0.02307f
C23934 _358_.A3 a_34308_24776# 0.00158f
C23935 a_41056_30669# uo_out[0] 0.17054f
C23936 a_59844_1636# a_59484_1592# 0.08707f
C23937 _370_.ZN VPWR 0.29474f
C23938 a_36996_2824# VPWR 0.20815f
C23939 a_54804_25156# clk 0.00151f
C23940 _270_.A2 a_58116_30344# 0.49961f
C23941 _459_.CLK a_17396_27912# 0.03533f
C23942 a_17036_23111# a_16948_23208# 0.28563f
C23943 a_20956_24679# a_20868_24776# 0.28563f
C23944 a_2724_24776# a_3172_24776# 0.01328f
C23945 a_66564_9096# a_67012_9096# 0.01328f
C23946 _316_.A3 a_35816_21192# 0.01317f
C23947 a_4156_9432# VPWR 0.30552f
C23948 a_49852_14136# VPWR 0.32315f
C23949 a_55956_25940# vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN 0.00186f
C23950 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_55700_25156# 0.00628f
C23951 _400_.ZN _421_.A1 0.03977f
C23952 a_2276_18504# a_2724_18504# 0.01328f
C23953 _427_.A2 _281_.A1 0.05526f
C23954 a_33052_18407# a_33412_18504# 0.08717f
C23955 _304_.A1 a_36748_23544# 0.00672f
C23956 a_18044_29816# uio_out[7] 0.01475f
C23957 _281_.A1 a_51196_21543# 0.00736f
C23958 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN a_64188_27815# 0.02457f
C23959 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62844_27815# 0.00502f
C23960 a_4852_12232# VPWR 0.22733f
C23961 a_41700_15748# a_42148_15748# 0.01328f
C23962 _441_.ZN _441_.B 0.2587f
C23963 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_61836_23544# 0.00163f
C23964 a_36656_29123# uo_out[2] 0.00155f
C23965 _424_.A2 a_51332_24372# 0.34445f
C23966 _397_.A1 a_47297_25596# 0.00976f
C23967 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN _250_.B 0.32741f
C23968 a_17396_24776# VPWR 0.20348f
C23969 _244_.Z _251_.ZN 0.00544f
C23970 _245_.Z a_60604_26247# 0.01703f
C23971 _340_.A2 _342_.ZN 0.31134f
C23972 a_2812_2727# a_3172_2824# 0.08717f
C23973 a_39548_15704# VPWR 0.3289f
C23974 a_4940_19975# a_4852_20072# 0.28563f
C23975 _459_.CLK a_24304_26795# 0.01392f
C23976 _359_.B a_43916_29816# 0.00584f
C23977 a_47524_9476# a_47612_9432# 0.28563f
C23978 _451_.Q a_40244_18180# 0.28766f
C23979 _294_.ZN a_31484_26680# 0.00487f
C23980 _350_.A1 a_31088_30301# 0.01207f
C23981 _327_.A2 _450_.D 0.08215f
C23982 _444_.D a_37556_23588# 0.00285f
C23983 _265_.ZN a_43044_27912# 0.0053f
C23984 a_52764_2727# a_53212_2727# 0.0131f
C23985 a_53684_13800# a_53572_12612# 0.02666f
C23986 a_1468_12568# a_1916_12568# 0.0131f
C23987 a_4068_12612# a_3708_12568# 0.08717f
C23988 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I 0.79495f
C23989 _416_.A1 a_44948_28292# 0.10246f
C23990 a_47388_17272# VPWR 0.31389f
C23991 a_67324_1592# VPWR 0.3289f
C23992 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN a_53592_30344# 0.00174f
C23993 _437_.A1 _447_.Q 0.07693f
C23994 a_34172_1159# a_34084_1256# 0.28563f
C23995 a_67772_1592# a_67908_1256# 0.00168f
C23996 a_63852_12135# a_63764_12232# 0.28563f
C23997 _252_.B _245_.Z 0.55533f
C23998 _324_.C a_59572_29076# 0.00812f
C23999 a_1828_4392# a_1828_3204# 0.05841f
C24000 _378_.I a_21287_29076# 0.00433f
C24001 a_22884_1636# a_22524_1592# 0.08707f
C24002 a_22560_30288# a_23108_29860# 0.19548f
C24003 _287_.A1 a_36500_29860# 0.01106f
C24004 _311_.A2 a_36860_23111# 0.0069f
C24005 a_27900_21543# VPWR 0.31389f
C24006 _304_.B _234_.ZN 0.02577f
C24007 a_49540_17316# a_49988_17316# 0.01328f
C24008 _284_.A2 hold2.I 0.00516f
C24009 a_40452_23588# VPWR 0.0068f
C24010 a_59396_2824# VPWR 0.20348f
C24011 a_67772_11000# a_67660_10567# 0.02634f
C24012 a_53772_10567# a_54220_10567# 0.01288f
C24013 a_66340_1636# a_66788_1636# 0.01328f
C24014 a_64548_1636# a_64188_1592# 0.08717f
C24015 a_15604_23208# a_16052_23208# 0.01328f
C24016 _459_.Q a_29828_26344# 0.01102f
C24017 a_27900_23111# a_28260_23208# 0.08707f
C24018 a_60793_29860# VPWR 0.00574f
C24019 _452_.Q a_42796_23981# 0.00189f
C24020 a_54780_9432# VPWR 0.31143f
C24021 VPWR uio_out[1] 0.40442f
C24022 _399_.ZN a_47948_23111# 0.02717f
C24023 a_24228_2824# a_24316_1159# 0.0027f
C24024 a_65444_14180# VPWR 0.21032f
C24025 a_22300_21543# a_22748_21543# 0.01288f
C24026 a_1020_21543# a_932_21640# 0.28563f
C24027 _330_.A1 _331_.ZN 0.29936f
C24028 _336_.A1 a_28796_23111# 0.02761f
C24029 _304_.B a_41476_26344# 0.06203f
C24030 _324_.C a_44571_26841# 0.01363f
C24031 _384_.A3 _427_.B1 0.00975f
C24032 _230_.I a_60156_27815# 0.01875f
C24033 a_66228_12232# VPWR 0.22482f
C24034 a_37084_2727# a_37220_1636# 0.00154f
C24035 a_53572_2824# a_54244_2824# 0.00347f
C24036 a_42460_20452# VPWR 0.01049f
C24037 a_20308_27912# a_21044_27508# 0.00395f
C24038 a_35292_30951# a_35652_31048# 0.08674f
C24039 vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN 0.00271f
C24040 _287_.A1 _462_.D 0.01874f
C24041 _268_.A2 a_53212_27815# 0.00198f
C24042 a_7628_30951# a_7652_29860# 0.0016f
C24043 uio_oe[3] uio_oe[2] 0.0383f
C24044 a_36172_24463# VPWR 0.39641f
C24045 _303_.ZN a_40780_21543# 0.0122f
C24046 a_4068_18884# VPWR 0.2157f
C24047 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.65903f
C24048 a_14236_2727# a_14148_2824# 0.28563f
C24049 a_54432_31128# vgaringosc.ro_inv4.inv_array_notouch_\[3\].I 0.00203f
C24050 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.00154f
C24051 a_53212_15704# VPWR 0.32982f
C24052 _448_.D a_35988_18504# 0.00291f
C24053 a_37360_19325# a_37892_17316# 0.00165f
C24054 _251_.A1 a_56720_26344# 0.01162f
C24055 a_52900_9476# a_53348_9476# 0.01328f
C24056 _397_.A1 _412_.ZN 0.2018f
C24057 _252_.ZN a_61748_26724# 0.0018f
C24058 _324_.C _257_.B 0.01234f
C24059 a_49764_14180# a_49740_13703# 0.00172f
C24060 a_45820_14136# a_45820_13703# 0.05841f
C24061 a_59820_14136# a_60268_14136# 0.01255f
C24062 a_2276_20452# a_2364_20408# 0.28563f
C24063 a_30388_28776# a_32476_28776# 0.01212f
C24064 _460_.Q _359_.ZN 0.40261f
C24065 _355_.C _378_.ZN 0.5567f
C24066 a_57244_27815# VPWR 0.35116f
C24067 _452_.Q a_40452_18180# 0.00179f
C24068 a_48420_12612# a_48060_12568# 0.08707f
C24069 a_14708_24776# a_14708_23588# 0.05841f
C24070 _260_.ZN _448_.Q 0.0657f
C24071 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN a_62060_20408# 0.02545f
C24072 a_45148_1159# a_45508_1256# 0.08717f
C24073 a_60628_12232# a_61076_12232# 0.01328f
C24074 _363_.Z a_35008_27533# 0.55291f
C24075 a_22300_1159# VPWR 0.3289f
C24076 _304_.B _284_.A2 2.06351f
C24077 a_25796_1636# a_25884_1592# 0.28563f
C24078 a_29380_1636# a_29828_1636# 0.01328f
C24079 a_24900_21640# VPWR 0.20614f
C24080 _234_.ZN VPWR 0.43587f
C24081 _424_.B1 a_52512_19715# 0.02316f
C24082 a_51956_26183# a_52304_26399# 0.00277f
C24083 a_51084_10567# a_50996_10664# 0.28563f
C24084 a_49044_28292# VPWR 0.00714f
C24085 _325_.A2 a_40220_19975# 0.00494f
C24086 _424_.B1 a_51428_23340# 0.00118f
C24087 a_33164_24679# a_33524_24776# 0.08674f
C24088 a_63764_23208# VPWR 0.2058f
C24089 a_14796_23544# VPWR 0.30073f
C24090 a_65756_9432# VPWR 0.31505f
C24091 a_2364_2727# VPWR 0.30029f
C24092 a_52428_13703# VPWR 0.31431f
C24093 _459_.CLK a_23912_27967# 0.00137f
C24094 a_67996_6296# VPWR 0.35142f
C24095 a_20956_21543# a_21316_21640# 0.08707f
C24096 a_66004_20072# a_66452_20072# 0.01328f
C24097 a_41476_26344# VPWR 0.21479f
C24098 _441_.A3 a_39985_24372# 0.00631f
C24099 _337_.A3 a_27004_27815# 0.06314f
C24100 _336_.A2 _336_.A1 1.09428f
C24101 a_41664_22020# VPWR 0.01528f
C24102 a_47836_15704# a_48284_15704# 0.01288f
C24103 a_47612_11000# VPWR 0.29679f
C24104 a_31068_28292# VPWR 0.0086f
C24105 a_51780_15748# a_51868_15704# 0.28563f
C24106 _243_.A1 a_58228_27912# 0.00206f
C24107 _439_.ZN _434_.ZN 0.36133f
C24108 _437_.ZN _441_.B 0.11539f
C24109 _304_.ZN a_43156_20452# 0.01212f
C24110 _416_.A1 hold1.Z 0.0029f
C24111 _459_.D a_31348_25156# 0.00261f
C24112 a_3172_26724# VPWR 0.20993f
C24113 _345_.A2 a_23920_27555# 0.00201f
C24114 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN 0.65656f
C24115 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN 0.00793f
C24116 a_58500_26344# VPWR 0.16308f
C24117 a_15156_26344# VPWR 0.20348f
C24118 a_47164_30951# vgaringosc.workerclkbuff_notouch_.I 0.00613f
C24119 a_25212_2727# a_25572_2824# 0.08717f
C24120 _245_.Z a_60013_26344# 0.00353f
C24121 _474_.Q a_49672_19668# 0.00152f
C24122 a_62284_23544# clk 0.00613f
C24123 _460_.Q a_35552_27216# 0.00258f
C24124 a_58500_9476# a_58588_9432# 0.28563f
C24125 a_2812_28248# VPWR 0.30213f
C24126 a_67236_14180# a_67324_14136# 0.28563f
C24127 a_53212_14136# a_53324_13703# 0.02634f
C24128 a_1380_3204# a_1468_3160# 0.28563f
C24129 a_16140_20408# a_16588_20408# 0.0131f
C24130 a_17844_20452# a_18516_20452# 0.00347f
C24131 _409_.ZN uio_in[1] 0.00242f
C24132 _379_.A2 a_19328_28733# 0.00279f
C24133 a_35008_22461# _317_.A2 0.00598f
C24134 _416_.A1 a_45396_25156# 0.0096f
C24135 _465_.D uio_out[6] 0.26849f
C24136 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.01415f
C24137 a_55252_23588# a_54892_23544# 0.08717f
C24138 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN a_59172_23588# 0.00228f
C24139 a_4068_1636# VPWR 0.21569f
C24140 a_65084_30951# vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN 0.00621f
C24141 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN _274_.A2 0.02651f
C24142 a_54916_12612# a_55364_12612# 0.01328f
C24143 a_50996_28292# a_51084_28248# 0.28563f
C24144 _474_.CLK vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.01614f
C24145 _459_.CLK a_24864_29931# 0.01299f
C24146 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN 0.09274f
C24147 a_44700_1159# VPWR 0.29679f
C24148 a_1828_11044# a_1916_11000# 0.28563f
C24149 a_56572_1159# a_56484_1256# 0.28563f
C24150 _284_.A2 VPWR 1.5295f
C24151 a_62532_18884# VPWR 0.20348f
C24152 _281_.ZN _419_.Z 0.00295f
C24153 _362_.ZN _294_.ZN 0.07496f
C24154 _424_.A2 a_52408_19759# 0.01874f
C24155 _373_.ZN a_26970_29480# 0.02521f
C24156 a_61612_10567# a_61972_10664# 0.08707f
C24157 a_47524_10664# a_47972_10664# 0.01328f
C24158 _467_.D a_16588_27815# 0.04913f
C24159 _281_.ZN _399_.A2 0.00143f
C24160 a_16700_1159# a_17148_1159# 0.0131f
C24161 a_57156_1636# a_57020_1159# 0.00168f
C24162 a_17956_2824# a_17956_1636# 0.05841f
C24163 a_18760_29032# _378_.I 0.02388f
C24164 a_55700_23588# a_56148_23588# 0.01328f
C24165 _252_.B a_60013_26344# 0.02793f
C24166 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN 0.08971f
C24167 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I 0.64925f
C24168 _242_.Z a_56516_26344# 0.23952f
C24169 a_15692_21976# VPWR 0.29679f
C24170 _331_.ZN a_40040_17675# 0.00197f
C24171 _452_.Q _435_.ZN 0.11685f
C24172 a_46180_13800# VPWR 0.20348f
C24173 a_46628_2824# a_46716_1159# 0.0027f
C24174 a_31932_21543# a_31844_21640# 0.28563f
C24175 a_19524_21640# a_19972_21640# 0.01328f
C24176 a_24764_2727# VPWR 0.31143f
C24177 a_63068_15271# a_63516_15271# 0.0131f
C24178 a_1916_29816# VPWR 0.297f
C24179 a_55004_21543# a_55140_20452# 0.00154f
C24180 _383_.ZN a_49044_28292# 0.00183f
C24181 a_61412_11044# VPWR 0.20595f
C24182 a_3260_23111# VPWR 0.30487f
C24183 _370_.B _370_.ZN 0.0998f
C24184 _451_.Q _302_.Z 0.01854f
C24185 _402_.ZN a_46156_26031# 0.00108f
C24186 a_25884_27815# a_26556_27815# 0.00544f
C24187 a_66652_15704# a_67100_15704# 0.01255f
C24188 _452_.Q a_43380_20452# 0.00169f
C24189 a_3620_27912# VPWR 0.22347f
C24190 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I 0.10733f
C24191 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN a_62508_23111# 0.00298f
C24192 a_56484_23208# a_56932_23208# 0.01328f
C24193 a_63852_23111# a_63764_23208# 0.28563f
C24194 _274_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I 0.0237f
C24195 a_36636_2727# a_36548_2824# 0.28563f
C24196 _327_.A2 a_41460_22020# 0.00494f
C24197 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I 0.02743f
C24198 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN a_52676_27912# 0.00213f
C24199 a_63740_9432# a_64324_9476# 0.01675f
C24200 a_16948_23588# a_17396_23588# 0.01328f
C24201 a_17508_1256# a_17956_1256# 0.01328f
C24202 a_54356_20072# a_54804_20072# 0.01328f
C24203 _324_.C vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I 0.07002f
C24204 a_64772_6340# a_64860_6296# 0.28563f
C24205 a_66564_6340# a_67012_6340# 0.01328f
C24206 a_65668_7908# a_66116_7908# 0.01328f
C24207 _327_.Z a_38971_18559# 0.00118f
C24208 a_4964_4772# a_4940_4295# 0.00172f
C24209 a_65668_4772# a_65756_4728# 0.28563f
C24210 a_67460_4772# a_67908_4772# 0.01328f
C24211 a_46716_13703# a_47164_13703# 0.0131f
C24212 a_64412_3160# a_64860_3160# 0.0131f
C24213 a_66564_3204# a_66652_3160# 0.28563f
C24214 _452_.CLK a_33948_19975# 0.00866f
C24215 vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I 0.67041f
C24216 a_10092_30951# a_10452_31048# 0.08674f
C24217 a_7964_29383# a_8636_29383# 0.00544f
C24218 _448_.Q _311_.Z 0.00844f
C24219 _452_.CLK a_35628_18407# 0.00854f
C24220 a_62172_17272# a_62284_16839# 0.02634f
C24221 a_10204_1592# VPWR 0.33263f
C24222 a_64884_13800# a_64972_12135# 0.00151f
C24223 _355_.C uio_out[6] 0.716f
C24224 a_61164_20408# a_61276_19975# 0.02634f
C24225 _436_.B _442_.ZN 0.06418f
C24226 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_62420_23208# 0.00593f
C24227 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I 0.03753f
C24228 a_44612_31048# vgaringosc.workerclkbuff_notouch_.I 0.00533f
C24229 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I 0.61661f
C24230 _229_.I vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN 0.15205f
C24231 a_67548_1159# a_67908_1256# 0.08674f
C24232 a_2276_9096# VPWR 0.20634f
C24233 a_31708_19975# VPWR 0.31436f
C24234 a_67100_1159# VPWR 0.3289f
C24235 a_4068_5960# VPWR 0.22146f
C24236 _452_.CLK a_31732_22020# 0.00239f
C24237 a_49764_11044# a_50212_11044# 0.01328f
C24238 a_33052_18407# VPWR 0.29736f
C24239 a_46180_11044# a_46268_11000# 0.28563f
C24240 a_7652_1636# a_7516_1159# 0.00168f
C24241 a_3708_1592# a_3708_1159# 0.05841f
C24242 a_35516_1592# a_35964_1592# 0.01288f
C24243 a_39460_1636# a_39548_1592# 0.28563f
C24244 a_61748_23588# a_61836_23544# 0.28563f
C24245 a_32964_16936# a_33412_16936# 0.01328f
C24246 _399_.ZN a_48529_22460# 0.00171f
C24247 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_55956_25940# 0.05116f
C24248 a_56964_26724# vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I 0.00394f
C24249 _319_.A2 _325_.A2 0.00447f
C24250 _330_.A1 _470_.D 0.98524f
C24251 a_16252_30951# uio_oe[0] 0.03219f
C24252 _257_.B _252_.ZN 0.01196f
C24253 a_39256_28292# VPWR 0.60322f
C24254 a_35008_27533# a_35660_27508# 0.00587f
C24255 _294_.A2 a_31484_30951# 0.00616f
C24256 _459_.CLK a_32132_27912# 0.0079f
C24257 a_29356_21976# VPWR 0.31547f
C24258 a_34980_22895# _316_.A3 0.00125f
C24259 a_23084_28248# VPWR 0.30527f
C24260 _256_.A2 _247_.ZN 0.00864f
C24261 _465_.D a_20250_31048# 0.02753f
C24262 _325_.A2 _325_.B 0.42737f
C24263 _304_.B a_52452_24072# 0.06196f
C24264 a_44252_30951# a_44700_30951# 0.0131f
C24265 a_47164_2727# VPWR 0.31143f
C24266 _276_.A2 _268_.A1 0.01246f
C24267 a_68020_13800# VPWR 0.21406f
C24268 a_37360_19325# a_37067_19001# 0.49319f
C24269 a_58063_30644# _272_.B1 0.00592f
C24270 a_14796_26247# a_15156_26344# 0.08717f
C24271 a_34708_29860# VPWR 0.01593f
C24272 a_15580_29816# VPWR 0.29679f
C24273 _421_.B a_46476_20937# 0.00855f
C24274 a_65332_16936# a_65308_15704# 0.0016f
C24275 a_48060_10567# VPWR 0.29679f
C24276 a_33500_15271# a_33860_15368# 0.08717f
C24277 _281_.ZN _424_.A1 0.00755f
C24278 a_932_23208# VPWR 0.22176f
C24279 a_49764_26724# a_49952_26724# 0.0101f
C24280 _284_.B _260_.A2 0.00514f
C24281 a_46252_19759# a_46596_20127# 0.00275f
C24282 _359_.B _358_.A3 0.1173f
C24283 a_1828_28292# a_2276_28292# 0.01328f
C24284 a_47612_2727# a_47972_2824# 0.08717f
C24285 a_63876_17316# a_63964_17272# 0.28563f
C24286 a_54892_19975# a_55252_20072# 0.08663f
C24287 a_54192_22851# a_54604_23263# 0.00275f
C24288 a_56124_23111# a_56036_23208# 0.28563f
C24289 a_2276_16936# a_2276_15748# 0.05841f
C24290 a_67100_9432# a_67100_8999# 0.05841f
C24291 a_15604_25156# a_16052_25156# 0.01328f
C24292 a_1020_7431# a_932_7528# 0.28563f
C24293 a_41056_30669# a_41264_30669# 0.00372f
C24294 a_35204_31048# VPWR 0.23867f
C24295 _287_.A2 _294_.ZN 0.04066f
C24296 a_4156_13703# a_4068_13800# 0.28563f
C24297 _369_.ZN _337_.ZN 0.19519f
C24298 a_66787_30600# a_67237_31198# 0.00209f
C24299 a_27116_20408# a_27564_20408# 0.0131f
C24300 a_29268_20452# a_28908_20408# 0.08717f
C24301 a_65220_18504# a_65220_17316# 0.05841f
C24302 a_46356_24072# a_46580_23588# 0.01342f
C24303 a_54804_24776# a_54804_23588# 0.05841f
C24304 a_30812_16839# a_30724_16936# 0.28563f
C24305 _419_.Z a_50660_20452# 0.0106f
C24306 _441_.ZN _452_.Q 0.05162f
C24307 a_17786_29480# uio_out[7] 0.00151f
C24308 a_61500_12568# a_61948_12568# 0.01288f
C24309 a_23868_1592# VPWR 0.32517f
C24310 a_37756_1592# a_37892_1256# 0.00168f
C24311 a_65444_12612# a_65084_12568# 0.08707f
C24312 _304_.B a_40692_27912# 0.00141f
C24313 _381_.Z _397_.A4 0.02663f
C24314 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN 0.01244f
C24315 a_42820_1636# a_42460_1592# 0.08707f
C24316 a_51892_12232# a_51980_10567# 0.00151f
C24317 _362_.ZN a_33140_29860# 0.00494f
C24318 a_39100_1159# a_39548_1159# 0.0131f
C24319 a_12356_29860# uio_oe[3] 0.00519f
C24320 _402_.A1 _324_.B 0.02693f
C24321 a_5052_20408# VPWR 0.33516f
C24322 a_52452_24072# VPWR 0.30323f
C24323 _452_.CLK _312_.ZN 0.00111f
C24324 a_4852_27912# a_4940_26247# 0.00151f
C24325 a_63540_16936# a_63988_16936# 0.01328f
C24326 a_49404_12568# VPWR 0.32055f
C24327 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN rst_n 0.00617f
C24328 _284_.ZN a_39300_29480# 0.00911f
C24329 a_21424_25987# a_22059_26399# 0.02112f
C24330 a_20496_26344# a_22352_25987# 0.02307f
C24331 a_43044_15368# a_43492_15368# 0.01328f
C24332 _355_.C a_20250_31048# 0.00869f
C24333 a_6620_29383# a_6532_29480# 0.28563f
C24334 _452_.CLK a_38971_18559# 0.024f
C24335 a_55676_27815# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I 0.00505f
C24336 a_2276_10664# VPWR 0.20634f
C24337 a_44924_15271# a_44836_15368# 0.28563f
C24338 _416_.A2 a_47612_18407# 0.00109f
C24339 a_31844_23208# VPWR 0.20622f
C24340 _435_.ZN a_40357_24776# 0.04128f
C24341 _324_.C a_51332_24072# 0.39279f
C24342 _304_.B a_41160_29083# 0.076f
C24343 _459_.CLK a_18264_29480# 0.00343f
C24344 _272_.B1 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I 0.00343f
C24345 a_20672_30301# _375_.Z 0.00608f
C24346 a_46492_15271# a_46940_15271# 0.0131f
C24347 a_16500_28292# a_16140_28248# 0.08663f
C24348 _237_.A1 _272_.A2 0.01907f
C24349 _336_.A1 a_29136_25641# 0.00157f
C24350 _447_.Q a_43750_23544# 0.06493f
C24351 a_59036_2727# a_58948_2824# 0.28563f
C24352 a_17844_22020# a_18292_22020# 0.01328f
C24353 _459_.Q a_31820_23544# 0.00111f
C24354 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN 0.08406f
C24355 a_2812_16839# a_3260_16839# 0.0131f
C24356 _300_.ZN a_39324_19975# 0.00147f
C24357 _416_.A1 clkbuf_1_0__f_clk.I 0.11988f
C24358 a_67460_15748# VPWR 0.20622f
C24359 _245_.I1 a_62560_25112# 0.02473f
C24360 _358_.A3 a_32144_26724# 0.00135f
C24361 a_36996_21640# a_37444_21640# 0.01328f
C24362 a_43356_30951# a_43268_31048# 0.28563f
C24363 a_35988_16936# a_36100_15748# 0.02666f
C24364 a_46316_29977# VPWR 0.00246f
C24365 a_24452_23208# a_24540_21543# 0.00151f
C24366 _332_.Z a_41048_17341# 0.00372f
C24367 a_17732_31048# VPWR 0.20878f
C24368 a_39908_1256# a_40356_1256# 0.01328f
C24369 a_27924_23588# a_27564_23544# 0.08674f
C24370 a_24428_23544# a_24876_23544# 0.0131f
C24371 a_1468_7864# VPWR 0.29679f
C24372 a_11684_1256# VPWR 0.24201f
C24373 _448_.Q a_39780_22805# 0.00201f
C24374 _384_.ZN a_48859_29076# 0.01006f
C24375 a_23060_26724# VPWR 0.01385f
C24376 a_3260_4728# VPWR 0.30487f
C24377 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I 0.0181f
C24378 a_58063_30644# VPWR 0.8339f
C24379 a_18940_2727# a_19388_2727# 0.0131f
C24380 a_54668_13703# a_55028_13800# 0.08707f
C24381 a_2364_29383# VPWR 0.30029f
C24382 a_932_13800# a_1380_13800# 0.01328f
C24383 _370_.B a_31068_28292# 0.00303f
C24384 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN 0.73688f
C24385 a_2364_17272# a_2364_16839# 0.05841f
C24386 a_55700_25156# a_55340_25112# 0.08663f
C24387 _327_.Z a_40636_18180# 0.00207f
C24388 a_62564_29032# a_61940_29076# 0.00587f
C24389 a_59796_29480# a_59572_29076# 0.01751f
C24390 a_41452_16839# a_41812_16936# 0.08663f
C24391 a_48420_10664# a_48420_9476# 0.05841f
C24392 _284_.A2 a_44744_26355# 0.00123f
C24393 a_57132_10567# a_57156_9476# 0.0016f
C24394 a_2276_16936# VPWR 0.20634f
C24395 a_37668_1636# VPWR 0.2085f
C24396 a_19276_23544# a_19164_23111# 0.02634f
C24397 _460_.Q a_35108_28776# 0.00106f
C24398 a_5860_1636# a_5500_1592# 0.08707f
C24399 a_40692_27912# VPWR 0.1242f
C24400 a_4068_29860# a_4516_29860# 0.01328f
C24401 a_45800_30345# _393_.ZN 0.00828f
C24402 a_1468_17272# a_1916_17272# 0.0131f
C24403 a_4068_17316# a_3708_17272# 0.08717f
C24404 _296_.ZN VPWR 0.95874f
C24405 _229_.I a_60852_28292# 0.01594f
C24406 a_59844_11044# a_59932_11000# 0.28563f
C24407 a_55900_11000# a_56348_11000# 0.01288f
C24408 a_49316_1636# a_49764_1636# 0.01328f
C24409 a_55788_25112# VPWR 0.3101f
C24410 vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN 0.62756f
C24411 a_3172_20072# a_3172_18884# 0.05841f
C24412 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN a_54444_18407# 0.00105f
C24413 a_47076_18504# a_47052_16839# 0.00131f
C24414 a_62172_18407# VPWR 0.29679f
C24415 a_1020_25112# VPWR 0.30073f
C24416 a_63876_18884# a_63516_18840# 0.08717f
C24417 a_17484_27815# a_17932_27815# 0.0131f
C24418 a_3260_27815# a_3620_27912# 0.08717f
C24419 a_25100_20408# VPWR 0.31143f
C24420 a_4964_15748# a_5052_15704# 0.28563f
C24421 a_63204_12612# VPWR 0.20595f
C24422 a_19972_2824# a_20420_2824# 0.01328f
C24423 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I a_66004_20072# 0.00184f
C24424 a_58656_27912# VPWR 0.00723f
C24425 a_61300_15748# VPWR 0.20924f
C24426 _311_.A2 a_36212_23588# 0.0107f
C24427 a_64860_8999# a_64772_9096# 0.28563f
C24428 a_55340_24679# clk 0.01858f
C24429 a_53460_24776# a_53908_24776# 0.01328f
C24430 a_63764_10664# VPWR 0.20674f
C24431 a_65756_7431# a_65668_7528# 0.28563f
C24432 _371_.A1 a_33764_27208# 0.00889f
C24433 a_66652_5863# a_66564_5960# 0.28563f
C24434 a_55900_15271# a_56260_15368# 0.08717f
C24435 _287_.A2 a_30778_31048# 0.02497f
C24436 a_67548_4295# a_67460_4392# 0.28563f
C24437 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I 0.72199f
C24438 a_41160_29083# VPWR 1.0095f
C24439 a_37220_15368# VPWR 0.20348f
C24440 _457_.D a_25236_23588# 0.00167f
C24441 _257_.B a_59796_29480# 0.00238f
C24442 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_56236_24679# 0.03116f
C24443 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I VPWR 0.79501f
C24444 a_40668_15271# VPWR 0.32938f
C24445 hold2.Z a_41476_24776# 0.00141f
C24446 a_1468_14136# a_1916_14136# 0.0131f
C24447 a_4068_14180# a_3708_14136# 0.08717f
C24448 a_64860_17272# VPWR 0.31855f
C24449 a_39124_16936# a_39100_15704# 0.0016f
C24450 a_42932_16936# a_43044_15748# 0.02666f
C24451 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN VPWR 0.72566f
C24452 _324_.C a_42587_25940# 0.0093f
C24453 a_34084_1256# VPWR 0.20902f
C24454 _448_.Q a_39796_22504# 0.15337f
C24455 a_65868_13703# a_65780_13800# 0.28563f
C24456 _455_.D a_20928_26399# 0.00245f
C24457 a_17820_30951# VPWR 0.31143f
C24458 a_57244_27815# a_57156_27912# 0.28563f
C24459 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I a_59732_14180# 0.00504f
C24460 _416_.A1 a_46580_28292# 0.00253f
C24461 a_61860_30736# ui_in[1] 0.03592f
C24462 a_52652_16839# a_52564_16936# 0.28563f
C24463 a_67796_18504# VPWR 0.2115f
C24464 a_64300_10567# a_64324_9476# 0.0016f
C24465 a_11324_1159# a_11684_1256# 0.08717f
C24466 a_49204_16936# VPWR 0.21075f
C24467 _229_.I _238_.I 0.08647f
C24468 a_43804_1592# VPWR 0.29679f
C24469 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN 0.00209f
C24470 a_55564_12135# a_56012_12135# 0.01288f
C24471 a_1916_12135# a_2276_12232# 0.08717f
C24472 a_8772_1636# a_8860_1592# 0.28563f
C24473 a_12356_1636# a_12804_1636# 0.01328f
C24474 a_4740_29480# a_5188_29480# 0.01328f
C24475 _411_.A2 a_50792_26344# 0.1336f
C24476 a_61636_20072# a_61724_18407# 0.0027f
C24477 _424_.A2 a_45564_21236# 0.00939f
C24478 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I VPWR 0.7662f
C24479 a_33860_17316# a_33500_17272# 0.08707f
C24480 a_39536_26795# a_40092_27209# 0.8399f
C24481 a_63204_11044# a_63292_11000# 0.28563f
C24482 _330_.A1 a_39324_26247# 0.00359f
C24483 _442_.ZN a_40464_27165# 0.00761f
C24484 a_14148_2824# VPWR 0.20348f
C24485 _371_.A1 uo_out[6] 0.16778f
C24486 a_37084_26680# VPWR 0.29679f
C24487 _459_.CLK a_19524_26344# 0.00809f
C24488 a_17932_24679# a_18716_24679# 0.00443f
C24489 a_61276_1159# a_61948_1159# 0.00544f
C24490 a_1020_19975# a_1468_19975# 0.0131f
C24491 _437_.A1 a_38523_27967# 0.06037f
C24492 _455_.Q a_23420_26247# 0.01486f
C24493 a_67684_15368# VPWR 0.20893f
C24494 a_2364_18407# a_2812_18407# 0.0131f
C24495 a_52639_30644# _267_.A2 0.00204f
C24496 a_23084_25112# VPWR 0.3262f
C24497 a_58924_18840# vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I 0.01358f
C24498 _334_.A1 a_32240_31048# 0.10749f
C24499 a_34756_15748# a_34844_15704# 0.28563f
C24500 a_30812_15704# a_31260_15704# 0.01288f
C24501 a_50188_12135# VPWR 0.32969f
C24502 a_52116_18504# a_52228_17316# 0.02666f
C24503 a_48420_18504# a_48284_17272# 0.00154f
C24504 a_22748_2727# a_22884_1636# 0.00154f
C24505 a_44795_29535# a_45080_29535# 0.00277f
C24506 _427_.A2 a_53704_23219# 0.0089f
C24507 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN 0.00143f
C24508 a_52639_30644# a_53212_29816# 0.01891f
C24509 a_3260_24679# VPWR 0.30487f
C24510 a_27228_26247# a_27676_26247# 0.01222f
C24511 _450_.D VPWR 0.78817f
C24512 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN ui_in[7] 0.00758f
C24513 _474_.CLK _276_.A2 0.72683f
C24514 _436_.B _441_.ZN 0.00243f
C24515 a_43156_20452# _328_.A2 0.00127f
C24516 a_32964_15748# VPWR 0.20348f
C24517 _355_.C a_27924_24776# 0.00688f
C24518 _362_.ZN _362_.B 0.01229f
C24519 a_25796_27912# VPWR 0.1658f
C24520 _324_.C _303_.ZN 0.00256f
C24521 a_46268_18407# a_46716_18407# 0.0131f
C24522 a_27924_22020# a_28012_21976# 0.28563f
C24523 a_23980_21976# a_24428_21976# 0.01288f
C24524 _304_.B _419_.A4 0.00433f
C24525 a_48420_14180# a_48060_14136# 0.08707f
C24526 a_49740_16839# a_50412_16839# 0.00544f
C24527 _452_.CLK a_37084_17272# 0.00599f
C24528 _350_.A2 a_28928_29123# 0.00583f
C24529 a_44364_16839# VPWR 0.29679f
C24530 a_52360_26355# a_52744_26031# 1.16391f
C24531 _275_.ZN _409_.ZN 0.00314f
C24532 a_21204_31048# uio_out[5] 0.03327f
C24533 a_62308_1256# a_62756_1256# 0.01328f
C24534 _325_.A1 a_41776_20072# 0.01051f
C24535 a_56484_1256# VPWR 0.20488f
C24536 _346_.ZN a_21600_26725# 0.01027f
C24537 a_41340_2727# a_41788_2727# 0.0131f
C24538 a_54020_21640# a_53884_20408# 0.00154f
C24539 a_62420_13800# a_62868_13800# 0.01328f
C24540 a_44364_17272# a_44364_16839# 0.05841f
C24541 a_34844_17272# VPWR 0.35856f
C24542 a_34716_20937# _319_.A2 0.00193f
C24543 a_57604_1636# VPWR 0.21525f
C24544 a_22748_1159# a_22660_1256# 0.28563f
C24545 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I 0.00753f
C24546 a_52876_12135# a_52788_12232# 0.28563f
C24547 a_61940_29076# _250_.B 0.01434f
C24548 _362_.ZN a_32628_26725# 0.09042f
C24549 a_14148_29860# a_14236_29816# 0.28563f
C24550 a_10204_29816# a_10652_29816# 0.01288f
C24551 a_44276_17316# a_44724_17316# 0.01328f
C24552 a_2812_10567# a_3260_10567# 0.0131f
C24553 a_29232_29931# VPWR 1.10884f
C24554 a_60380_11000# a_60268_10567# 0.02634f
C24555 a_54356_25156# clk 0.00147f
C24556 a_36548_2824# VPWR 0.20815f
C24557 _237_.A1 _228_.ZN 0.17599f
C24558 a_59396_1636# a_59484_1592# 0.28563f
C24559 a_35876_1636# a_35740_1159# 0.00168f
C24560 _324_.C _397_.A4 1.94007f
C24561 _274_.A3 a_52756_29076# 0.03372f
C24562 a_28796_23111# a_29244_23111# 0.01288f
C24563 _459_.CLK a_16948_27912# 0.02618f
C24564 a_16588_23111# a_16948_23208# 0.08717f
C24565 a_20508_24679# a_20868_24776# 0.08707f
C24566 _455_.Q _346_.ZN 0.91659f
C24567 a_3708_9432# VPWR 0.33374f
C24568 a_1916_21543# a_2364_21543# 0.0131f
C24569 a_53124_2824# a_52988_1592# 0.00154f
C24570 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_55252_25156# 0.00142f
C24571 a_55956_25940# a_55700_25156# 0.00121f
C24572 _316_.A3 a_35268_21640# 0.02114f
C24573 a_49404_14136# VPWR 0.32055f
C24574 _400_.ZN a_45128_26031# 0.00698f
C24575 _279_.Z clk 0.03699f
C24576 _251_.A1 a_63180_26680# 0.00799f
C24577 a_33052_18407# a_32964_18504# 0.28563f
C24578 _335_.ZN VPWR 2.70082f
C24579 a_37556_23588# _439_.ZN 0.0029f
C24580 _304_.A1 a_36300_23544# 0.0152f
C24581 _350_.A2 _336_.Z 0.00257f
C24582 a_17596_29816# uio_out[7] 0.00448f
C24583 a_35728_29480# uo_out[2] 0.00171f
C24584 a_4068_12232# VPWR 0.22146f
C24585 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62396_27815# 0.04095f
C24586 a_50972_15704# a_51108_15368# 0.00168f
C24587 a_42148_2824# a_42820_2824# 0.00347f
C24588 _474_.CLK _395_.A1 0.00416f
C24589 _363_.Z _365_.ZN 0.83704f
C24590 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I VPWR 1.25873f
C24591 a_16948_24776# VPWR 0.20348f
C24592 _340_.A2 a_24864_29931# 0.15543f
C24593 a_41188_18840# a_41804_19376# 0.00478f
C24594 a_2812_2727# a_2724_2824# 0.28563f
C24595 a_39100_15704# VPWR 0.3289f
C24596 a_4156_19975# a_4852_20072# 0.01227f
C24597 a_5300_20072# a_5388_18407# 0.0027f
C24598 _459_.CLK a_21600_26725# 0.04722f
C24599 a_45372_9432# a_45820_9432# 0.0131f
C24600 a_47524_9476# a_47164_9432# 0.08717f
C24601 _451_.Q a_39264_18147# 0.1934f
C24602 _324_.C a_43788_29167# 0.00665f
C24603 _350_.A1 a_29788_30345# 0.02988f
C24604 a_54916_14180# a_55364_14180# 0.01328f
C24605 _419_.A4 VPWR 1.23624f
C24606 _327_.A2 a_41776_20072# 0.00123f
C24607 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_56036_28292# 0.00315f
C24608 _444_.D a_37108_23588# 0.00308f
C24609 _265_.ZN a_42596_27912# 0.01784f
C24610 _304_.B a_56124_27815# 0.00116f
C24611 _435_.A3 a_39587_24372# 0.00116f
C24612 a_3620_12612# a_3708_12568# 0.28563f
C24613 a_53548_18407# a_53572_17316# 0.0016f
C24614 _281_.ZN _399_.ZN 0.105f
C24615 a_36212_23588# a_36660_23588# 0.01328f
C24616 a_51420_17272# a_51308_16839# 0.02634f
C24617 _336_.A2 a_27676_26247# 0.00972f
C24618 a_29156_23208# a_29268_22020# 0.02666f
C24619 a_46940_17272# VPWR 0.31389f
C24620 a_25348_23208# a_25324_21976# 0.0016f
C24621 _331_.ZN _332_.Z 0.5231f
C24622 a_33724_1159# a_34084_1256# 0.08717f
C24623 a_66876_1592# VPWR 0.3289f
C24624 _378_.I a_21103_29076# 0.00367f
C24625 a_63404_12135# a_63764_12232# 0.08707f
C24626 _282_.ZN a_46794_25156# 0.02503f
C24627 _252_.B a_59172_26724# 0.00702f
C24628 a_18492_1592# a_18940_1592# 0.01288f
C24629 a_22436_1636# a_22524_1592# 0.28563f
C24630 a_49652_12232# a_50100_12232# 0.01328f
C24631 _287_.A1 a_35818_29860# 0.00303f
C24632 a_27452_21543# VPWR 0.32285f
C24633 a_18044_29816# _459_.CLK 0.07874f
C24634 _304_.B a_40038_28720# 0.00315f
C24635 _352_.A2 a_31116_26020# 0.00187f
C24636 _459_.CLK _455_.Q 0.4914f
C24637 a_39760_23588# VPWR 0.01382f
C24638 a_58948_2824# VPWR 0.20348f
C24639 a_64100_1636# a_64188_1592# 0.28563f
C24640 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I 0.00107f
C24641 a_3620_2824# a_3620_1636# 0.05841f
C24642 _428_.Z _427_.A2 0.08852f
C24643 a_27900_23111# a_27812_23208# 0.28563f
C24644 a_22660_24776# a_23108_24776# 0.01328f
C24645 _452_.CLK a_45920_20523# 0.01004f
C24646 _452_.Q a_41488_24072# 0.51975f
C24647 a_54332_9432# VPWR 0.31143f
C24648 a_64996_14180# VPWR 0.20816f
C24649 _304_.B a_41028_26344# 0.00796f
C24650 _324_.C a_44864_27165# 0.00203f
C24651 _287_.A2 _362_.B 0.00591f
C24652 _350_.A2 uio_out[0] 0.00188f
C24653 _281_.A1 a_54020_21640# 0.00183f
C24654 _402_.A1 uo_out[1] 0.00135f
C24655 _416_.A1 a_45732_18884# 0.0015f
C24656 a_65780_12232# VPWR 0.22327f
C24657 a_44476_15704# a_44924_15704# 0.01288f
C24658 _325_.A2 a_40416_18885# 0.00411f
C24659 a_35292_30951# a_35204_31048# 0.28563f
C24660 a_63516_18840# a_63516_18407# 0.05841f
C24661 a_67908_18884# a_67884_18407# 0.00172f
C24662 _303_.ZN a_40332_21543# 0.00838f
C24663 a_36544_24419# VPWR 0.18864f
C24664 a_3620_18884# VPWR 0.22347f
C24665 a_13788_2727# a_14148_2824# 0.08717f
C24666 a_52764_15704# VPWR 0.32975f
C24667 a_66092_19975# a_66540_19975# 0.01255f
C24668 _251_.A1 a_56368_26344# 0.00208f
C24669 _252_.ZN a_60828_26680# 0.00571f
C24670 _324_.C a_52756_29076# 0.0057f
C24671 a_48732_17272# a_48644_15748# 0.00151f
C24672 a_2276_20452# a_1916_20408# 0.08717f
C24673 a_4068_20452# a_4516_20452# 0.01328f
C24674 _384_.ZN clkload0.Z 0.083f
C24675 _355_.C a_17472_28363# 0.06392f
C24676 _294_.A2 a_33476_27912# 0.00164f
C24677 a_56124_27815# VPWR 0.30114f
C24678 _336_.Z a_29804_23544# 0.01171f
C24679 _229_.I VPWR 2.03774f
C24680 a_47972_12612# a_48060_12568# 0.28563f
C24681 a_63740_2727# a_64188_2727# 0.0131f
C24682 a_51556_12612# a_52004_12612# 0.01328f
C24683 a_21852_1159# VPWR 0.3289f
C24684 a_66116_9096# a_66116_7908# 0.05841f
C24685 a_45148_1159# a_45060_1256# 0.28563f
C24686 a_32516_20072# a_32964_20072# 0.01328f
C24687 a_67012_7528# a_67012_6340# 0.05841f
C24688 a_64188_12568# a_64100_11044# 0.00151f
C24689 _304_.B a_51048_26680# 0.00571f
C24690 a_25796_1636# a_25436_1592# 0.08707f
C24691 a_24452_21640# VPWR 0.20614f
C24692 a_37532_26247# a_37980_26247# 0.012f
C24693 a_40038_28720# VPWR 0.79818f
C24694 _424_.B1 a_52024_20083# 0.03823f
C24695 a_52316_17272# a_52764_17272# 0.01288f
C24696 a_64300_10567# a_64972_10567# 0.00544f
C24697 a_50636_10567# a_50996_10664# 0.08707f
C24698 a_5276_1159# a_5724_1159# 0.0131f
C24699 _402_.A1 a_49172_27508# 0.00146f
C24700 _325_.A2 a_39772_19975# 0.00839f
C24701 a_48820_28292# VPWR 0.01425f
C24702 a_26468_23208# a_26916_23208# 0.01328f
C24703 _424_.B1 a_50732_23233# 0.00293f
C24704 a_63316_23208# VPWR 0.20348f
C24705 a_33164_24679# a_33076_24776# 0.28563f
C24706 _474_.CLK _397_.A1 0.27168f
C24707 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN 0.00631f
C24708 a_21876_23588# VPWR 0.21241f
C24709 a_67548_6296# VPWR 0.29679f
C24710 a_19524_26344# a_19612_24679# 0.00151f
C24711 a_20956_21543# a_20868_21640# 0.28563f
C24712 a_65308_9432# VPWR 0.30378f
C24713 a_32828_21543# a_33276_21543# 0.01288f
C24714 _379_.Z a_18028_28777# 0.00467f
C24715 a_35204_2824# a_35292_1159# 0.0027f
C24716 a_1916_2727# VPWR 0.297f
C24717 a_51980_13703# VPWR 0.31431f
C24718 _441_.A3 a_39781_24372# 0.00263f
C24719 _337_.A3 a_26556_27815# 0.01707f
C24720 _455_.Q _371_.A3 0.01381f
C24721 a_41028_26344# VPWR 0.21024f
C24722 _365_.ZN uo_out[3] 0.00678f
C24723 _359_.B uo_out[1] 0.05549f
C24724 _279_.Z _416_.A3 0.00102f
C24725 _301_.Z a_38340_21327# 0.21679f
C24726 a_47164_11000# VPWR 0.29679f
C24727 a_41460_22020# VPWR 0.00709f
C24728 a_51780_15748# a_51420_15704# 0.08707f
C24729 a_14684_29816# a_14684_29383# 0.05841f
C24730 a_30596_28292# VPWR 0.02076f
C24731 _476_.Q _474_.D 0.16493f
C24732 _395_.A1 _398_.C 0.13515f
C24733 _437_.ZN a_38759_24072# 0.00513f
C24734 a_64548_2824# a_64996_2824# 0.01328f
C24735 _459_.D a_31124_25156# 0.00883f
C24736 a_2724_26724# VPWR 0.20782f
C24737 _304_.ZN a_42728_20452# 0.00117f
C24738 _223_.I a_31396_26724# 0.03595f
C24739 a_14908_30951# a_15044_29860# 0.00154f
C24740 _250_.ZN _250_.A2 0.25725f
C24741 _345_.A2 a_23627_27967# 0.00691f
C24742 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62756_27912# 0.00728f
C24743 a_32180_20452# a_32156_19975# 0.00172f
C24744 a_62084_15748# a_62532_15748# 0.01328f
C24745 _459_.CLK _330_.A1 0.00104f
C24746 a_14708_26344# VPWR 0.22176f
C24747 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I a_58252_18407# 0.00769f
C24748 a_25212_2727# a_25124_2824# 0.28563f
C24749 a_46716_30951# vgaringosc.workerclkbuff_notouch_.I 0.00613f
C24750 _245_.Z a_59397_26344# 0.00217f
C24751 a_61836_23544# clk 0.00613f
C24752 _365_.ZN a_35660_27508# 0.38386f
C24753 _416_.A1 a_44476_27815# 0.04368f
C24754 a_6084_1256# a_6532_1256# 0.01328f
C24755 _442_.ZN _261_.ZN 0.00819f
C24756 a_2364_28248# VPWR 0.30029f
C24757 a_1380_23588# a_1828_23588# 0.01328f
C24758 a_58500_9476# a_58140_9432# 0.08717f
C24759 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN 0.79547f
C24760 a_2276_4772# a_2724_4772# 0.01328f
C24761 _436_.B a_42148_27912# 0.0019f
C24762 _393_.ZN a_45088_29123# 0.00458f
C24763 a_7092_31048# a_7540_31048# 0.01328f
C24764 a_1380_6340# a_1828_6340# 0.01328f
C24765 a_1380_3204# a_1020_3160# 0.08717f
C24766 a_3172_3204# a_3620_3204# 0.01328f
C24767 a_67236_14180# a_66876_14136# 0.08707f
C24768 a_63292_14136# a_63740_14136# 0.01288f
C24769 a_17844_20452# a_17932_20408# 0.28563f
C24770 a_34715_22137# a_34960_22505# 0.00232f
C24771 a_35008_22461# a_36148_21976# 0.00995f
C24772 a_54804_23588# a_54892_23544# 0.28563f
C24773 _416_.A1 a_44948_25156# 0.0065f
C24774 _258_.I _258_.ZN 0.60439f
C24775 _350_.A1 _288_.ZN 0.09914f
C24776 a_63616_31128# vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN 0.00346f
C24777 a_3620_1636# VPWR 0.22347f
C24778 _343_.A2 VPWR 1.43764f
C24779 a_53684_13800# a_53772_12135# 0.00151f
C24780 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN 0.00116f
C24781 a_56124_1159# a_56484_1256# 0.08717f
C24782 a_44252_1159# VPWR 0.29679f
C24783 a_5948_29816# a_6084_29480# 0.00168f
C24784 a_3620_11044# a_4068_11044# 0.01328f
C24785 a_1828_11044# a_1468_11000# 0.08717f
C24786 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I VPWR 0.80678f
C24787 a_64076_16839# a_64524_16839# 0.0131f
C24788 a_51048_26680# VPWR 0.31071f
C24789 a_32292_1636# a_32740_1636# 0.01328f
C24790 a_62084_18884# VPWR 0.22588f
C24791 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN 0.00239f
C24792 _435_.ZN _433_.ZN 0.08253f
C24793 a_42236_27815# a_42684_27815# 0.01255f
C24794 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_59732_13800# 0.00123f
C24795 _424_.A2 a_52512_19715# 0.0208f
C24796 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I 0.0042f
C24797 _467_.D a_16140_27815# 0.01312f
C24798 a_62196_23588# a_62060_23111# 0.00168f
C24799 a_61612_10567# a_61524_10664# 0.28563f
C24800 a_4068_18504# a_4068_17316# 0.05841f
C24801 VPWR rst_n 0.64989f
C24802 a_54916_21640# a_55364_21640# 0.01328f
C24803 a_15244_21976# VPWR 0.29679f
C24804 _252_.B a_59397_26344# 0.10877f
C24805 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN a_65668_23208# 0.0063f
C24806 _304_.B _381_.A2 0.17867f
C24807 a_29716_23588# VPWR 0.1307f
C24808 a_31484_21543# a_31844_21640# 0.08707f
C24809 _475_.D a_47531_21258# 0.00602f
C24810 a_24316_2727# VPWR 0.31143f
C24811 a_4604_18840# a_5052_18840# 0.01222f
C24812 a_45732_13800# VPWR 0.20348f
C24813 a_60276_29032# a_59572_29076# 0.00142f
C24814 a_1468_29816# VPWR 0.29679f
C24815 a_60964_11044# VPWR 0.2267f
C24816 _383_.ZN a_48820_28292# 0.0063f
C24817 _324_.B a_42982_21730# 0.00204f
C24818 _438_.A2 _435_.A3 0.20486f
C24819 a_20084_22020# a_20060_21543# 0.00172f
C24820 a_16140_21976# a_16140_21543# 0.05841f
C24821 a_50972_2727# a_51108_1636# 0.00154f
C24822 a_2812_23111# VPWR 0.30213f
C24823 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN VPWR 0.96003f
C24824 _452_.Q a_43156_20452# 0.00401f
C24825 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN a_62560_25112# 0.07943f
C24826 a_3172_27912# VPWR 0.20993f
C24827 _424_.A2 _282_.ZN 0.09109f
C24828 _393_.A3 _395_.A1 0.33145f
C24829 a_36188_2727# a_36548_2824# 0.08717f
C24830 a_63404_23111# a_63764_23208# 0.08717f
C24831 _460_.Q _371_.A1 1.30955f
C24832 _478_.D a_54420_21976# 0.00807f
C24833 _319_.A3 a_36008_20569# 0.00142f
C24834 _370_.B _335_.ZN 0.01111f
C24835 _324_.C a_64324_29860# 0.00135f
C24836 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN a_52228_27912# 0.0026f
C24837 a_1468_6296# a_1468_5863# 0.05841f
C24838 a_64772_6340# a_64412_6296# 0.08717f
C24839 _397_.A2 _281_.ZN 0.66088f
C24840 a_2364_4728# a_2364_4295# 0.05841f
C24841 a_65668_4772# a_65308_4728# 0.08717f
C24842 a_66564_3204# a_66204_3160# 0.08717f
C24843 a_3260_3160# a_3260_2727# 0.05841f
C24844 a_23220_20452# a_23668_20452# 0.01328f
C24845 a_10092_30951# a_10004_31048# 0.28563f
C24846 _244_.Z vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I 0.08124f
C24847 a_66116_17316# a_66092_16839# 0.00172f
C24848 _379_.A2 uio_out[7] 0.93732f
C24849 _452_.CLK a_35180_18407# 0.0147f
C24850 a_9756_1592# VPWR 0.32966f
C24851 a_57692_12568# a_58140_12568# 0.01288f
C24852 _223_.I VPWR 1.42952f
C24853 a_39884_27815# _442_.ZN 0.00103f
C24854 _436_.B a_39536_26795# 0.0883f
C24855 a_66988_19975# a_67012_18884# 0.0016f
C24856 a_44164_31048# vgaringosc.workerclkbuff_notouch_.I 0.00557f
C24857 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN a_58164_18504# 0.00315f
C24858 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_61972_23208# 0.03719f
C24859 a_46180_11044# a_45820_11000# 0.08707f
C24860 a_31260_19975# VPWR 0.31436f
C24861 a_66652_1159# VPWR 0.3289f
C24862 a_1828_9096# VPWR 0.20348f
C24863 a_3620_5960# VPWR 0.22347f
C24864 a_67548_1159# a_67460_1256# 0.28563f
C24865 _443_.D VPWR 0.468f
C24866 a_32604_18407# VPWR 0.29679f
C24867 a_39460_1636# a_39100_1592# 0.08663f
C24868 _452_.CLK a_31284_22020# 0.0012f
C24869 _397_.A1 a_52988_26680# 0.0107f
C24870 a_15460_31048# uio_oe[0] 0.00329f
C24871 a_40580_20452# _325_.A2 0.00242f
C24872 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I a_57940_20452# 0.07119f
C24873 _330_.A1 a_44961_27912# 0.15206f
C24874 a_44388_27912# _470_.D 0.00268f
C24875 _238_.ZN _247_.ZN 0.19973f
C24876 _257_.B a_60276_29032# 0.2304f
C24877 a_27676_1159# a_28124_1159# 0.0131f
C24878 a_58388_10664# a_58836_10664# 0.01328f
C24879 _255_.ZN _243_.ZN 0.00322f
C24880 a_38772_28292# VPWR 0.00943f
C24881 a_35008_27533# a_35216_27533# 0.00372f
C24882 a_20420_24776# a_20508_23111# 0.00151f
C24883 _416_.A1 _408_.ZN 0.00561f
C24884 a_1916_26680# a_1916_26247# 0.05841f
C24885 _381_.A2 VPWR 2.10015f
C24886 a_28908_21976# VPWR 0.31547f
C24887 a_55788_25112# a_55788_24679# 0.05841f
C24888 _268_.A2 _258_.I 0.12155f
C24889 a_22636_28248# VPWR 0.33306f
C24890 _397_.A1 _398_.C 0.11635f
C24891 _325_.A2 a_37772_19759# 0.00122f
C24892 a_46716_2727# VPWR 0.31605f
C24893 a_34260_29860# VPWR 0.01552f
C24894 a_67572_13800# VPWR 0.20595f
C24895 a_57380_2824# a_57468_1159# 0.0027f
C24896 a_30052_21640# a_30500_21640# 0.01328f
C24897 a_35504_18955# a_36384_19369# 0.00306f
C24898 a_60156_27815# _244_.Z 0.00154f
C24899 a_14796_26247# a_14708_26344# 0.28563f
C24900 _270_.A2 ui_in[2] 0.00265f
C24901 _237_.A1 ui_in[3] 0.08127f
C24902 a_31620_15368# a_32068_15368# 0.01328f
C24903 _330_.A1 uo_out[7] 0.0021f
C24904 a_15132_29816# VPWR 0.29679f
C24905 a_20003_29611# uio_out[6] 0.55731f
C24906 a_27028_22020# a_27004_21543# 0.00172f
C24907 a_47612_10567# VPWR 0.29679f
C24908 a_23084_21976# a_23196_21543# 0.02634f
C24909 a_33500_15271# a_33412_15368# 0.28563f
C24910 _251_.A1 _243_.A1 0.00828f
C24911 _474_.Q _476_.Q 0.84024f
C24912 a_33724_23111# VPWR 0.35211f
C24913 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN 0.00195f
C24914 a_35068_15271# a_35516_15271# 0.0131f
C24915 a_47552_19715# a_48776_20204# 0.00164f
C24916 a_62196_26724# a_62644_26724# 0.01328f
C24917 a_2276_22020# a_2724_22020# 0.01328f
C24918 a_47612_2727# a_47524_2824# 0.28563f
C24919 a_54892_19975# a_54804_20072# 0.28563f
C24920 a_67460_17316# a_67908_17316# 0.01328f
C24921 a_63876_17316# a_63516_17272# 0.08717f
C24922 _275_.A2 uio_in[1] 0.00112f
C24923 _436_.ZN _432_.ZN 0.1883f
C24924 _261_.ZN _435_.ZN 0.32955f
C24925 _480_.Q _330_.A1 0.00224f
C24926 a_3708_8999# a_4156_8999# 0.0131f
C24927 a_60828_26680# a_60964_26344# 0.00168f
C24928 a_28484_1256# a_28932_1256# 0.01328f
C24929 a_19724_23544# a_20172_23544# 0.01288f
C24930 a_4940_7431# a_5388_7431# 0.01222f
C24931 a_64412_5863# a_64860_5863# 0.0131f
C24932 a_67212_20408# a_67348_20072# 0.00168f
C24933 a_3708_13703# a_4068_13800# 0.08717f
C24934 a_65308_4295# a_65756_4295# 0.0131f
C24935 a_7516_2727# a_7964_2727# 0.0131f
C24936 a_57580_13703# a_58028_13703# 0.01288f
C24937 _267_.A2 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.05971f
C24938 a_66787_30600# a_67741_30600# 0.00337f
C24939 a_39572_16936# a_39772_15271# 0.00119f
C24940 a_28820_20452# a_28908_20408# 0.28563f
C24941 _311_.A2 a_36548_21640# 0.00131f
C24942 _324_.B a_43400_18909# 0.00148f
C24943 a_23420_1592# VPWR 0.32982f
C24944 _419_.Z a_50212_20452# 0.0071f
C24945 a_64996_12612# a_65084_12568# 0.28563f
C24946 a_11091_30644# a_11548_30951# 0.00916f
C24947 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN 0.0102f
C24948 a_2812_23544# a_2812_23111# 0.05841f
C24949 _325_.A1 _325_.ZN 0.31488f
C24950 a_57580_17272# a_57468_16839# 0.02634f
C24951 _362_.B a_35008_27533# 0.00906f
C24952 a_54332_20408# a_54444_19975# 0.02634f
C24953 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN _231_.I 0.0021f
C24954 a_62084_18504# a_62532_18504# 0.01328f
C24955 a_52540_11000# a_53124_11044# 0.01675f
C24956 _296_.ZN a_41056_30669# 0.00543f
C24957 a_932_15368# a_932_14180# 0.05841f
C24958 _304_.A1 _324_.B 0.00883f
C24959 a_43828_16936# a_44276_16936# 0.01328f
C24960 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN a_58924_18840# 0.00117f
C24961 a_45956_1636# a_46404_1636# 0.01328f
C24962 a_42372_1636# a_42460_1592# 0.28563f
C24963 _452_.D a_42404_17433# 0.00159f
C24964 a_3708_26680# a_4156_26680# 0.0131f
C24965 a_24952_29032# VPWR 0.30737f
C24966 _362_.ZN a_32916_29860# 0.01306f
C24967 a_31844_2824# a_31708_1592# 0.00154f
C24968 a_4604_20408# VPWR 0.33016f
C24969 _255_.ZN _258_.ZN 0.11893f
C24970 _452_.CLK a_33636_23208# 0.00961f
C24971 a_48956_12568# VPWR 0.33349f
C24972 a_21424_25987# a_21052_26031# 0.10745f
C24973 a_20496_26344# a_22059_26399# 0.41635f
C24974 a_8548_2824# a_8996_2824# 0.01328f
C24975 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN 0.10373f
C24976 a_6172_29383# a_6532_29480# 0.08717f
C24977 _452_.CLK a_37964_18191# 0.026f
C24978 _397_.A1 _393_.A3 0.06765f
C24979 a_2812_28248# a_2812_27815# 0.05841f
C24980 a_44476_15271# a_44836_15368# 0.08717f
C24981 a_1828_10664# VPWR 0.20348f
C24982 _416_.A2 a_47164_18407# 0.02579f
C24983 a_31396_23208# VPWR 0.20622f
C24984 a_20379_29977# _375_.Z 0.02592f
C24985 _459_.CLK a_17786_29480# 0.00484f
C24986 a_14796_28248# a_15244_28248# 0.01255f
C24987 a_16052_28292# a_16140_28248# 0.28563f
C24988 _419_.Z a_51240_19624# 0.01376f
C24989 _447_.Q a_43126_24119# 0.00817f
C24990 a_67012_15748# VPWR 0.20622f
C24991 a_58588_2727# a_58948_2824# 0.08717f
C24992 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN a_64412_29816# 0.00531f
C24993 _245_.I1 a_61836_25515# 0.62001f
C24994 a_42908_30951# a_43268_31048# 0.08717f
C24995 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN 0.00619f
C24996 a_62084_15368# a_62532_15368# 0.01328f
C24997 _459_.Q a_31372_23544# 0.00111f
C24998 a_45360_29977# VPWR 0.00204f
C24999 _441_.A2 _302_.Z 0.00303f
C25000 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I VPWR 0.73205f
C25001 a_27476_23588# a_27564_23544# 0.28563f
C25002 a_54356_18504# a_54804_18504# 0.01328f
C25003 _452_.CLK a_42596_27912# 0.0128f
C25004 a_18380_25112# a_18828_25112# 0.01288f
C25005 a_11236_1256# VPWR 0.21187f
C25006 a_1020_7864# VPWR 0.30073f
C25007 a_2812_4728# VPWR 0.30213f
C25008 a_17284_31048# VPWR 0.20981f
C25009 a_32156_18840# a_32156_18407# 0.05841f
C25010 a_54668_13703# a_54580_13800# 0.28563f
C25011 a_50772_16936# a_50748_15271# 0.00134f
C25012 a_34160_20523# _319_.ZN 0.24766f
C25013 a_1916_29383# VPWR 0.297f
C25014 _370_.B a_30596_28292# 0.00101f
C25015 a_28124_30600# _371_.ZN 0.03282f
C25016 a_41140_27912# a_41392_27165# 0.0031f
C25017 a_44028_27815# a_43564_27209# 0.00104f
C25018 a_41452_16839# a_41364_16936# 0.28563f
C25019 a_55252_25156# a_55340_25112# 0.28563f
C25020 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN 0.12206f
C25021 _327_.A2 _325_.ZN 0.06315f
C25022 a_37220_1636# VPWR 0.2085f
C25023 a_1828_16936# VPWR 0.20348f
C25024 a_4940_12135# a_5388_12135# 0.01222f
C25025 _474_.CLK _389_.ZN 0.0011f
C25026 a_39796_27912# VPWR 0.12977f
C25027 a_5412_1636# a_5500_1592# 0.28563f
C25028 a_1468_1592# a_1916_1592# 0.01288f
C25029 a_58063_30644# a_58116_30344# 0.00171f
C25030 a_38576_22504# VPWR 0.81136f
C25031 a_55228_28248# a_55228_27815# 0.05841f
C25032 a_3620_17316# a_3708_17272# 0.28563f
C25033 _229_.I a_60404_28292# 0.0095f
C25034 a_59844_11044# a_59484_11000# 0.08707f
C25035 a_21540_1636# a_21404_1159# 0.00168f
C25036 a_17596_1592# a_17596_1159# 0.05841f
C25037 a_62420_12232# a_62508_10567# 0.00151f
C25038 a_55340_25112# VPWR 0.29679f
C25039 a_58836_17316# a_58924_17272# 0.28563f
C25040 a_60940_15704# a_60964_14180# 0.00144f
C25041 _424_.A2 a_53348_18884# 0.00803f
C25042 a_44459_18559# a_44744_18559# 0.00277f
C25043 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_56720_26344# 0.00164f
C25044 _237_.A1 _267_.A2 0.06187f
C25045 a_49852_1159# a_50524_1159# 0.00544f
C25046 _470_.Q a_44571_26841# 0.00257f
C25047 _475_.Q _419_.Z 0.10151f
C25048 a_61724_18407# VPWR 0.32947f
C25049 a_63428_18884# a_63516_18840# 0.28563f
C25050 a_67460_18884# a_67908_18884# 0.01328f
C25051 a_4964_25156# VPWR 0.21167f
C25052 _229_.I a_61689_29860# 0.00149f
C25053 a_3260_27815# a_3172_27912# 0.28563f
C25054 a_24652_20408# VPWR 0.31143f
C25055 a_51988_24776# a_51332_24372# 0.01565f
C25056 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I a_67684_21640# 0.05286f
C25057 _436_.ZN _260_.A1 0.00444f
C25058 _311_.A2 _444_.D 0.1274f
C25059 _441_.ZN _261_.ZN 0.17354f
C25060 a_62756_12612# VPWR 0.20595f
C25061 a_62560_25112# a_62864_25156# 0.00736f
C25062 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I a_62404_25156# 0.00138f
C25063 a_2364_15704# a_2812_15704# 0.0131f
C25064 _417_.A2 _421_.B 0.01169f
C25065 _399_.A2 _475_.Q 0.00594f
C25066 a_4964_15748# a_4604_15704# 0.08674f
C25067 a_60852_15748# VPWR 0.14831f
C25068 a_36636_15704# a_36772_15368# 0.00168f
C25069 a_54020_15368# a_54468_15368# 0.01328f
C25070 _379_.Z _467_.D 0.39119f
C25071 _311_.A2 a_34939_23705# 0.00992f
C25072 a_38564_15748# a_38428_15271# 0.00168f
C25073 a_63316_10664# VPWR 0.20641f
C25074 a_54892_24679# clk 0.01873f
C25075 a_64412_8999# a_64772_9096# 0.08717f
C25076 _350_.A2 _287_.A1 0.04083f
C25077 a_66204_5863# a_66564_5960# 0.08717f
C25078 a_55900_15271# a_55812_15368# 0.28563f
C25079 a_65308_7431# a_65668_7528# 0.08717f
C25080 a_31372_21976# a_31396_21640# 0.00172f
C25081 a_67100_4295# a_67460_4392# 0.08717f
C25082 a_22748_21543# a_22772_20452# 0.0016f
C25083 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN 0.00275f
C25084 a_37584_29123# VPWR 0.70601f
C25085 a_36772_15368# VPWR 0.20348f
C25086 _457_.D a_24788_23588# 0.00167f
C25087 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_55788_24679# 0.00379f
C25088 _448_.Q _304_.ZN 0.02866f
C25089 _386_.A4 _403_.ZN 0.00109f
C25090 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I VPWR 0.83726f
C25091 a_58700_16839# VPWR 0.34536f
C25092 a_20620_21976# a_21068_21976# 0.01288f
C25093 _243_.A1 a_58020_27508# 0.22382f
C25094 vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I 0.00413f
C25095 a_3620_14180# a_3708_14136# 0.28563f
C25096 a_38764_16839# a_39212_16839# 0.01288f
C25097 a_40220_15271# VPWR 0.32938f
C25098 a_28012_23544# a_27924_22020# 0.00151f
C25099 a_64412_17272# VPWR 0.31695f
C25100 _268_.A2 _255_.ZN 0.00197f
C25101 _432_.ZN _439_.ZN 0.15673f
C25102 a_33636_1256# VPWR 0.20713f
C25103 VPWR uio_oe[1] 0.09161f
C25104 a_50884_1256# a_51332_1256# 0.01328f
C25105 a_52920_22760# _427_.B2 0.03151f
C25106 a_29916_2727# a_30364_2727# 0.0131f
C25107 a_65420_13703# a_65780_13800# 0.08717f
C25108 a_49292_13703# a_49316_12612# 0.0016f
C25109 a_51444_13800# a_51892_13800# 0.01328f
C25110 _346_.B a_21652_29480# 0.00885f
C25111 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I a_59284_14180# 0.02898f
C25112 a_60909_30600# ui_in[1] 0.0072f
C25113 a_33148_25641# a_33492_25273# 0.00275f
C25114 a_17372_30951# VPWR 0.31184f
C25115 _395_.A2 a_50084_24328# 0.03711f
C25116 a_67348_18504# VPWR 0.20595f
C25117 _359_.B _362_.ZN 0.16898f
C25118 _365_.ZN _294_.ZN 0.00327f
C25119 a_52204_16839# a_52564_16936# 0.08717f
C25120 a_43356_1592# VPWR 0.29679f
C25121 a_44632_30206# a_45012_29816# 0.49319f
C25122 a_55476_10664# a_55588_9476# 0.02666f
C25123 a_51644_1592# a_51780_1256# 0.00168f
C25124 a_11324_1159# a_11236_1256# 0.28563f
C25125 a_1916_12135# a_1828_12232# 0.28563f
C25126 a_48756_16936# VPWR 0.20885f
C25127 a_8188_1592# a_8860_1592# 0.00544f
C25128 _452_.CLK _442_.ZN 0.02537f
C25129 a_26668_23544# a_26556_23111# 0.02634f
C25130 a_6844_29816# a_7292_29816# 0.01288f
C25131 a_56484_29480# VPWR 0.17205f
C25132 a_28054_30196# _349_.A4 0.0026f
C25133 a_33412_17316# a_33500_17272# 0.28563f
C25134 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I 0.05466f
C25135 _424_.A2 a_45156_21236# 0.00194f
C25136 a_36996_17316# a_37444_17316# 0.01328f
C25137 a_49092_15368# a_48956_14136# 0.00154f
C25138 _470_.D a_43440_26841# 0.00165f
C25139 a_52092_1592# a_52540_1592# 0.01288f
C25140 _424_.A1 a_51240_19624# 0.00503f
C25141 a_66340_11044# a_66788_11044# 0.01328f
C25142 a_63204_11044# a_62844_11000# 0.08707f
C25143 a_39536_26795# a_40464_27165# 1.16391f
C25144 a_13700_2824# VPWR 0.20348f
C25145 a_30388_28776# uo_out[6] 0.02326f
C25146 a_63852_23111# vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I 0.00134f
C25147 _275_.ZN _390_.ZN 0.00151f
C25148 a_36636_26680# VPWR 0.29679f
C25149 a_17484_23111# a_17932_23111# 0.0131f
C25150 _384_.A3 _417_.A2 0.34319f
C25151 _330_.A1 a_34396_21543# 0.00957f
C25152 _459_.CLK a_19076_26344# 0.00688f
C25153 _437_.A1 a_37516_27599# 0.00707f
C25154 a_5052_6296# a_4964_4772# 0.00151f
C25155 a_67236_15368# VPWR 0.20348f
C25156 _455_.Q a_22352_25987# 0.17593f
C25157 a_22636_25112# VPWR 0.3185f
C25158 _223_.I _370_.B 0.17678f
C25159 _325_.A2 _331_.ZN 0.03833f
C25160 a_58476_18840# vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I 0.00268f
C25161 a_34756_15748# a_34396_15704# 0.08707f
C25162 a_49740_12135# VPWR 0.32073f
C25163 _358_.A3 _459_.D 0.04327f
C25164 a_30724_2824# a_31396_2824# 0.00347f
C25165 _311_.A2 a_34715_22137# 0.01264f
C25166 a_56036_28292# vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I 0.00236f
C25167 a_45372_15704# a_45372_15271# 0.05841f
C25168 a_2812_24679# VPWR 0.30213f
C25169 a_41776_20072# VPWR 0.01501f
C25170 a_21316_21640# a_21292_20408# 0.0016f
C25171 a_52639_30644# _276_.A2 0.021f
C25172 a_53212_29816# ui_in[7] 0.00182f
C25173 _300_.ZN a_39684_20452# 0.13599f
C25174 a_32516_15748# VPWR 0.20348f
C25175 a_2724_9476# a_3172_9476# 0.01328f
C25176 a_27924_22020# a_27564_21976# 0.08707f
C25177 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN 0.84533f
C25178 _303_.ZN a_39772_20408# 0.00323f
C25179 a_51556_14180# a_52004_14180# 0.01328f
C25180 a_47972_14180# a_48060_14136# 0.28563f
C25181 _325_.A1 _438_.ZN 0.52658f
C25182 a_54332_18840# a_54780_18840# 0.01222f
C25183 _384_.ZN _404_.A1 0.14795f
C25184 a_43916_16839# VPWR 0.31223f
C25185 _350_.A2 a_28000_29480# 0.03913f
C25186 a_49652_16936# a_49540_15748# 0.02666f
C25187 a_52360_26355# a_52848_25987# 0.8399f
C25188 _325_.A1 a_41572_20072# 0.00162f
C25189 a_56036_1256# VPWR 0.20348f
C25190 a_46180_13800# a_46180_12612# 0.05841f
C25191 a_65980_14136# a_65892_12612# 0.00151f
C25192 a_44752_18147# a_45172_17316# 0.01617f
C25193 a_34396_17272# VPWR 0.33851f
C25194 _231_.ZN _231_.I 0.47744f
C25195 a_62868_10664# a_62756_9476# 0.02666f
C25196 a_61076_10664# a_61052_9432# 0.0016f
C25197 a_35088_20893# _319_.A2 0.00271f
C25198 a_22300_1159# a_22660_1256# 0.08717f
C25199 a_66316_12135# a_66764_12135# 0.0131f
C25200 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I _249_.A2 0.04177f
C25201 a_52428_12135# a_52788_12232# 0.08707f
C25202 a_57156_1636# VPWR 0.2129f
C25203 a_25324_23544# a_25348_23208# 0.00172f
C25204 a_15492_29480# a_16164_29480# 0.00347f
C25205 _402_.A1 _421_.A1 0.5219f
C25206 a_15132_1592# a_15580_1592# 0.01288f
C25207 _325_.B a_42896_18504# 0.07421f
C25208 a_14148_29860# a_13788_29816# 0.08707f
C25209 _358_.A3 a_33524_24776# 0.00157f
C25210 a_36100_2824# VPWR 0.20815f
C25211 a_59396_1636# a_59036_1592# 0.08707f
C25212 a_58911_30644# _255_.I 0.00557f
C25213 a_53908_25156# clk 0.00151f
C25214 _459_.CLK a_16500_27912# 0.00496f
C25215 _370_.B a_32508_30644# 0.00878f
C25216 a_20508_24679# a_20420_24776# 0.28563f
C25217 a_2276_24776# a_2724_24776# 0.01328f
C25218 a_16588_23111# a_16500_23208# 0.28563f
C25219 _371_.A1 a_29184_25597# 0.00114f
C25220 _455_.Q a_20308_27912# 0.00231f
C25221 a_3260_9432# VPWR 0.30487f
C25222 a_66116_9096# a_66564_9096# 0.01328f
C25223 a_45396_28292# _403_.ZN 0.00195f
C25224 a_67012_7528# a_67460_7528# 0.01328f
C25225 a_48956_14136# VPWR 0.33349f
C25226 _316_.A3 a_35044_21640# 0.00294f
C25227 _412_.A1 a_51332_24372# 0.17246f
C25228 _251_.A1 a_62732_26680# 0.02325f
C25229 _400_.ZN a_45232_25987# 0.04262f
C25230 _427_.A2 _476_.Q 0.00631f
C25231 a_1828_18504# a_2276_18504# 0.01328f
C25232 a_32604_18407# a_32964_18504# 0.08717f
C25233 a_56036_28292# vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.00201f
C25234 a_37556_23588# a_37644_23544# 0.28563f
C25235 _230_.I _250_.A2 0.50302f
C25236 _476_.Q a_51196_21543# 0.00312f
C25237 a_17148_29816# uio_out[7] 0.00127f
C25238 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_61948_27815# 0.01306f
C25239 _373_.A2 _349_.A4 0.02677f
C25240 _260_.A1 _439_.ZN 0.61557f
C25241 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.86475f
C25242 a_41252_15748# a_41700_15748# 0.01328f
C25243 a_3620_12232# VPWR 0.22347f
C25244 a_55956_25940# VPWR 0.56662f
C25245 a_16500_24776# VPWR 0.20348f
C25246 _475_.Q _416_.A2 0.01272f
C25247 a_41188_18840# a_41600_19376# 0.00705f
C25248 _422_.ZN _424_.ZN 0.0119f
C25249 a_2364_2727# a_2724_2824# 0.08717f
C25250 a_38652_15704# VPWR 0.33352f
C25251 a_4156_19975# a_4068_20072# 0.28563f
C25252 _334_.A1 _287_.A1 0.74467f
C25253 _436_.ZN _260_.A2 0.04951f
C25254 _287_.A2 _359_.B 0.03094f
C25255 a_44571_26841# a_44816_27209# 0.00232f
C25256 _451_.Q a_38971_18559# 0.01886f
C25257 a_47076_9476# a_47164_9432# 0.28563f
C25258 _324_.C a_44160_29123# 0.00196f
C25259 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_55588_28292# 0.03625f
C25260 _350_.A1 a_30160_30301# 0.06727f
C25261 _327_.A2 a_41572_20072# 0.00387f
C25262 _444_.D a_36660_23588# 0.00308f
C25263 uio_out[1] uio_out[0] 0.06083f
C25264 _265_.ZN a_42148_27912# 0.042f
C25265 _304_.B a_55676_27815# 0.00224f
C25266 a_3620_12612# a_3260_12568# 0.08717f
C25267 a_52316_2727# a_52764_2727# 0.0131f
C25268 a_53236_13800# a_53124_12612# 0.02666f
C25269 a_1020_12568# a_1468_12568# 0.0131f
C25270 a_61297_30300# vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I 0.00247f
C25271 _355_.ZN a_27760_25273# 0.00242f
C25272 a_29184_25597# a_30476_25112# 0.00295f
C25273 _424_.A2 _324_.B 1.01954f
C25274 _331_.ZN a_40244_18180# 0.01863f
C25275 a_46492_17272# VPWR 0.31945f
C25276 a_66428_1592# VPWR 0.33479f
C25277 a_67324_1592# a_67460_1256# 0.00168f
C25278 a_33724_1159# a_33636_1256# 0.28563f
C25279 a_22436_1636# a_22076_1592# 0.08707f
C25280 a_63404_12135# a_63316_12232# 0.28563f
C25281 _287_.A1 a_35156_29860# 0.00199f
C25282 a_1380_4392# a_1380_3204# 0.05841f
C25283 a_27004_21543# VPWR 0.34756f
C25284 a_17596_29816# _459_.CLK 0.02874f
C25285 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I _324_.C 0.04283f
C25286 a_20672_30301# a_22560_30288# 0.01012f
C25287 _416_.A1 _473_.Q 0.1188f
C25288 a_49092_17316# a_49540_17316# 0.01328f
C25289 a_17844_26344# a_17844_25156# 0.05841f
C25290 _459_.CLK a_24392_28248# 0.0321f
C25291 a_39536_23588# VPWR 0.01391f
C25292 _274_.ZN a_52964_29480# 0.01355f
C25293 a_53324_10567# a_53772_10567# 0.01288f
C25294 a_67324_11000# a_67212_10567# 0.02634f
C25295 a_64100_1636# a_63740_1592# 0.08717f
C25296 a_65892_1636# a_66340_1636# 0.01328f
C25297 _389_.ZN _393_.A3 0.62461f
C25298 a_58500_2824# VPWR 0.21417f
C25299 _428_.Z a_51332_24072# 0.0328f
C25300 a_56036_27912# vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.06797f
C25301 a_15156_23208# a_15604_23208# 0.01328f
C25302 a_27452_23111# a_27812_23208# 0.08707f
C25303 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I VPWR 0.87857f
C25304 _337_.ZN a_31964_28292# 0.01071f
C25305 _229_.I _248_.B1 0.24464f
C25306 _284_.ZN _437_.A1 0.01357f
C25307 a_53884_9432# VPWR 0.31143f
C25308 a_64548_14180# VPWR 0.21283f
C25309 a_21852_21543# a_22300_21543# 0.01288f
C25310 _336_.A2 a_28796_23111# 0.00239f
C25311 _324_.C a_43564_27209# 0.01446f
C25312 a_65332_12232# VPWR 0.21224f
C25313 _427_.B2 a_53003_22504# 0.00927f
C25314 _330_.A1 _313_.ZN 0.68931f
C25315 _409_.ZN _402_.A1 0.00623f
C25316 a_53124_2824# a_53572_2824# 0.01328f
C25317 a_36636_2727# a_36772_1636# 0.00154f
C25318 a_7180_30951# a_7204_29860# 0.0016f
C25319 _334_.A1 _293_.A2 0.89304f
C25320 _229_.I vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN 0.81868f
C25321 a_35616_24776# VPWR 1.11125f
C25322 a_3172_18884# VPWR 0.20993f
C25323 _311_.A2 _301_.Z 0.21257f
C25324 _412_.ZN clk 0.07953f
C25325 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_55588_27912# 0.00251f
C25326 a_13788_2727# a_13700_2824# 0.28563f
C25327 a_52316_15704# VPWR 0.32971f
C25328 _275_.A2 _275_.ZN 0.83882f
C25329 a_52316_9432# a_52900_9476# 0.01675f
C25330 _252_.ZN a_59620_27208# 0.04444f
C25331 _416_.A1 _475_.D 0.50641f
C25332 a_24080_25227# a_24340_23588# 0.00105f
C25333 a_59372_14136# a_59820_14136# 0.01255f
C25334 a_49316_14180# a_49292_13703# 0.00172f
C25335 a_45372_14136# a_45372_13703# 0.05841f
C25336 a_62508_23111# clk 0.00239f
C25337 a_1828_20452# a_1916_20408# 0.28563f
C25338 _384_.ZN a_48384_26724# 0.04949f
C25339 a_55676_27815# VPWR 0.29679f
C25340 _336_.Z a_29028_24072# 0.00183f
C25341 _392_.A2 _381_.Z 0.00364f
C25342 a_47972_12612# a_47612_12568# 0.08707f
C25343 a_21404_1159# VPWR 0.3289f
C25344 a_44700_1159# a_45060_1256# 0.08717f
C25345 a_60180_12232# a_60628_12232# 0.01328f
C25346 a_25348_1636# a_25436_1592# 0.28563f
C25347 a_28932_1636# a_29380_1636# 0.01328f
C25348 a_38316_20408# a_38764_20408# 0.01222f
C25349 a_24004_21640# VPWR 0.20614f
C25350 _352_.ZN a_25936_25597# 0.00296f
C25351 a_38584_28292# VPWR 0.31423f
C25352 a_64188_11000# a_64212_10664# 0.00172f
C25353 a_50636_10567# a_50548_10664# 0.28563f
C25354 _325_.ZN a_44756_19001# 0.00195f
C25355 _325_.A2 a_39324_19975# 0.00839f
C25356 a_48596_28292# VPWR 0.01382f
C25357 _424_.B1 a_50420_23233# 0.00175f
C25358 a_62868_23208# VPWR 0.20869f
C25359 a_55252_20072# vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN 0.00294f
C25360 a_32096_24419# a_33076_24776# 0.00702f
C25361 a_41392_27165# a_41476_26344# 0.00101f
C25362 a_21428_23588# VPWR 0.20622f
C25363 a_64860_9432# VPWR 0.30145f
C25364 a_20508_21543# a_20868_21640# 0.08707f
C25365 a_1468_2727# VPWR 0.29679f
C25366 a_51532_13703# VPWR 0.31431f
C25367 a_67100_6296# VPWR 0.29679f
C25368 a_40580_26344# VPWR 0.20512f
C25369 _337_.A3 a_25884_27815# 0.01608f
C25370 _441_.A3 a_39587_24372# 0.00201f
C25371 _455_.Q a_27004_27815# 0.00229f
C25372 _447_.Q _323_.A3 0.01165f
C25373 a_35740_30951# uo_out[3] 0.00876f
C25374 _330_.A1 _316_.ZN 0.5656f
C25375 a_51332_15748# a_51420_15704# 0.28563f
C25376 a_46716_11000# VPWR 0.29679f
C25377 a_47388_15704# a_47836_15704# 0.01288f
C25378 _437_.ZN a_38575_24072# 0.00403f
C25379 a_29575_28293# VPWR 0.56551f
C25380 a_2276_26724# VPWR 0.20634f
C25381 _245_.Z a_61748_26724# 0.00743f
C25382 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62308_27912# 0.03753f
C25383 _250_.ZN a_60940_28248# 0.00779f
C25384 _237_.A1 _256_.A2 0.09942f
C25385 _345_.A2 a_22620_27599# 0.03425f
C25386 a_46044_30951# vgaringosc.workerclkbuff_notouch_.I 0.00613f
C25387 a_5300_26344# VPWR 0.21406f
C25388 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I a_57580_18407# 0.00168f
C25389 _452_.CLK _441_.ZN 0.00178f
C25390 a_24764_2727# a_25124_2824# 0.08717f
C25391 _473_.Q a_46389_21236# 0.00918f
C25392 _438_.A2 _430_.ZN 0.20518f
C25393 _350_.A2 a_29620_30345# 0.00122f
C25394 a_1916_28248# VPWR 0.297f
C25395 _260_.A2 _439_.ZN 0.07684f
C25396 a_58052_9476# a_58140_9432# 0.28563f
C25397 _393_.ZN a_44795_29535# 0.00156f
C25398 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I _250_.B 0.01085f
C25399 a_66788_14180# a_66876_14136# 0.28563f
C25400 a_49600_30180# uio_in[1] 0.00224f
C25401 a_17844_20452# a_17484_20408# 0.08717f
C25402 _336_.Z a_29356_21976# 0.00131f
C25403 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN a_63105_28293# 0.00356f
C25404 a_15692_20408# a_16140_20408# 0.0131f
C25405 _416_.A1 a_44500_25156# 0.0046f
C25406 a_54804_23588# a_54444_23544# 0.08717f
C25407 _258_.I a_56572_29383# 0.05977f
C25408 a_63616_31128# a_65084_30951# 0.0058f
C25409 a_54468_12612# a_54916_12612# 0.01328f
C25410 a_23084_29383# VPWR 0.33665f
C25411 a_3172_1636# VPWR 0.20993f
C25412 _397_.A2 a_47636_25940# 0.06444f
C25413 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN _248_.B1 0.01436f
C25414 _459_.CLK a_23644_29816# 0.0288f
C25415 a_55140_20452# VPWR 0.20962f
C25416 _433_.ZN a_40880_23588# 0.01051f
C25417 a_43804_1159# VPWR 0.29679f
C25418 _441_.ZN a_40316_23233# 0.00436f
C25419 a_56124_1159# a_56036_1256# 0.28563f
C25420 _416_.A1 _381_.Z 0.00334f
C25421 a_1380_11044# a_1468_11000# 0.28563f
C25422 _424_.A2 a_52024_20083# 0.02952f
C25423 a_47076_10664# a_47524_10664# 0.01328f
C25424 _467_.D a_15692_27815# 0.0048f
C25425 a_61164_10567# a_61524_10664# 0.08707f
C25426 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_59284_13800# 0.00157f
C25427 a_56708_1636# a_56572_1159# 0.00168f
C25428 a_16252_1159# a_16700_1159# 0.0131f
C25429 _474_.Q _397_.Z 0.793f
C25430 _260_.A1 _303_.ZN 0.10068f
C25431 _448_.Q _441_.B 0.00209f
C25432 _452_.Q a_40656_23588# 0.00147f
C25433 a_17508_2824# a_17508_1636# 0.05841f
C25434 a_55252_23588# a_55700_23588# 0.01328f
C25435 a_14796_21976# VPWR 0.30073f
C25436 a_42610_21812# VPWR 0.00514f
C25437 _365_.ZN a_36284_29167# 0.01143f
C25438 a_28820_24072# VPWR 0.30822f
C25439 a_19076_21640# a_19524_21640# 0.01328f
C25440 a_31484_21543# a_31396_21640# 0.28563f
C25441 a_23868_2727# VPWR 0.31605f
C25442 a_45284_13800# VPWR 0.22176f
C25443 _304_.B _427_.B2 0.29081f
C25444 a_62620_15271# a_63068_15271# 0.0131f
C25445 a_1020_29816# VPWR 0.30073f
C25446 a_19744_30301# uio_out[6] 0.00118f
C25447 _383_.ZN a_48596_28292# 0.0063f
C25448 a_54556_21543# a_54692_20452# 0.00154f
C25449 a_60380_11000# VPWR 0.34427f
C25450 _365_.ZN _362_.B 0.07746f
C25451 a_67908_15748# a_67772_15271# 0.00168f
C25452 a_2364_23111# VPWR 0.30029f
C25453 _230_.I a_59172_27912# 0.03404f
C25454 a_64412_29816# VPWR 0.33894f
C25455 _452_.Q a_42728_20452# 0.0087f
C25456 _325_.A1 a_40692_21640# 0.00331f
C25457 a_2724_27912# VPWR 0.20782f
C25458 a_66204_15704# a_66652_15704# 0.01255f
C25459 a_36188_2727# a_36100_2824# 0.28563f
C25460 a_63404_23111# a_63316_23208# 0.28563f
C25461 _383_.A2 _392_.A2 0.07588f
C25462 a_53348_18884# a_54244_18884# 0.0023f
C25463 _268_.A1 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.20966f
C25464 a_63292_9432# a_63740_9432# 0.0131f
C25465 a_16500_23588# a_16948_23588# 0.01328f
C25466 a_65220_7908# a_65668_7908# 0.01328f
C25467 a_17060_1256# a_17508_1256# 0.01328f
C25468 _290_.ZN a_34586_27912# 0.02369f
C25469 a_65220_4772# a_65308_4728# 0.28563f
C25470 a_67012_4772# a_67460_4772# 0.01328f
C25471 a_64324_6340# a_64412_6296# 0.28563f
C25472 a_66116_6340# a_66564_6340# 0.01328f
C25473 _363_.Z VPWR 1.83945f
C25474 _355_.C a_27140_26344# 0.00925f
C25475 a_46268_13703# a_46716_13703# 0.0131f
C25476 a_66116_3204# a_66204_3160# 0.28563f
C25477 _244_.Z a_59652_25640# 0.00507f
C25478 a_59036_26247# _231_.ZN 0.05994f
C25479 a_7516_29383# a_7964_29383# 0.0131f
C25480 a_9635_30644# a_10004_31048# 0.02397f
C25481 _246_.B2 _250_.ZN 0.01051f
C25482 _282_.ZN clkbuf_1_0__f_clk.I 0.00149f
C25483 a_9308_1592# VPWR 0.3289f
C25484 a_64212_13800# a_64300_12135# 0.00151f
C25485 a_31396_31048# VPWR 0.2323f
C25486 a_43716_31048# vgaringosc.workerclkbuff_notouch_.I 0.00544f
C25487 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_61524_23208# 0.05202f
C25488 a_66204_1159# VPWR 0.34855f
C25489 a_36960_27912# VPWR 1.10363f
C25490 a_67100_1159# a_67460_1256# 0.08674f
C25491 a_1380_9096# VPWR 0.20348f
C25492 a_30812_19975# VPWR 0.32017f
C25493 a_7204_1636# a_7068_1159# 0.00168f
C25494 a_3260_1592# a_3260_1159# 0.05841f
C25495 a_35068_1592# a_35516_1592# 0.01288f
C25496 a_39012_1636# a_39100_1592# 0.28563f
C25497 a_37084_25112# a_37532_25112# 0.012f
C25498 a_3172_5960# VPWR 0.20993f
C25499 a_45732_11044# a_45820_11000# 0.28563f
C25500 a_49316_11044# a_49764_11044# 0.01328f
C25501 a_32516_16936# a_32964_16936# 0.01328f
C25502 _409_.ZN _424_.B1 0.08202f
C25503 a_32156_18407# VPWR 0.29679f
C25504 _399_.ZN _475_.Q 0.01011f
C25505 a_40132_20452# _325_.A2 0.00208f
C25506 a_43296_28733# a_43936_27165# 0.00107f
C25507 _330_.ZN a_37892_17316# 0.02213f
C25508 a_28460_21976# VPWR 0.31547f
C25509 _384_.ZN _399_.A2 0.17813f
C25510 a_22996_28292# VPWR 0.20521f
C25511 a_36432_19325# a_37067_19001# 0.02112f
C25512 a_35504_18955# a_35892_19369# 0.00393f
C25513 a_43804_30951# a_44252_30951# 0.0131f
C25514 _448_.Q _300_.A2 0.69787f
C25515 _249_.A2 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN 0.01254f
C25516 a_67124_13800# VPWR 0.20595f
C25517 a_33812_29860# VPWR 0.0179f
C25518 _427_.B2 VPWR 0.85102f
C25519 a_46044_2727# VPWR 0.33981f
C25520 _441_.A2 a_43750_23544# 0.01487f
C25521 hold2.Z _452_.Q 0.01963f
C25522 _304_.B _400_.ZN 0.6845f
C25523 a_14684_29816# VPWR 0.29679f
C25524 a_64884_16936# a_64860_15704# 0.0016f
C25525 a_47164_10567# VPWR 0.29679f
C25526 a_33052_15271# a_33412_15368# 0.08717f
C25527 _327_.A2 a_40692_21640# 0.00476f
C25528 a_33276_23111# VPWR 0.32289f
C25529 _379_.A2 _459_.CLK 0.00603f
C25530 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN a_58836_17316# 0.00102f
C25531 _274_.ZN _274_.A1 0.46361f
C25532 _352_.A2 _355_.B 1.1419f
C25533 a_1380_28292# a_1828_28292# 0.01328f
C25534 a_47164_2727# a_47524_2824# 0.08717f
C25535 _325_.ZN VPWR 0.37449f
C25536 a_50436_30689# uio_in[1] 0.49261f
C25537 a_63428_17316# a_63516_17272# 0.28563f
C25538 a_54444_19975# a_54804_20072# 0.08674f
C25539 a_31920_29480# a_33776_29123# 0.02307f
C25540 a_32848_29123# a_33483_29535# 0.02112f
C25541 _304_.B uo_out[3] 0.44117f
C25542 a_1828_16936# a_1828_15748# 0.05841f
C25543 _349_.A4 a_25867_26841# 0.00175f
C25544 _459_.Q a_33188_25940# 0.00789f
C25545 a_67436_18407# a_67884_18407# 0.012f
C25546 a_15156_25156# a_15604_25156# 0.01328f
C25547 a_66652_9432# a_66652_8999# 0.05841f
C25548 _284_.ZN a_43492_27912# 0.03769f
C25549 a_66787_30600# a_67117_30600# 0.53809f
C25550 _358_.A3 _359_.ZN 0.35295f
C25551 a_3708_13703# a_3620_13800# 0.28563f
C25552 a_26668_20408# a_27116_20408# 0.0131f
C25553 a_28820_20452# a_28460_20408# 0.08717f
C25554 _325_.ZN a_44364_17272# 0.0036f
C25555 _416_.A1 _383_.A2 0.05987f
C25556 a_64772_18504# a_64772_17316# 0.05841f
C25557 a_54356_24776# a_54356_23588# 0.05841f
C25558 a_5388_16839# a_5300_16936# 0.28563f
C25559 a_46984_23588# _397_.Z 0.24544f
C25560 a_37308_1592# a_37444_1256# 0.00168f
C25561 _419_.Z a_49068_20408# 0.39284f
C25562 a_22972_1592# VPWR 0.3289f
C25563 a_64996_12612# a_64636_12568# 0.08707f
C25564 a_61052_12568# a_61500_12568# 0.01288f
C25565 a_4964_23588# a_4940_23111# 0.00172f
C25566 _438_.A2 _441_.A3 0.02513f
C25567 _324_.C _392_.A2 0.5444f
C25568 _325_.A1 a_43784_19369# 0.03562f
C25569 _470_.Q _397_.A4 1.39951f
C25570 a_51444_12232# a_51532_10567# 0.00151f
C25571 a_42372_1636# a_42012_1592# 0.08707f
C25572 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN a_59708_23111# 0.00114f
C25573 a_24304_29480# VPWR 0.01383f
C25574 a_38428_1159# a_39100_1159# 0.00544f
C25575 _346_.B a_20396_27815# 0.10696f
C25576 a_4156_20408# VPWR 0.30552f
C25577 _452_.CLK a_33188_23208# 0.02982f
C25578 a_932_2824# VPWR 0.22176f
C25579 a_48508_12568# VPWR 0.29679f
C25580 a_63092_16936# a_63540_16936# 0.01328f
C25581 a_20496_26344# a_21052_26031# 0.8399f
C25582 a_6172_29383# a_6084_29480# 0.28563f
C25583 _251_.A1 _250_.C 0.04343f
C25584 a_42596_15368# a_43044_15368# 0.01328f
C25585 _452_.CLK a_38336_18147# 0.01371f
C25586 _400_.ZN VPWR 0.5809f
C25587 a_4964_28292# a_4940_27815# 0.00172f
C25588 a_1380_10664# VPWR 0.20348f
C25589 a_44476_15271# a_44388_15368# 0.28563f
C25590 a_30948_23208# VPWR 0.20622f
C25591 a_35816_21192# a_36204_21327# 0.00334f
C25592 _324_.C a_50532_24072# 0.00928f
C25593 _257_.B _252_.B 0.00609f
C25594 a_58164_18504# a_58028_17272# 0.00154f
C25595 a_46044_15271# a_46492_15271# 0.0131f
C25596 _375_.Z _455_.Q 0.00125f
C25597 _255_.I _243_.A1 0.11708f
C25598 a_16052_28292# a_15692_28248# 0.0869f
C25599 a_17396_22020# a_17844_22020# 0.01328f
C25600 a_58588_2727# a_58500_2824# 0.28563f
C25601 _419_.Z a_48776_20204# 0.00146f
C25602 a_66564_15748# VPWR 0.20904f
C25603 a_42908_30951# a_42820_31048# 0.28563f
C25604 _231_.I clk 0.04465f
C25605 VPWR uo_out[3] 0.87345f
C25606 a_36548_21640# a_36996_21640# 0.01328f
C25607 a_2364_16839# a_2812_16839# 0.0131f
C25608 a_62308_26344# a_61836_25515# 0.00201f
C25609 _358_.A3 a_35552_27216# 0.00152f
C25610 a_35540_16936# a_35652_15748# 0.02666f
C25611 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I a_61300_16936# 0.00103f
C25612 a_62420_22020# VPWR 0.14846f
C25613 a_24004_23208# a_24092_21543# 0.00151f
C25614 a_10788_1256# VPWR 0.20914f
C25615 a_4964_7908# VPWR 0.21167f
C25616 a_16164_31048# VPWR 0.23282f
C25617 a_39460_1256# a_39908_1256# 0.01328f
C25618 a_27476_23588# a_27116_23544# 0.0869f
C25619 a_23980_23544# a_24428_23544# 0.0131f
C25620 a_2364_4728# VPWR 0.30029f
C25621 a_21876_25156# a_22548_25156# 0.00347f
C25622 a_1468_29383# VPWR 0.29679f
C25623 a_18492_2727# a_18940_2727# 0.0131f
C25624 a_54220_13703# a_54580_13800# 0.08707f
C25625 a_29828_26344# _358_.A2 0.08881f
C25626 a_27668_31048# _371_.ZN 0.00155f
C25627 _370_.B a_29575_28293# 0.10406f
C25628 a_1916_17272# a_1916_16839# 0.05841f
C25629 a_41004_16839# a_41364_16936# 0.08707f
C25630 a_55252_25156# a_54892_25112# 0.0869f
C25631 a_47972_10664# a_47972_9476# 0.05841f
C25632 _327_.A2 a_43784_19369# 0.00344f
C25633 _284_.A2 a_44340_26183# 0.02644f
C25634 _251_.A1 _245_.I1 0.32225f
C25635 _311_.A2 _439_.ZN 0.10268f
C25636 a_1380_16936# VPWR 0.20348f
C25637 a_36772_1636# VPWR 0.2085f
C25638 a_35660_27508# VPWR 0.00417f
C25639 a_5412_1636# a_5052_1592# 0.08707f
C25640 hold1.Z _324_.B 0.08075f
C25641 a_18828_23544# a_18716_23111# 0.02634f
C25642 a_3620_29860# a_4068_29860# 0.01328f
C25643 _384_.ZN a_49316_23588# 0.00494f
C25644 a_45904_30180# _393_.ZN 0.23284f
C25645 a_1020_17272# a_1468_17272# 0.0131f
C25646 a_3620_17316# a_3260_17272# 0.08717f
C25647 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I VPWR 0.806f
C25648 _370_.ZN a_28000_29480# 0.02475f
C25649 a_55452_11000# a_55900_11000# 0.01288f
C25650 a_59396_11044# a_59484_11000# 0.28563f
C25651 a_48868_1636# a_49316_1636# 0.01328f
C25652 a_54356_16936# a_54804_16936# 0.01328f
C25653 _352_.A2 a_25643_25273# 0.07269f
C25654 _416_.A1 _324_.C 3.36223f
C25655 a_54892_25112# VPWR 0.29679f
C25656 a_58836_17316# a_58476_17272# 0.08674f
C25657 a_2724_20072# a_2724_18884# 0.05841f
C25658 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_56368_26344# 0.00167f
C25659 _371_.A2 VPWR 2.96303f
C25660 a_46628_18504# a_46604_16839# 0.00131f
C25661 _470_.Q a_44864_27165# 0.17715f
C25662 a_63428_18884# a_63068_18840# 0.08717f
C25663 a_4516_25156# VPWR 0.20862f
C25664 a_17036_27815# a_17484_27815# 0.0131f
C25665 a_2812_27815# a_3172_27912# 0.08717f
C25666 a_51540_24776# a_51332_24372# 0.02745f
C25667 a_24204_20408# VPWR 0.31143f
C25668 a_37532_25112# _444_.D 0.0256f
C25669 a_57468_16839# vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN 0.00564f
C25670 a_62560_25112# a_62404_25156# 0.00399f
C25671 a_61836_25515# a_62864_25156# 0.00128f
C25672 a_4516_15748# a_4604_15704# 0.28563f
C25673 _416_.A1 _416_.ZN 0.83487f
C25674 a_62308_12612# VPWR 0.20595f
C25675 _284_.ZN a_43600_25640# 0.00176f
C25676 a_19300_2824# a_19972_2824# 0.00347f
C25677 a_17148_29383# _467_.D 0.01468f
C25678 VPWR uio_in[1] 0.5508f
C25679 _304_.B _438_.ZN 0.42423f
C25680 _311_.A2 a_35232_24029# 0.02731f
C25681 a_55452_15271# a_55812_15368# 0.08717f
C25682 vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN a_56684_17272# 0.00643f
C25683 a_65308_7431# a_65220_7528# 0.28563f
C25684 a_62868_10664# VPWR 0.20641f
C25685 a_64412_8999# a_64324_9096# 0.28563f
C25686 a_54444_24679# clk 0.01873f
C25687 a_67100_4295# a_67012_4392# 0.28563f
C25688 a_66204_5863# a_66116_5960# 0.28563f
C25689 _284_.B _474_.Q 0.03191f
C25690 a_37291_29535# VPWR 0.36874f
C25691 a_36324_15368# VPWR 0.20348f
C25692 a_58252_16839# VPWR 0.38006f
C25693 _350_.A1 _352_.A2 1.17322f
C25694 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I 0.24216f
C25695 uio_oe[2] uio_oe[1] 0.07417f
C25696 a_39772_15271# VPWR 0.32938f
C25697 a_1020_14136# a_1468_14136# 0.0131f
C25698 a_3620_14180# a_3260_14136# 0.08717f
C25699 a_42484_16936# a_42596_15748# 0.02666f
C25700 a_38676_16936# a_38652_15704# 0.0016f
C25701 a_63964_17272# VPWR 0.31389f
C25702 a_932_7528# VPWR 0.22176f
C25703 a_33188_1256# VPWR 0.2051f
C25704 a_27328_25227# _355_.ZN 0.24767f
C25705 a_65420_13703# a_65332_13800# 0.28563f
C25706 a_33948_17272# a_33948_16839# 0.05841f
C25707 a_16916_31048# VPWR 0.35948f
C25708 a_37892_17316# a_37868_16839# 0.00172f
C25709 a_60285_30600# ui_in[1] 0.00257f
C25710 a_52204_16839# a_52116_16936# 0.28563f
C25711 _474_.CLK vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.02904f
C25712 _268_.A2 _267_.A1 0.03692f
C25713 a_4068_23208# a_4068_22020# 0.05841f
C25714 a_66900_18504# VPWR 0.20595f
C25715 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I a_51457_29861# 0.02819f
C25716 a_42908_1592# VPWR 0.31296f
C25717 a_10876_1159# a_11236_1256# 0.08717f
C25718 a_48308_16936# VPWR 0.20703f
C25719 a_44632_30206# a_43916_29816# 0.00341f
C25720 a_4068_29480# a_4740_29480# 0.00347f
C25721 a_55116_12135# a_55564_12135# 0.01288f
C25722 a_1468_12135# a_1828_12232# 0.08717f
C25723 a_11908_1636# a_12356_1636# 0.01328f
C25724 _452_.CLK a_39536_26795# 0.05015f
C25725 a_23084_25112# a_23196_24679# 0.02634f
C25726 _417_.A2 _417_.Z 0.33329f
C25727 a_26427_29977# _349_.A4 0.03189f
C25728 a_33412_17316# a_33052_17272# 0.08707f
C25729 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN a_64188_27815# 0.05037f
C25730 a_62756_11044# a_62844_11000# 0.28563f
C25731 _231_.I a_59260_23544# 0.00693f
C25732 _474_.CLK _384_.A1 0.01977f
C25733 a_13252_2824# VPWR 0.20348f
C25734 _330_.A1 _438_.A2 0.37716f
C25735 _250_.B vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN 0.02218f
C25736 a_63404_23111# vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I 0.00328f
C25737 _363_.Z _370_.B 0.25255f
C25738 a_36188_26680# VPWR 0.29533f
C25739 a_17484_24679# a_17932_24679# 0.0131f
C25740 _459_.CLK a_18628_26344# 0.00651f
C25741 a_60828_1159# a_61276_1159# 0.0131f
C25742 _437_.A1 a_37888_27555# 0.01923f
C25743 a_38576_22504# a_39796_22504# 0.00203f
C25744 _455_.Q a_22059_26399# 0.00106f
C25745 a_66788_15368# VPWR 0.20348f
C25746 a_1916_18407# a_2364_18407# 0.0131f
C25747 a_22996_25156# VPWR 0.20939f
C25748 _223_.I a_32240_31048# 0.01027f
C25749 a_31396_31048# _370_.B 0.00237f
C25750 a_49292_12135# VPWR 0.32402f
C25751 a_58028_18840# vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I 0.00135f
C25752 a_34308_15748# a_34396_15704# 0.28563f
C25753 _358_.A3 a_31732_25156# 0.07283f
C25754 a_22300_2727# a_22436_1636# 0.00154f
C25755 a_47972_18504# a_47836_17272# 0.00154f
C25756 a_51668_18504# a_51780_17316# 0.02666f
C25757 a_43788_29167# a_44132_29535# 0.00275f
C25758 _438_.ZN VPWR 0.97728f
C25759 _427_.A2 a_53300_23047# 0.04904f
C25760 _474_.Q _474_.D 0.13463f
C25761 a_2364_24679# VPWR 0.30029f
C25762 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_61612_23111# 0.00266f
C25763 a_41572_20072# VPWR 0.0072f
C25764 a_52639_30644# a_52871_31198# 0.00209f
C25765 a_52415_31220# _276_.A2 0.01923f
C25766 a_57132_17272# vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN 0.00199f
C25767 a_32068_15748# VPWR 0.20348f
C25768 _384_.ZN a_49212_26369# 0.00616f
C25769 _293_.A2 _234_.ZN 0.03579f
C25770 a_42460_20452# _328_.A2 0.00118f
C25771 _300_.ZN a_38676_20452# 0.0042f
C25772 _409_.ZN _407_.A1 0.58505f
C25773 _276_.A2 ui_in[7] 0.08937f
C25774 a_65072_29860# rst_n 0.43433f
C25775 _438_.ZN a_41012_23208# 0.01899f
C25776 a_45820_18407# a_46268_18407# 0.0131f
C25777 a_27476_22020# a_27564_21976# 0.28563f
C25778 _319_.A3 _448_.D 0.07782f
C25779 _452_.Q _448_.Q 0.1712f
C25780 a_23532_21976# a_23980_21976# 0.01288f
C25781 _285_.Z uo_out[2] 0.04235f
C25782 a_49292_16839# a_49740_16839# 0.012f
C25783 _243_.B2 a_58052_26724# 0.00379f
C25784 a_47972_14180# a_47612_14136# 0.08707f
C25785 _452_.CLK a_36188_17272# 0.00111f
C25786 _229_.I a_60740_26724# 0.00202f
C25787 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN 0.04773f
C25788 a_48708_29816# a_49496_30345# 0.02112f
C25789 a_43468_16839# VPWR 0.31366f
C25790 a_51956_26183# a_52744_26031# 0.02112f
C25791 a_55588_1256# VPWR 0.20348f
C25792 a_61860_1256# a_62308_1256# 0.01328f
C25793 a_40892_2727# a_41340_2727# 0.0131f
C25794 a_61972_13800# a_62420_13800# 0.01328f
C25795 a_44752_18147# a_44724_17316# 0.00687f
C25796 a_59955_30600# VPWR 0.3126f
C25797 a_21764_23208# a_21876_22020# 0.02666f
C25798 a_33948_17272# VPWR 0.30233f
C25799 a_56708_1636# VPWR 0.21139f
C25800 a_22300_1159# a_22212_1256# 0.28563f
C25801 a_52428_12135# a_52340_12232# 0.28563f
C25802 _402_.A1 a_45128_26031# 0.00323f
C25803 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN a_65072_29860# 0.015f
C25804 a_13700_29860# a_13788_29816# 0.28563f
C25805 a_9756_29816# a_10204_29816# 0.01288f
C25806 a_61836_26680# a_61836_25515# 0.00151f
C25807 _358_.A3 a_33076_24776# 0.00181f
C25808 a_35428_1636# a_35292_1159# 0.00168f
C25809 a_58948_1636# a_59036_1592# 0.28563f
C25810 a_62532_1636# a_62980_1636# 0.01328f
C25811 a_2364_10567# a_2812_10567# 0.0131f
C25812 a_59932_11000# a_59820_10567# 0.02634f
C25813 a_35652_2824# VPWR 0.20815f
C25814 VPWR uio_in[7] 0.0019f
C25815 a_28348_23111# a_28796_23111# 0.01288f
C25816 a_16140_23111# a_16500_23208# 0.08717f
C25817 _459_.CLK a_16052_27912# 0.0054f
C25818 vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN VPWR 0.73788f
C25819 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN ui_in[0] 0.02822f
C25820 a_20060_24679# a_20420_24776# 0.08707f
C25821 _455_.Q a_19860_27912# 0.0011f
C25822 a_1468_21543# a_1916_21543# 0.0131f
C25823 a_2812_9432# VPWR 0.30213f
C25824 a_48508_14136# VPWR 0.29679f
C25825 a_52676_2824# a_52540_1592# 0.00154f
C25826 _442_.ZN a_40668_26247# 0.0064f
C25827 a_32604_18407# a_32516_18504# 0.28563f
C25828 a_39536_26795# a_41116_26247# 0.00516f
C25829 _251_.A1 a_62284_26680# 0.01487f
C25830 _400_.ZN a_44744_26355# 0.04335f
C25831 a_37556_23588# a_37196_23544# 0.0869f
C25832 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN a_64972_26680# 0.00394f
C25833 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_61500_27815# 0.0048f
C25834 a_3172_12232# VPWR 0.20993f
C25835 a_55364_21640# a_55340_19975# 0.00131f
C25836 a_54088_22895# a_54420_21976# 0.00422f
C25837 a_50996_28292# vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.00412f
C25838 a_50524_15704# a_50660_15368# 0.00168f
C25839 a_41700_2824# a_42148_2824# 0.01328f
C25840 a_16052_24776# VPWR 0.20348f
C25841 _475_.Q a_47860_21640# 0.00741f
C25842 a_2364_2727# a_2276_2824# 0.28563f
C25843 _350_.A2 _337_.ZN 1.35685f
C25844 a_3708_19975# a_4068_20072# 0.08717f
C25845 a_45732_15748# VPWR 0.21323f
C25846 a_4852_20072# a_4940_18407# 0.00151f
C25847 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN 0.01287f
C25848 a_5052_18840# a_4964_17316# 0.00151f
C25849 _438_.A2 _300_.ZN 0.03166f
C25850 a_47076_9476# a_46716_9432# 0.08717f
C25851 _311_.A2 _303_.ZN 0.03147f
C25852 _419_.A4 _279_.Z 0.57407f
C25853 a_54468_14180# a_54916_14180# 0.01328f
C25854 _327_.A2 a_40580_20072# 0.00156f
C25855 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_55140_28292# 0.02411f
C25856 _444_.D a_36212_23588# 0.00308f
C25857 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN 0.0024f
C25858 _390_.ZN _402_.A1 0.15046f
C25859 _304_.B a_55228_27815# 0.00447f
C25860 a_3172_12612# a_3260_12568# 0.28563f
C25861 a_53100_18407# a_53124_17316# 0.0016f
C25862 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I VPWR 0.70603f
C25863 _346_.A2 _455_.D 0.33149f
C25864 a_50972_17272# a_50860_16839# 0.02634f
C25865 a_29184_25597# a_30388_25156# 0.00345f
C25866 a_53572_17316# VPWR 0.21311f
C25867 a_24900_23208# a_24876_21976# 0.0016f
C25868 _459_.CLK vgaringosc.workerclkbuff_notouch_.I 0.00994f
C25869 a_65980_1592# VPWR 0.377f
C25870 _384_.ZN _411_.A2 0.4634f
C25871 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[3\].I 1.0811f
C25872 a_33276_1159# a_33636_1256# 0.08717f
C25873 a_4940_24679# a_4964_23588# 0.0016f
C25874 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN 0.09449f
C25875 a_29232_29931# a_30112_30345# 0.00306f
C25876 a_28708_23208# a_28820_22020# 0.02666f
C25877 a_49204_12232# a_49652_12232# 0.01328f
C25878 a_60380_12568# a_60292_11044# 0.00151f
C25879 a_62956_12135# a_63316_12232# 0.08707f
C25880 a_18044_1592# a_18492_1592# 0.01288f
C25881 a_21988_1636# a_22076_1592# 0.28563f
C25882 _324_.C a_63336_29480# 0.0021f
C25883 _229_.I a_62396_27815# 0.00468f
C25884 a_17148_29816# _459_.CLK 0.03553f
C25885 _287_.A1 a_34708_29860# 0.0021f
C25886 a_26556_21543# VPWR 0.32638f
C25887 a_39332_23588# VPWR 0.00683f
C25888 _398_.C _384_.A1 0.35925f
C25889 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN a_55228_28248# 0.00323f
C25890 a_58052_2824# VPWR 0.24545f
C25891 _284_.ZN a_43736_25896# 0.02289f
C25892 a_63652_1636# a_63740_1592# 0.28563f
C25893 a_42372_1636# a_42236_1159# 0.00168f
C25894 a_3172_2824# a_3172_1636# 0.05841f
C25895 clkbuf_1_0__f_clk.I _324_.B 0.01858f
C25896 a_55588_27912# vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.012f
C25897 a_64972_26680# VPWR 0.33187f
C25898 _337_.ZN a_31516_28292# 0.00909f
C25899 a_22212_24776# a_22660_24776# 0.01328f
C25900 a_27452_23111# a_27364_23208# 0.28563f
C25901 a_53436_9432# VPWR 0.31143f
C25902 a_64100_14180# VPWR 0.20967f
C25903 _324_.C a_43936_27165# 0.06035f
C25904 _267_.A2 a_52900_26724# 0.0015f
C25905 a_8996_31048# a_8860_29816# 0.00154f
C25906 a_64884_12232# VPWR 0.23091f
C25907 a_44028_15704# a_44476_15704# 0.01288f
C25908 _388_.B a_48141_29480# 0.02716f
C25909 a_37744_20452# VPWR 0.01415f
C25910 _287_.A1 a_35204_31048# 0.00145f
C25911 _251_.ZN vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN 0.3906f
C25912 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN 0.00301f
C25913 a_67460_18884# a_67436_18407# 0.00172f
C25914 a_63068_18840# a_63068_18407# 0.05841f
C25915 a_34756_24776# VPWR 0.22826f
C25916 _281_.ZN _395_.A3 0.01458f
C25917 a_2724_18884# VPWR 0.20782f
C25918 _459_.D a_30796_24463# 0.22196f
C25919 a_13340_2727# a_13700_2824# 0.08717f
C25920 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_55140_27912# 0.05354f
C25921 a_51868_15704# VPWR 0.32971f
C25922 _370_.B _371_.A2 0.00695f
C25923 a_65308_19975# a_66092_19975# 0.00443f
C25924 _324_.B a_42252_20936# 0.00161f
C25925 _355_.C _352_.ZN 0.13676f
C25926 _230_.I _246_.B2 0.2467f
C25927 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN 0.09948f
C25928 a_62060_23111# clk 0.00239f
C25929 a_48284_17272# a_48196_15748# 0.00151f
C25930 a_1828_20452# a_1468_20408# 0.08717f
C25931 a_3620_20452# a_4068_20452# 0.01328f
C25932 _355_.C a_21540_28292# 0.08159f
C25933 _294_.A2 a_32580_27912# 0.00164f
C25934 a_55228_27815# VPWR 0.29679f
C25935 _336_.Z a_29716_23588# 0.11276f
C25936 a_16028_1592# a_16164_1256# 0.00168f
C25937 a_62532_30736# vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN 0.02628f
C25938 a_47524_12612# a_47612_12568# 0.28563f
C25939 a_51108_12612# a_51556_12612# 0.01328f
C25940 a_63292_2727# a_63740_2727# 0.0131f
C25941 _245_.I1 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN 0.02639f
C25942 _384_.ZN _399_.ZN 0.22943f
C25943 a_65668_9096# a_65668_7908# 0.05841f
C25944 a_44700_1159# a_44612_1256# 0.28563f
C25945 a_63740_12568# a_63652_11044# 0.00151f
C25946 a_66564_7528# a_66564_6340# 0.05841f
C25947 a_32068_20072# a_32516_20072# 0.01328f
C25948 a_20956_1159# VPWR 0.3289f
C25949 a_25348_1636# a_24988_1592# 0.08707f
C25950 a_67460_5960# a_67460_4772# 0.05841f
C25951 a_48384_26724# clkload0.Z 0.93071f
C25952 a_23556_21640# VPWR 0.20614f
C25953 a_49112_29885# a_50032_30345# 0.00306f
C25954 a_37084_26247# a_37532_26247# 0.01222f
C25955 _424_.B1 a_51620_19911# 0.001f
C25956 a_51868_17272# a_52316_17272# 0.01288f
C25957 _325_.ZN a_44300_19001# 0.00125f
C25958 _474_.CLK clk 0.32421f
C25959 a_50188_10567# a_50548_10664# 0.08707f
C25960 a_4828_1159# a_5276_1159# 0.0131f
C25961 a_63852_10567# a_64300_10567# 0.012f
C25962 a_47924_28292# VPWR 0.00683f
C25963 _325_.A2 a_38876_19975# 0.00839f
C25964 a_62420_23208# VPWR 0.20348f
C25965 a_25796_23208# a_26468_23208# 0.00347f
C25966 a_54804_20072# vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN 0.00131f
C25967 _294_.ZN VPWR 1.06995f
C25968 a_19328_28733# uio_out[5] 0.02152f
C25969 _304_.B a_40692_21640# 0.01393f
C25970 a_19076_26344# a_19164_24679# 0.00151f
C25971 a_61524_23208# vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN 0.00129f
C25972 a_66652_6296# VPWR 0.29679f
C25973 a_64412_9432# VPWR 0.30448f
C25974 a_20980_23588# VPWR 0.20622f
C25975 a_32380_21543# a_32828_21543# 0.01288f
C25976 a_1020_2727# VPWR 0.30073f
C25977 a_51084_13703# VPWR 0.31431f
C25978 a_20508_21543# a_20420_21640# 0.28563f
C25979 a_65220_20072# a_66004_20072# 0.00276f
C25980 _459_.CLK a_23920_27555# 0.05733f
C25981 a_40132_26344# VPWR 0.2069f
C25982 _250_.B a_64220_29098# 0.00594f
C25983 _455_.Q a_26556_27815# 0.02518f
C25984 _330_.A1 a_33152_22091# 0.00622f
C25985 a_29351_28293# VPWR 0.0067f
C25986 a_46268_11000# VPWR 0.29679f
C25987 a_14236_29816# a_14236_29383# 0.05841f
C25988 a_51332_15748# a_50972_15704# 0.08707f
C25989 _395_.A1 _384_.A3 0.00526f
C25990 a_64100_2824# a_64548_2824# 0.01328f
C25991 _223_.I _336_.Z 0.00111f
C25992 a_1828_26724# VPWR 0.20348f
C25993 a_14460_30951# a_14596_29860# 0.00154f
C25994 _245_.Z a_60828_26680# 0.00937f
C25995 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_61860_27912# 0.00857f
C25996 _250_.ZN a_60492_28248# 0.0037f
C25997 a_61388_15704# a_62084_15748# 0.01227f
C25998 _345_.A2 a_22992_27555# 0.03995f
C25999 a_31732_20452# a_31708_19975# 0.00172f
C26000 _346_.A2 _454_.D 0.07624f
C26001 a_4852_26344# VPWR 0.22733f
C26002 a_56720_26344# VPWR 0.01026f
C26003 a_45596_30951# vgaringosc.workerclkbuff_notouch_.I 0.00613f
C26004 a_24764_2727# a_24676_2824# 0.28563f
C26005 _451_.Q a_42784_25640# 0.00133f
C26006 _438_.A2 a_38616_24328# 0.41738f
C26007 a_58052_9476# a_57692_9432# 0.08717f
C26008 a_59396_9476# a_59844_9476# 0.01328f
C26009 a_932_23588# a_1380_23588# 0.01328f
C26010 a_1468_28248# VPWR 0.29679f
C26011 a_5636_1256# a_6084_1256# 0.01328f
C26012 _436_.B a_41140_27912# 0.01104f
C26013 _287_.A1 _296_.ZN 0.05144f
C26014 _365_.ZN _359_.B 0.06275f
C26015 a_62844_14136# a_63292_14136# 0.01288f
C26016 a_1828_4772# a_2276_4772# 0.01328f
C26017 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I a_63952_29480# 0.01477f
C26018 a_2724_3204# a_3172_3204# 0.01328f
C26019 a_49112_29885# uio_in[1] 0.00473f
C26020 a_66788_14180# a_66428_14136# 0.08707f
C26021 a_17396_20452# a_17484_20408# 0.28563f
C26022 _336_.Z a_28908_21976# 0.00118f
C26023 _330_.A1 _402_.ZN 0.00315f
C26024 _451_.Q a_40452_18180# 0.00291f
C26025 _416_.A1 a_44028_25156# 0.00277f
C26026 a_54356_23588# a_54444_23544# 0.28563f
C26027 a_22636_29383# VPWR 0.32072f
C26028 a_2724_1636# VPWR 0.20782f
C26029 a_22972_1592# a_23108_1256# 0.00168f
C26030 a_53236_13800# a_53324_12135# 0.00151f
C26031 a_36748_23544# a_36772_23208# 0.00172f
C26032 a_23556_29860# a_23644_29816# 0.28563f
C26033 _459_.CLK a_23196_29816# 0.02822f
C26034 _416_.A1 a_47028_18884# 0.01262f
C26035 _395_.A2 _474_.Q 0.02522f
C26036 a_5500_29816# a_5636_29480# 0.00168f
C26037 _441_.ZN a_40004_23233# 0.02381f
C26038 _433_.ZN a_40656_23588# 0.00449f
C26039 a_43356_1159# VPWR 0.29679f
C26040 a_3172_11044# a_3620_11044# 0.01328f
C26041 a_1380_11044# a_1020_11000# 0.08717f
C26042 a_55676_1159# a_56036_1256# 0.08717f
C26043 a_54692_20452# VPWR 0.20894f
C26044 a_31708_1592# a_32292_1636# 0.01675f
C26045 _251_.ZN vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN 0.00945f
C26046 a_63628_16839# a_64076_16839# 0.0131f
C26047 vgaringosc.workerclkbuff_notouch_.I _480_.Q 0.00155f
C26048 a_41228_27815# a_42236_27815# 0.00323f
C26049 _229_.I a_62756_27912# 0.0025f
C26050 _467_.D a_15244_27815# 0.00241f
C26051 a_61748_23588# a_61612_23111# 0.00168f
C26052 a_61164_10567# a_61076_10664# 0.28563f
C26053 a_3620_18504# a_3620_17316# 0.05841f
C26054 _474_.Q a_46984_23588# 0.05344f
C26055 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I 0.00905f
C26056 a_21876_22020# VPWR 0.21241f
C26057 a_54468_21640# a_54916_21640# 0.01328f
C26058 a_40692_21640# VPWR 0.20948f
C26059 _365_.ZN a_36656_29123# 0.00441f
C26060 a_28460_23544# VPWR 0.31757f
C26061 a_5300_13800# VPWR 0.21406f
C26062 a_4156_18840# a_4604_18840# 0.01222f
C26063 a_31036_21543# a_31396_21640# 0.08707f
C26064 a_23196_2727# VPWR 0.33981f
C26065 a_22996_31048# a_23084_29383# 0.00151f
C26066 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN 0.64692f
C26067 _447_.Q _437_.ZN 0.39381f
C26068 a_18816_29931# uio_out[6] 0.02354f
C26069 a_8100_29860# VPWR 0.21466f
C26070 _275_.ZN VPWR 0.42713f
C26071 _412_.A1 _282_.ZN 0.0215f
C26072 a_59932_11000# VPWR 0.31547f
C26073 a_19636_22020# a_19612_21543# 0.00172f
C26074 a_64412_15704# a_64412_15271# 0.05841f
C26075 a_15692_21976# a_15692_21543# 0.05841f
C26076 a_53996_24679# _384_.A1 0.00102f
C26077 _337_.A3 a_29828_26344# 0.00107f
C26078 a_50524_2727# a_50660_1636# 0.00154f
C26079 a_1916_23111# VPWR 0.297f
C26080 vgaringosc.workerclkbuff_notouch_.I uio_in[0] 0.01502f
C26081 _452_.Q a_42460_20452# 0.00763f
C26082 a_50120_26476# a_50308_26476# 0.00257f
C26083 a_2276_27912# VPWR 0.20634f
C26084 _296_.ZN _293_.A2 0.0377f
C26085 a_62956_23111# a_63316_23208# 0.08717f
C26086 _424_.A2 _421_.A1 0.0077f
C26087 a_35740_2727# a_36100_2824# 0.08717f
C26088 a_53348_18884# a_53436_18840# 0.28563f
C26089 _251_.A1 _258_.I 0.21262f
C26090 _355_.C _345_.A2 0.31666f
C26091 a_1020_6296# a_1020_5863# 0.05841f
C26092 a_1916_4728# a_1916_4295# 0.05841f
C26093 a_65220_4772# a_64860_4728# 0.08717f
C26094 _355_.C a_26746_26344# 0.00505f
C26095 a_2812_3160# a_2812_2727# 0.05841f
C26096 a_66116_3204# a_65756_3160# 0.08717f
C26097 a_22772_20452# a_23220_20452# 0.01328f
C26098 _251_.A1 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN 0.08357f
C26099 a_9084_30951# a_10004_31048# 0.00794f
C26100 a_59036_26247# a_58948_26344# 0.28563f
C26101 a_9635_30644# a_8996_31048# 0.00397f
C26102 a_8860_1592# VPWR 0.33352f
C26103 _319_.A2 _323_.A3 0.01632f
C26104 a_57244_12568# a_57692_12568# 0.01288f
C26105 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN 0.10648f
C26106 a_30778_31048# VPWR 0.01425f
C26107 _337_.A3 a_27328_25227# 0.00232f
C26108 a_66540_19975# a_66564_18884# 0.0016f
C26109 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_61076_23208# 0.08244f
C26110 a_43268_31048# vgaringosc.workerclkbuff_notouch_.I 0.01359f
C26111 _359_.B a_29856_29123# 0.01552f
C26112 _416_.A1 a_51457_29861# 0.05417f
C26113 a_67100_1159# a_67012_1256# 0.28563f
C26114 a_5388_19975# VPWR 0.35526f
C26115 a_65756_1159# VPWR 0.35108f
C26116 a_2724_5960# VPWR 0.20782f
C26117 a_31708_18407# VPWR 0.29679f
C26118 a_45732_11044# a_45372_11000# 0.08707f
C26119 a_39012_1636# a_38652_1592# 0.08707f
C26120 _293_.A2 a_41160_29083# 0.01138f
C26121 a_39684_20452# _325_.A2 0.00227f
C26122 a_43492_27912# _470_.D 0.0014f
C26123 a_28556_29167# _371_.A2 0.00148f
C26124 _398_.C clk 0.99551f
C26125 a_25524_26344# VPWR 0.00698f
C26126 a_57940_10664# a_58388_10664# 0.01328f
C26127 _330_.ZN a_37444_17316# 0.00465f
C26128 a_37408_18504# a_37892_17316# 0.00263f
C26129 a_27004_1159# a_27676_1159# 0.00544f
C26130 a_19972_24776# a_20060_23111# 0.00151f
C26131 _381_.A2 _279_.Z 0.02776f
C26132 a_1468_26680# a_1468_26247# 0.05841f
C26133 a_28012_21976# VPWR 0.31547f
C26134 a_55340_25112# a_55340_24679# 0.05841f
C26135 a_22548_28292# VPWR 0.22567f
C26136 _397_.A1 _384_.A3 0.0984f
C26137 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I 0.66074f
C26138 a_45596_2727# VPWR 0.31143f
C26139 a_66676_13800# VPWR 0.20595f
C26140 a_35504_18955# a_37067_19001# 0.41635f
C26141 a_29604_21640# a_30052_21640# 0.01328f
C26142 a_56932_2824# a_57020_1159# 0.0027f
C26143 a_33140_29860# VPWR 0.00664f
C26144 a_5388_26247# a_5300_26344# 0.28563f
C26145 _441_.A2 a_43126_24119# 0.07236f
C26146 a_31172_15368# a_31620_15368# 0.01328f
C26147 a_14236_29816# VPWR 0.29679f
C26148 _475_.Q a_47483_20569# 0.00215f
C26149 a_67796_16936# a_67908_15748# 0.02666f
C26150 a_46716_10567# VPWR 0.29679f
C26151 a_33052_15271# a_32964_15368# 0.28563f
C26152 a_57468_2727# a_57604_1636# 0.00154f
C26153 a_26580_22020# a_26556_21543# 0.00172f
C26154 a_22636_21976# a_22748_21543# 0.02634f
C26155 _452_.Q a_41664_22020# 0.00241f
C26156 a_32828_23111# VPWR 0.3279f
C26157 a_34620_15271# a_35068_15271# 0.0131f
C26158 _352_.A2 a_28804_27208# 0.00113f
C26159 _304_.A1 _305_.A2 0.00263f
C26160 a_47259_20127# a_47552_19715# 0.49319f
C26161 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN 0.74631f
C26162 a_61748_26724# a_62196_26724# 0.01328f
C26163 a_47164_2727# a_47076_2824# 0.28563f
C26164 a_1828_22020# a_2276_22020# 0.01328f
C26165 a_67012_17316# a_67460_17316# 0.01328f
C26166 a_63428_17316# a_63068_17272# 0.08717f
C26167 a_41056_30669# uo_out[3] 0.05418f
C26168 a_49852_30951# uio_in[1] 0.01264f
C26169 _304_.B _388_.B 0.7353f
C26170 a_43784_19369# VPWR 0.18854f
C26171 a_32848_29123# a_32476_29167# 0.10745f
C26172 a_31920_29480# a_33483_29535# 0.41635f
C26173 _349_.A4 a_26160_27165# 0.00106f
C26174 _480_.Q a_43940_27912# 0.0016f
C26175 a_19276_23544# a_19724_23544# 0.01288f
C26176 a_3260_8999# a_3708_8999# 0.0131f
C26177 _428_.Z a_52852_24372# 0.38933f
C26178 _284_.ZN a_43044_27912# 0.00857f
C26179 a_4156_7431# a_4940_7431# 0.00443f
C26180 a_66764_20408# a_66900_20072# 0.00168f
C26181 a_67548_7864# a_67548_7431# 0.05841f
C26182 a_28036_1256# a_28484_1256# 0.01328f
C26183 a_34404_31048# VPWR 0.01937f
C26184 a_64860_4295# a_65308_4295# 0.0131f
C26185 _325_.ZN a_43932_17800# 0.00997f
C26186 a_3260_13703# a_3620_13800# 0.08717f
C26187 a_39124_16936# a_39324_15271# 0.00119f
C26188 a_7068_2727# a_7516_2727# 0.0131f
C26189 a_28372_20452# a_28460_20408# 0.28563f
C26190 a_57132_13703# a_57580_13703# 0.01288f
C26191 _397_.A2 _384_.ZN 0.38969f
C26192 a_4940_16839# a_5300_16936# 0.08674f
C26193 _411_.A2 a_51576_25896# 0.00991f
C26194 a_22524_1592# VPWR 0.3289f
C26195 a_64548_12612# a_64636_12568# 0.28563f
C26196 a_2364_23544# a_2364_23111# 0.05841f
C26197 a_10540_30951# a_11091_30644# 0.03643f
C26198 _325_.A1 a_43888_19204# 0.03293f
C26199 a_61636_18504# a_62084_18504# 0.01328f
C26200 _287_.A1 _335_.ZN 0.05868f
C26201 _304_.B a_52452_21236# 0.02317f
C26202 a_67772_15271# a_67684_15368# 0.28563f
C26203 a_43380_16936# a_43828_16936# 0.01328f
C26204 a_52092_11000# a_52540_11000# 0.012f
C26205 a_41924_1636# a_42012_1592# 0.28563f
C26206 a_45508_1636# a_45956_1636# 0.01328f
C26207 _304_.A1 a_41440_23208# 0.00306f
C26208 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN a_59260_23111# 0.00244f
C26209 a_3260_26680# a_3708_26680# 0.0131f
C26210 _265_.ZN hold2.Z 0.04616f
C26211 a_24100_29480# VPWR 0.00666f
C26212 _395_.A2 a_50196_22805# 0.01735f
C26213 _336_.A1 a_29348_25940# 0.00152f
C26214 a_31396_2824# a_31260_1592# 0.00154f
C26215 a_5300_21640# a_5388_19975# 0.0027f
C26216 _346_.B a_19948_27815# 0.004f
C26217 a_3708_20408# VPWR 0.33374f
C26218 _452_.CLK a_32740_23208# 0.04879f
C26219 _474_.Q a_51196_21543# 0.01933f
C26220 _388_.B a_47972_31048# 0.00115f
C26221 a_48060_12568# VPWR 0.29679f
C26222 a_67996_2727# VPWR 0.31806f
C26223 a_7876_2824# a_8548_2824# 0.00347f
C26224 a_7964_2727# a_8100_1636# 0.00154f
C26225 _251_.A1 a_62148_29505# 0.00316f
C26226 a_20496_26344# a_21424_25987# 1.16391f
C26227 a_5724_29383# a_6084_29480# 0.08717f
C26228 a_55228_27815# a_55252_26724# 0.0016f
C26229 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I 0.0439f
C26230 a_2364_28248# a_2364_27815# 0.05841f
C26231 a_932_10664# VPWR 0.22176f
C26232 _274_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.88142f
C26233 a_44028_15271# a_44388_15368# 0.08717f
C26234 a_32268_21976# a_32380_21543# 0.02634f
C26235 a_30500_23208# VPWR 0.20622f
C26236 _370_.B _294_.ZN 0.13783f
C26237 a_15604_28292# a_15692_28248# 0.28563f
C26238 _336_.A1 a_28891_25273# 0.1251f
C26239 a_58140_2727# a_58500_2824# 0.08717f
C26240 a_61636_15368# a_62084_15368# 0.01328f
C26241 _388_.B VPWR 1.92721f
C26242 a_66116_15748# VPWR 0.23915f
C26243 _328_.A2 _450_.D 0.11859f
C26244 a_61860_26344# a_61836_25515# 0.03254f
C26245 a_53908_18504# a_54356_18504# 0.01328f
C26246 a_14820_31048# VPWR 0.21092f
C26247 a_17932_25112# a_18380_25112# 0.01288f
C26248 a_21876_25156# a_21964_25112# 0.28563f
C26249 a_27028_23588# a_27116_23544# 0.28563f
C26250 a_4516_7908# VPWR 0.20862f
C26251 a_10340_1256# VPWR 0.20722f
C26252 _448_.Q a_38131_22804# 0.0025f
C26253 a_1916_4728# VPWR 0.297f
C26254 _452_.CLK _316_.A3 0.00232f
C26255 a_31708_18840# a_31708_18407# 0.05841f
C26256 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.00267f
C26257 a_1020_29383# VPWR 0.30073f
C26258 a_54220_13703# a_54132_13800# 0.28563f
C26259 a_33164_20408# _319_.ZN 0.00144f
C26260 _370_.B a_29351_28293# 0.02873f
C26261 a_50324_16936# a_50300_15271# 0.00134f
C26262 a_27004_30951# _371_.ZN 0.00207f
C26263 a_27668_31048# a_28124_30600# 0.02301f
C26264 a_54804_25156# a_54892_25112# 0.28563f
C26265 a_41004_16839# a_40916_16936# 0.28563f
C26266 a_40692_27912# a_40092_27209# 0.01033f
C26267 _311_.A2 a_37644_23544# 0.00619f
C26268 _251_.A1 a_62308_26344# 0.05744f
C26269 _327_.A2 a_43888_19204# 0.00728f
C26270 a_932_16936# VPWR 0.22176f
C26271 a_36324_1636# VPWR 0.2085f
C26272 a_4156_12135# a_4940_12135# 0.00443f
C26273 a_1020_1592# a_1468_1592# 0.01288f
C26274 a_4964_1636# a_5052_1592# 0.28563f
C26275 _460_.Q a_34084_28776# 0.25428f
C26276 _231_.ZN _251_.ZN 0.16585f
C26277 a_45416_29885# _393_.ZN 0.25115f
C26278 a_45904_30180# a_45800_30345# 0.10745f
C26279 a_52452_21236# VPWR 0.82545f
C26280 a_3172_17316# a_3260_17272# 0.28563f
C26281 _384_.ZN a_48308_23588# 0.02651f
C26282 a_61972_12232# a_62060_10567# 0.00151f
C26283 _352_.A2 a_25936_25597# 0.03653f
C26284 a_59396_11044# a_59036_11000# 0.08707f
C26285 a_17148_1592# a_17148_1159# 0.05841f
C26286 a_21092_1636# a_20956_1159# 0.00168f
C26287 a_54444_25112# VPWR 0.29679f
C26288 a_58388_17316# a_58476_17272# 0.28563f
C26289 _419_.A4 a_48888_19243# 0.0014f
C26290 _251_.A1 _255_.ZN 0.11652f
C26291 a_58140_26680# vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I 0.00115f
C26292 a_49404_1159# a_49852_1159# 0.0131f
C26293 a_43452_18191# a_43796_18559# 0.00275f
C26294 a_38340_2824# a_38204_1592# 0.00154f
C26295 a_15156_27912# a_15156_26724# 0.05841f
C26296 a_4068_25156# VPWR 0.2157f
C26297 a_67012_18884# a_67460_18884# 0.01328f
C26298 a_62980_18884# a_63068_18840# 0.28563f
C26299 a_2812_27815# a_2724_27912# 0.28563f
C26300 a_23756_20408# VPWR 0.31143f
C26301 a_61836_25515# a_62404_25156# 0.03324f
C26302 _229_.I ui_in[2] 0.00218f
C26303 _416_.A1 a_45696_20072# 0.0447f
C26304 a_37084_25112# _444_.D 0.01584f
C26305 a_4516_15748# a_4156_15704# 0.08674f
C26306 a_1916_15704# a_2364_15704# 0.0131f
C26307 a_61860_12612# VPWR 0.20595f
C26308 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I a_65756_26247# 0.00442f
C26309 a_36188_15704# a_36324_15368# 0.00168f
C26310 a_16700_29383# _467_.D 0.01771f
C26311 a_53572_15368# a_54020_15368# 0.01328f
C26312 a_17148_29383# a_17060_29480# 0.28563f
C26313 _324_.C _243_.ZN 0.00588f
C26314 a_62420_10664# VPWR 0.20641f
C26315 a_53996_24679# clk 0.01873f
C26316 a_932_9096# a_1380_9096# 0.01328f
C26317 a_30924_21976# a_30948_21640# 0.00172f
C26318 a_65756_5863# a_66116_5960# 0.08717f
C26319 _371_.A1 a_28596_26725# 0.00417f
C26320 a_64860_7431# a_65220_7528# 0.08717f
C26321 a_55452_15271# a_55364_15368# 0.28563f
C26322 _304_.B a_40580_20072# 0.00157f
C26323 a_66652_4295# a_67012_4392# 0.08717f
C26324 a_22300_21543# a_22324_20452# 0.0016f
C26325 a_36284_29167# VPWR 0.39596f
C26326 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN a_65644_23544# 0.0016f
C26327 a_35876_15368# VPWR 0.20348f
C26328 a_56796_15271# vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN 0.00402f
C26329 a_20172_21976# a_20620_21976# 0.01288f
C26330 a_57468_16839# VPWR 0.34384f
C26331 _474_.CLK a_49652_29480# 0.00457f
C26332 a_39324_15271# VPWR 0.32938f
C26333 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN 0.17736f
C26334 a_27564_23544# a_27476_22020# 0.00151f
C26335 a_3172_14180# a_3260_14136# 0.28563f
C26336 a_38316_16839# a_38764_16839# 0.01288f
C26337 _362_.B VPWR 2.35896f
C26338 a_63516_17272# VPWR 0.31389f
C26339 a_32740_1256# VPWR 0.20348f
C26340 a_50436_1256# a_50884_1256# 0.01328f
C26341 a_67548_7431# VPWR 0.32135f
C26342 a_31820_23544# a_32268_23544# 0.012f
C26343 _260_.ZN a_43192_22504# 0.00179f
C26344 a_50996_13800# a_51444_13800# 0.01328f
C26345 _384_.ZN _330_.A1 0.02452f
C26346 a_37067_19001# a_37408_18504# 0.00242f
C26347 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN 0.00288f
C26348 a_64972_13703# a_65332_13800# 0.08717f
C26349 a_29468_2727# a_29916_2727# 0.0131f
C26350 _234_.ZN _436_.B 0.49364f
C26351 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN 0.74383f
C26352 a_16252_30951# VPWR 0.32936f
C26353 a_51756_16839# a_52116_16936# 0.08717f
C26354 a_55028_10664# a_55140_9476# 0.02666f
C26355 a_66452_18504# VPWR 0.21172f
C26356 _268_.A2 a_52640_29860# 0.00544f
C26357 a_10876_1159# a_10788_1256# 0.28563f
C26358 a_51196_1592# a_51332_1256# 0.00168f
C26359 a_43828_29860# a_43916_29816# 0.28563f
C26360 a_47860_16936# VPWR 0.20703f
C26361 _388_.B _383_.ZN 0.17902f
C26362 a_42460_1592# VPWR 0.35102f
C26363 a_58476_20408# a_58388_18884# 0.00251f
C26364 _452_.D a_42148_15748# 0.0019f
C26365 a_1468_12135# a_1380_12232# 0.28563f
C26366 vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I 0.64261f
C26367 a_26720_30301# _349_.A4 0.20675f
C26368 _390_.ZN _407_.A1 0.04748f
C26369 a_26427_29977# a_26672_30345# 0.00232f
C26370 a_6396_29816# a_6844_29816# 0.01288f
C26371 a_36548_17316# a_36996_17316# 0.01328f
C26372 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I 0.0025f
C26373 a_32964_17316# a_33052_17272# 0.28563f
C26374 a_48644_15368# a_48508_14136# 0.00154f
C26375 a_23084_30951# uio_out[4] 0.00623f
C26376 a_52452_15368# a_52452_14180# 0.05841f
C26377 _459_.CLK _437_.A1 0.00212f
C26378 _436_.B a_41476_26344# 0.00725f
C26379 a_62756_11044# a_62396_11000# 0.08707f
C26380 a_65892_11044# a_66340_11044# 0.01328f
C26381 a_63952_29480# vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN 0.00349f
C26382 a_12804_2824# VPWR 0.20348f
C26383 a_51644_1592# a_52092_1592# 0.01288f
C26384 _363_.Z a_32240_31048# 0.10862f
C26385 a_32628_26725# VPWR 0.59766f
C26386 a_17036_23111# a_17484_23111# 0.0131f
C26387 _459_.CLK a_17844_26344# 0.00641f
C26388 _455_.Q a_21052_26031# 0.00278f
C26389 a_4604_6296# a_4516_4772# 0.0027f
C26390 a_66340_15368# VPWR 0.21266f
C26391 a_22548_25156# VPWR 0.22672f
C26392 a_17396_27912# a_17844_27912# 0.01328f
C26393 a_34308_15748# a_33948_15704# 0.08707f
C26394 a_48508_12135# VPWR 0.31817f
C26395 a_30276_2824# a_30724_2824# 0.01328f
C26396 a_44795_29535# a_45088_29123# 0.49319f
C26397 _268_.A2 _274_.A3 0.13648f
C26398 _433_.ZN _448_.Q 0.03594f
C26399 a_1916_24679# VPWR 0.297f
C26400 a_44924_15704# a_44924_15271# 0.05841f
C26401 a_55588_28292# a_56036_28292# 0.01328f
C26402 a_59708_23111# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I 0.00455f
C26403 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_61164_23111# 0.00933f
C26404 a_40580_20072# VPWR 0.20765f
C26405 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN 0.06974f
C26406 a_20868_21640# a_20844_20408# 0.0016f
C26407 _452_.CLK a_45260_16839# 0.00207f
C26408 a_31620_15748# VPWR 0.20348f
C26409 _293_.A2 a_40038_28720# 0.02702f
C26410 _324_.C _258_.ZN 0.01122f
C26411 _384_.ZN a_48988_26369# 0.00188f
C26412 a_2276_9476# a_2724_9476# 0.01328f
C26413 _319_.A3 a_35716_20072# 0.02085f
C26414 a_27476_22020# a_27116_21976# 0.08707f
C26415 _459_.CLK _340_.ZN 0.63517f
C26416 a_67908_22020# a_67772_21543# 0.00168f
C26417 a_47524_14180# a_47612_14136# 0.28563f
C26418 a_51108_14180# a_51556_14180# 0.01328f
C26419 _424_.B1 _399_.A1 0.00986f
C26420 a_49204_16936# a_49092_15748# 0.02666f
C26421 a_43020_16839# VPWR 0.33033f
C26422 _462_.D _288_.ZN 0.10692f
C26423 a_55140_1256# VPWR 0.20348f
C26424 a_65532_14136# a_65444_12612# 0.00151f
C26425 a_45732_13800# a_45732_12612# 0.05841f
C26426 _416_.A3 a_47636_18884# 0.04883f
C26427 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I 0.00107f
C26428 a_58911_30644# VPWR 0.31359f
C26429 _459_.CLK a_32180_23588# 0.00176f
C26430 a_33500_17272# VPWR 0.30042f
C26431 a_62420_10664# a_62308_9476# 0.02666f
C26432 a_60628_10664# a_60604_9432# 0.0016f
C26433 a_29692_23111# a_29716_22020# 0.0016f
C26434 _416_.A2 a_47552_19715# 0.05241f
C26435 a_64412_29816# a_65072_29860# 0.01375f
C26436 a_31844_26344# a_32292_26344# 0.01328f
C26437 a_56260_1636# VPWR 0.2085f
C26438 a_21852_1159# a_22212_1256# 0.08717f
C26439 a_51980_12135# a_52340_12232# 0.08707f
C26440 a_14684_1592# a_15132_1592# 0.01288f
C26441 _404_.A1 a_48384_26724# 0.0011f
C26442 a_24876_23544# a_24900_23208# 0.00172f
C26443 _402_.A1 a_45232_25987# 0.00386f
C26444 a_15044_29480# a_15492_29480# 0.01328f
C26445 a_65868_12135# a_66316_12135# 0.0131f
C26446 a_13700_29860# a_13340_29816# 0.08707f
C26447 a_38616_24328# a_39004_24463# 0.00334f
C26448 a_4940_26247# a_4964_25156# 0.0016f
C26449 a_35204_2824# VPWR 0.23994f
C26450 a_58911_30644# a_59332_29816# 0.00234f
C26451 a_58948_1636# a_58588_1592# 0.08707f
C26452 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I 0.01311f
C26453 vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN 0.03158f
C26454 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN 0.00128f
C26455 a_16140_23111# a_16052_23208# 0.28563f
C26456 a_1828_24776# a_2276_24776# 0.01328f
C26457 a_20060_24679# a_19972_24776# 0.28563f
C26458 a_2364_9432# VPWR 0.30029f
C26459 a_65668_9096# a_66116_9096# 0.01328f
C26460 a_66564_7528# a_67012_7528# 0.01328f
C26461 a_48060_14136# VPWR 0.29679f
C26462 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN 0.68282f
C26463 _251_.A1 a_61836_26680# 0.00502f
C26464 a_24304_26795# _351_.ZN 0.24887f
C26465 a_1380_18504# a_1828_18504# 0.01328f
C26466 a_32156_18407# a_32516_18504# 0.08717f
C26467 _442_.ZN a_40220_26247# 0.01697f
C26468 a_37108_23588# a_37196_23544# 0.28563f
C26469 _230_.I a_60492_28248# 0.01316f
C26470 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN a_63180_26680# 0.00151f
C26471 a_17956_29860# uio_out[7] 0.01285f
C26472 a_2724_12232# VPWR 0.20782f
C26473 a_40804_15748# a_41252_15748# 0.01328f
C26474 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_61052_27815# 0.00241f
C26475 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I a_62172_19975# 0.00224f
C26476 _424_.A2 _305_.A2 0.02093f
C26477 vgaringosc.workerclkbuff_notouch_.I _274_.ZN 0.47519f
C26478 a_15604_24776# VPWR 0.20348f
C26479 a_1916_2727# a_2276_2824# 0.08717f
C26480 a_45284_15748# VPWR 0.20703f
C26481 a_3708_19975# a_3620_20072# 0.28563f
C26482 _223_.I _287_.A1 0.01801f
C26483 _402_.A1 a_49740_29383# 0.01605f
C26484 a_46628_9476# a_46716_9432# 0.28563f
C26485 _337_.A3 a_24304_26795# 0.00726f
C26486 a_31820_21976# a_32268_21976# 0.012f
C26487 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.00943f
C26488 _438_.ZN a_39796_22504# 0.02744f
C26489 _419_.A4 a_47297_25596# 0.06292f
C26490 _438_.A2 a_38852_25156# 0.00202f
C26491 _267_.A2 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I 0.01466f
C26492 _304_.B a_53660_27815# 0.01816f
C26493 _223_.I a_31932_26247# 0.00448f
C26494 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN 0.02447f
C26495 a_51868_2727# a_52316_2727# 0.0131f
C26496 a_3172_12612# a_2812_12568# 0.08717f
C26497 _437_.A1 uo_out[7] 0.09348f
C26498 _346_.A2 a_20844_26680# 0.00155f
C26499 _247_.ZN _247_.B 0.0148f
C26500 a_35232_24029# a_36212_23588# 0.00702f
C26501 a_29232_29931# a_29620_30345# 0.00393f
C26502 a_53124_17316# VPWR 0.20692f
C26503 a_53212_29816# vgaringosc.ro_inv4.inv_array_notouch_\[3\].I 0.00435f
C26504 a_33276_1159# a_33188_1256# 0.28563f
C26505 a_66876_1592# a_67012_1256# 0.00168f
C26506 a_65532_1592# VPWR 0.33691f
C26507 a_62956_12135# a_62868_12232# 0.28563f
C26508 a_21988_1636# a_21628_1592# 0.08707f
C26509 _229_.I a_61948_27815# 0.00718f
C26510 _287_.A1 a_34260_29860# 0.00199f
C26511 a_20379_29977# a_20672_30301# 0.58767f
C26512 _268_.A2 _324_.C 0.03081f
C26513 _379_.A2 _375_.Z 0.35296f
C26514 a_16700_29816# _459_.CLK 0.00923f
C26515 a_25884_21543# VPWR 0.34806f
C26516 a_17396_26344# a_17396_25156# 0.05841f
C26517 a_48644_17316# a_49092_17316# 0.01328f
C26518 a_66876_11000# a_66764_10567# 0.02634f
C26519 a_52876_10567# a_53324_10567# 0.01288f
C26520 a_57380_2824# VPWR 0.21976f
C26521 a_63068_1592# a_63740_1592# 0.00544f
C26522 a_65444_1636# a_65892_1636# 0.01328f
C26523 _261_.ZN _448_.Q 0.47724f
C26524 clkbuf_1_0__f_clk.I a_47860_23208# 0.04077f
C26525 a_55140_27912# vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I 0.00316f
C26526 a_55588_27912# a_56036_27912# 0.01328f
C26527 _411_.A2 clkload0.Z 0.03389f
C26528 a_14708_23208# a_15156_23208# 0.01328f
C26529 a_27004_23111# a_27364_23208# 0.08707f
C26530 a_63180_26680# VPWR 0.32012f
C26531 a_27172_24328# a_27552_24397# 0.00372f
C26532 _337_.ZN a_31068_28292# 0.00653f
C26533 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN VPWR 0.74675f
C26534 a_52988_9432# VPWR 0.31605f
C26535 _281_.A1 a_54420_21976# 0.00576f
C26536 a_21404_21543# a_21852_21543# 0.01288f
C26537 a_63652_14180# VPWR 0.20952f
C26538 a_23108_2824# a_23196_1159# 0.0027f
C26539 _324_.C a_43008_26795# 0.05838f
C26540 _476_.Q a_53572_21640# 0.00208f
C26541 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN clk 0.00467f
C26542 a_64212_12232# VPWR 0.21343f
C26543 _399_.A1 _218_.ZN 0.2178f
C26544 a_36188_2727# a_36324_1636# 0.00154f
C26545 a_52676_2824# a_53124_2824# 0.01328f
C26546 a_36008_20569# VPWR 0.00204f
C26547 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN a_57020_23111# 0.00124f
C26548 _473_.Q a_49828_22020# 0.00494f
C26549 _251_.ZN a_58364_25112# 0.00236f
C26550 a_6723_30644# a_6756_29860# 0.02559f
C26551 _229_.I a_61297_30300# 0.56373f
C26552 a_34308_24776# VPWR 0.23398f
C26553 _397_.A4 _397_.Z 0.01076f
C26554 a_2276_18884# VPWR 0.20634f
C26555 _459_.D a_31168_24419# 0.00761f
C26556 _379_.Z a_17932_27815# 0.00154f
C26557 a_13340_2727# a_13252_2824# 0.28563f
C26558 a_58588_26247# clk 0.00109f
C26559 a_51420_15704# VPWR 0.32971f
C26560 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I a_53572_27912# 0.0054f
C26561 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I 0.00888f
C26562 _416_.A1 _260_.A1 0.27792f
C26563 _355_.C a_24316_26247# 0.0241f
C26564 a_51868_9432# a_52316_9432# 0.0131f
C26565 _301_.A1 _319_.A3 0.00742f
C26566 _416_.A1 a_47047_21640# 0.00406f
C26567 a_61612_23111# clk 0.00209f
C26568 a_58924_14136# a_59372_14136# 0.01255f
C26569 a_1380_20452# a_1468_20408# 0.28563f
C26570 _447_.Q a_39669_21236# 0.00497f
C26571 _355_.C a_19328_28733# 0.11499f
C26572 a_53660_27815# VPWR 0.33665f
C26573 _294_.A2 a_32132_27912# 0.00234f
C26574 _336_.Z a_28820_24072# 0.2848f
C26575 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I VPWR 0.88657f
C26576 a_47524_12612# a_47164_12568# 0.08707f
C26577 _231_.ZN vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I 0.03167f
C26578 _397_.A1 _402_.B 0.00117f
C26579 a_20508_1159# VPWR 0.3289f
C26580 a_44252_1159# a_44612_1256# 0.08717f
C26581 _234_.ZN a_40464_27165# 0.00337f
C26582 a_24900_1636# a_24988_1592# 0.28563f
C26583 a_28484_1636# a_28932_1636# 0.01328f
C26584 a_44476_27815# _403_.ZN 0.00617f
C26585 a_59732_12232# a_60180_12232# 0.01328f
C26586 a_23108_21640# VPWR 0.20614f
C26587 _435_.A3 a_40468_25157# 0.03106f
C26588 _452_.CLK hold2.Z 0.00826f
C26589 a_50188_10567# a_50100_10664# 0.28563f
C26590 a_63740_11000# a_63764_10664# 0.00172f
C26591 _402_.A1 a_48376_27508# 0.00113f
C26592 _325_.A2 a_37384_19624# 0.22881f
C26593 a_47700_28292# VPWR 0.01391f
C26594 _285_.Z uo_out[1] 0.97434f
C26595 a_54804_20072# a_54892_18407# 0.00151f
C26596 _451_.Q a_41488_24072# 0.00112f
C26597 a_61972_23208# VPWR 0.20567f
C26598 a_19035_28409# uio_out[5] 0.00338f
C26599 a_30240_24776# a_30628_24463# 0.00393f
C26600 _460_.Q a_33776_29123# 0.00742f
C26601 _304_.B a_40244_21640# 0.01693f
C26602 a_66204_6296# VPWR 0.31657f
C26603 a_20532_23588# VPWR 0.20622f
C26604 a_20060_21543# a_20420_21640# 0.08707f
C26605 a_67460_9476# VPWR 0.21296f
C26606 a_67996_3160# VPWR 0.31806f
C26607 a_50636_13703# VPWR 0.33817f
C26608 _459_.CLK a_23627_27967# 0.05371f
C26609 _412_.B2 _417_.A2 0.04033f
C26610 _455_.Q a_25884_27815# 0.01783f
C26611 a_39684_26344# VPWR 0.20587f
C26612 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN a_61276_19975# 0.00636f
C26613 _459_.CLK _355_.B 0.02336f
C26614 a_46940_15704# a_47388_15704# 0.01288f
C26615 a_45820_11000# VPWR 0.29679f
C26616 a_42784_22504# VPWR 0.00171f
C26617 a_50884_15748# a_50972_15704# 0.28563f
C26618 a_1380_26724# VPWR 0.20348f
C26619 _325_.A2 a_43796_18559# 0.00108f
C26620 _346_.A2 a_22064_27912# 0.01217f
C26621 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_61412_27912# 0.0036f
C26622 _245_.Z a_59620_27208# 0.46003f
C26623 a_45148_30951# vgaringosc.workerclkbuff_notouch_.I 0.00613f
C26624 a_4068_26344# VPWR 0.22146f
C26625 a_56368_26344# VPWR 0.00645f
C26626 a_24316_2727# a_24676_2824# 0.08717f
C26627 _324_.B a_42168_22504# 1.98935f
C26628 _451_.Q a_42376_25640# 0.00167f
C26629 _460_.Q a_36100_26724# 0.00683f
C26630 a_1020_28248# VPWR 0.30073f
C26631 a_57604_9476# a_57692_9432# 0.28563f
C26632 _436_.B a_40692_27912# 0.0319f
C26633 a_66340_14180# a_66428_14136# 0.28563f
C26634 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I 0.001f
C26635 a_15244_20408# a_15692_20408# 0.0131f
C26636 a_17396_20452# a_17036_20408# 0.08717f
C26637 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I 0.01734f
C26638 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN a_61076_23208# 0.00196f
C26639 a_54420_21976# a_54816_22505# 0.00232f
C26640 a_22188_29383# VPWR 0.32626f
C26641 a_2276_1636# VPWR 0.20634f
C26642 a_54020_12612# a_54468_12612# 0.01328f
C26643 _303_.ZN a_42392_19243# 0.00534f
C26644 a_23556_29860# a_23196_29816# 0.08674f
C26645 a_55676_1159# a_55588_1256# 0.28563f
C26646 a_42908_1159# VPWR 0.31729f
C26647 _416_.A1 _470_.Q 0.00807f
C26648 a_932_11044# a_1020_11000# 0.28563f
C26649 a_54244_20452# VPWR 0.20878f
C26650 vgaringosc.workerclkbuff_notouch_.I a_43232_29480# 0.01363f
C26651 _252_.B a_59620_27208# 0.23777f
C26652 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I a_58388_13800# 0.00198f
C26653 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN a_58500_21640# 0.07112f
C26654 _229_.I a_62308_27912# 0.00478f
C26655 a_46628_10664# a_47076_10664# 0.01328f
C26656 a_56260_1636# a_56124_1159# 0.00168f
C26657 a_15580_1159# a_16252_1159# 0.00544f
C26658 a_60716_10567# a_61076_10664# 0.08707f
C26659 a_17060_2824# a_17060_1636# 0.05841f
C26660 a_54804_23588# a_55252_23588# 0.01328f
C26661 a_21428_22020# VPWR 0.20622f
C26662 _287_.A1 a_37584_29123# 0.00377f
C26663 _365_.ZN a_35728_29480# 0.05954f
C26664 a_40244_21640# VPWR 0.13651f
C26665 a_28012_23544# VPWR 0.31547f
C26666 uio_out[5] uio_out[7] 0.03027f
C26667 a_31036_21543# a_30948_21640# 0.28563f
C26668 a_18628_21640# a_19076_21640# 0.01328f
C26669 a_22748_2727# VPWR 0.31143f
C26670 a_4852_13800# VPWR 0.22733f
C26671 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN VPWR 0.99049f
C26672 a_62172_15271# a_62620_15271# 0.0131f
C26673 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN a_58476_20408# 0.05535f
C26674 a_7652_29860# VPWR 0.20641f
C26675 a_48708_29816# VPWR 0.36686f
C26676 a_54108_21543# a_54244_20452# 0.00154f
C26677 a_59484_11000# VPWR 0.31547f
C26678 a_41564_26247# a_41476_26344# 0.28563f
C26679 a_67460_15748# a_67324_15271# 0.00168f
C26680 a_1468_23111# VPWR 0.29679f
C26681 _267_.A1 a_56124_28248# 0.00155f
C26682 a_65756_15704# a_66204_15704# 0.01255f
C26683 _296_.ZN a_37968_31048# 0.00253f
C26684 a_1828_27912# VPWR 0.20348f
C26685 _441_.B a_38576_22504# 0.00346f
C26686 a_35740_2727# a_35652_2824# 0.28563f
C26687 a_62956_23111# a_62868_23208# 0.28563f
C26688 _362_.B _360_.ZN 0.00224f
C26689 _371_.A3 _355_.B 0.0097f
C26690 a_49896_18909# a_51308_19369# 0.00393f
C26691 _251_.ZN clk 0.0041f
C26692 a_62844_9432# a_63292_9432# 0.0131f
C26693 _448_.Q _327_.Z 0.00827f
C26694 a_16052_23588# a_16500_23588# 0.01328f
C26695 a_64772_7908# a_65220_7908# 0.01328f
C26696 a_16612_1256# a_17060_1256# 0.01328f
C26697 a_65668_6340# a_66116_6340# 0.01328f
C26698 _334_.A1 _452_.CLK 0.00826f
C26699 a_67460_3204# a_67908_3204# 0.01328f
C26700 a_65668_3204# a_65756_3160# 0.28563f
C26701 a_4964_3204# a_4828_2727# 0.00168f
C26702 a_45820_13703# a_46268_13703# 0.0131f
C26703 a_66564_4772# a_67012_4772# 0.01328f
C26704 a_64772_4772# a_64860_4728# 0.28563f
C26705 _251_.A1 a_62396_26247# 0.04763f
C26706 a_7068_29383# a_7516_29383# 0.0131f
C26707 a_9084_30951# a_8996_31048# 0.28563f
C26708 a_58588_26247# a_58948_26344# 0.08674f
C26709 _421_.A1 clkbuf_1_0__f_clk.I 0.39614f
C26710 _275_.ZN _407_.ZN 0.0021f
C26711 _384_.ZN _393_.A1 0.44819f
C26712 _304_.B vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN 0.05767f
C26713 a_15940_1636# VPWR 0.21466f
C26714 a_63764_13800# a_63852_12135# 0.00151f
C26715 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I 0.04598f
C26716 _459_.CLK a_25643_25273# 0.00106f
C26717 _416_.A1 _260_.A2 0.11271f
C26718 _359_.B a_29563_29535# 0.01391f
C26719 a_42820_31048# vgaringosc.workerclkbuff_notouch_.I 0.00697f
C26720 _230_.I vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 0.00442f
C26721 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_59620_23208# 0.00236f
C26722 _330_.ZN a_38764_16839# 0.0059f
C26723 a_48868_11044# a_49316_11044# 0.01328f
C26724 a_45284_11044# a_45372_11000# 0.28563f
C26725 a_4940_19975# VPWR 0.31945f
C26726 a_65084_1159# VPWR 0.33093f
C26727 a_2276_5960# VPWR 0.20634f
C26728 a_66652_1159# a_67012_1256# 0.0869f
C26729 a_31260_18407# VPWR 0.29679f
C26730 a_6756_1636# a_6620_1159# 0.00168f
C26731 a_2812_1592# a_2812_1159# 0.05841f
C26732 a_34620_1592# a_35068_1592# 0.01288f
C26733 a_38564_1636# a_38652_1592# 0.28563f
C26734 a_32068_16936# a_32516_16936# 0.01328f
C26735 a_36636_25112# a_37084_25112# 0.01255f
C26736 a_32628_26725# _360_.ZN 0.00441f
C26737 _304_.B _402_.A1 1.47197f
C26738 _293_.A2 a_37584_29123# 0.01161f
C26739 a_38676_20452# _325_.A2 0.00242f
C26740 _330_.A1 a_36612_20072# 0.01262f
C26741 a_25300_26344# VPWR 0.01379f
C26742 a_28928_29123# _371_.A2 0.00144f
C26743 _330_.ZN a_36996_17316# 0.00224f
C26744 a_63616_31128# vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I 0.01211f
C26745 _381_.A2 a_47297_25596# 0.18651f
C26746 a_27564_21976# VPWR 0.32115f
C26747 _397_.A1 a_52900_26724# 0.06118f
C26748 a_21628_28248# VPWR 0.3424f
C26749 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I a_62508_21976# 0.0046f
C26750 a_43356_30951# a_43804_30951# 0.0131f
C26751 _433_.ZN a_41664_22020# 0.00621f
C26752 a_35008_22461# a_34160_20523# 0.00114f
C26753 a_45148_2727# VPWR 0.31143f
C26754 _316_.ZN a_34716_20937# 0.00206f
C26755 a_66228_13800# VPWR 0.22482f
C26756 a_35504_18955# a_37360_19325# 0.02307f
C26757 a_36432_19325# a_36060_19369# 0.10745f
C26758 a_32916_29860# VPWR 0.01378f
C26759 a_4940_26247# a_5300_26344# 0.08674f
C26760 a_19164_26247# a_19612_26247# 0.012f
C26761 _441_.A2 a_42796_23981# 0.0137f
C26762 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN 0.00916f
C26763 _475_.Q a_47776_20893# 0.22338f
C26764 a_13788_29816# VPWR 0.29679f
C26765 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN 0.27893f
C26766 a_64436_16936# a_64412_15704# 0.0016f
C26767 a_46268_10567# VPWR 0.29679f
C26768 a_32604_15271# a_32964_15368# 0.08717f
C26769 _447_.Q _316_.A3 0.06801f
C26770 a_32380_23111# VPWR 0.3158f
C26771 _350_.A1 _459_.CLK 0.04278f
C26772 a_62284_23544# a_62420_23208# 0.00168f
C26773 _452_.Q a_41460_22020# 0.0218f
C26774 _407_.A1 a_51317_27508# 0.00936f
C26775 _474_.D a_50280_19369# 0.01093f
C26776 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN 0.0205f
C26777 _324_.B _473_.Q 0.37606f
C26778 _352_.A2 a_28124_26680# 0.04606f
C26779 a_932_28292# a_1380_28292# 0.01328f
C26780 _246_.B2 _244_.Z 0.03437f
C26781 a_46716_2727# a_47076_2824# 0.08717f
C26782 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN 0.04138f
C26783 a_62980_17316# a_63068_17272# 0.28563f
C26784 a_49404_30951# uio_in[1] 0.00503f
C26785 a_31920_29480# a_32476_29167# 0.8399f
C26786 a_29563_29535# a_29808_29167# 0.00232f
C26787 a_43888_19204# VPWR 0.39816f
C26788 a_41056_30669# _388_.B 0.47908f
C26789 _459_.Q a_30932_26020# 0.00372f
C26790 a_1380_16936# a_1380_15748# 0.05841f
C26791 _349_.A4 a_24860_27209# 0.00106f
C26792 a_53300_23047# a_53648_23263# 0.00277f
C26793 a_66988_18407# a_67436_18407# 0.01255f
C26794 _395_.A3 _475_.Q 0.0551f
C26795 _428_.Z a_51332_24372# 0.03877f
C26796 a_38576_22504# _300_.A2 0.23809f
C26797 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN a_64860_26247# 0.00383f
C26798 a_66204_9432# a_66204_8999# 0.05841f
C26799 vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN 0.00791f
C26800 _284_.ZN a_42596_27912# 0.0036f
C26801 a_14708_25156# a_15156_25156# 0.01328f
C26802 a_1020_5863# a_932_5960# 0.28563f
C26803 a_33956_31048# VPWR 0.01438f
C26804 _474_.CLK _284_.A2 0.78572f
C26805 a_3260_13703# a_3172_13800# 0.28563f
C26806 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I 0.17423f
C26807 a_26220_20408# a_26668_20408# 0.0131f
C26808 _352_.A2 _369_.ZN 0.31933f
C26809 a_28372_20452# a_28012_20408# 0.08717f
C26810 _258_.I _255_.I 0.10605f
C26811 a_60285_30600# a_60276_29032# 0.00145f
C26812 a_64324_18504# a_64324_17316# 0.05841f
C26813 _411_.A2 a_50120_26476# 0.40032f
C26814 a_4940_16839# a_4852_16936# 0.28563f
C26815 _397_.A4 _284_.B 0.02667f
C26816 _324_.B a_42996_18840# 0.00126f
C26817 _363_.Z a_35204_26344# 0.00145f
C26818 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN VPWR 1.19537f
C26819 a_24864_29931# _342_.ZN 0.25068f
C26820 a_22076_1592# VPWR 0.3289f
C26821 a_36860_1592# a_36996_1256# 0.00168f
C26822 a_64548_12612# a_64188_12568# 0.08707f
C26823 _325_.A1 a_43400_18909# 0.11531f
C26824 _417_.A2 a_49448_20936# 0.00183f
C26825 a_50996_12232# a_51084_10567# 0.00151f
C26826 a_67324_15271# a_67684_15368# 0.08663f
C26827 _359_.B _304_.B 0.0364f
C26828 _304_.A1 a_41216_23208# 0.00161f
C26829 a_41924_1636# a_41564_1592# 0.08707f
C26830 _402_.A1 VPWR 3.52155f
C26831 _397_.A2 clkload0.Z 0.02811f
C26832 _304_.B a_53996_25112# 0.00191f
C26833 _304_.A1 _325_.A1 0.46731f
C26834 _336_.A1 a_29164_25940# 0.00401f
C26835 a_22996_29480# VPWR 0.20924f
C26836 a_37980_1159# a_38428_1159# 0.0131f
C26837 _346_.B a_19500_27815# 0.00202f
C26838 _371_.ZN a_28388_29167# 0.0014f
C26839 _340_.A2 _340_.ZN 0.41461f
C26840 a_3260_20408# VPWR 0.30487f
C26841 _452_.CLK a_32292_23208# 0.00857f
C26842 a_67908_2824# a_67996_1159# 0.0027f
C26843 a_62644_16936# a_63092_16936# 0.01328f
C26844 a_67548_2727# VPWR 0.29679f
C26845 a_47612_12568# VPWR 0.29679f
C26846 _267_.ZN a_52764_27815# 0.00146f
C26847 _452_.CLK _448_.Q 0.11388f
C26848 _243_.A1 VPWR 0.64045f
C26849 _251_.A1 a_60916_29612# 0.00161f
C26850 a_5724_29383# a_5636_29480# 0.28563f
C26851 a_42148_15368# a_42596_15368# 0.01328f
C26852 a_68108_10567# VPWR 0.35526f
C26853 a_44028_15271# a_43940_15368# 0.28563f
C26854 hold1.Z _305_.A2 0.05447f
C26855 a_30052_23208# VPWR 0.20862f
C26856 _390_.ZN a_52764_27815# 0.00189f
C26857 a_45372_15271# a_46044_15271# 0.00544f
C26858 a_55340_19975# vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN 0.00891f
C26859 _324_.C _241_.I0 0.01541f
C26860 a_15604_28292# a_15244_28248# 0.0869f
C26861 _336_.A1 a_29184_25597# 0.26108f
C26862 a_16948_22020# a_17396_22020# 0.01328f
C26863 _355_.C _352_.A2 1.25879f
C26864 a_65668_15748# VPWR 0.21723f
C26865 a_58140_2727# a_58052_2824# 0.28563f
C26866 a_14820_31048# uio_oe[2] 0.00296f
C26867 a_1916_16839# a_2364_16839# 0.0131f
C26868 _328_.A2 a_41776_20072# 0.01407f
C26869 _459_.Q a_32180_23588# 0.002f
C26870 a_35092_16936# a_35204_15748# 0.02666f
C26871 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I a_63404_20408# 0.00103f
C26872 a_33483_29535# uo_out[6] 0.02377f
C26873 a_27028_23588# a_26668_23544# 0.0869f
C26874 a_23556_23208# a_23644_21543# 0.00151f
C26875 a_23532_23544# a_23980_23544# 0.0131f
C26876 _350_.A1 _371_.A3 0.0155f
C26877 vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I 0.69584f
C26878 a_1468_4728# VPWR 0.29679f
C26879 a_14372_31048# VPWR 0.20952f
C26880 a_21876_25156# a_21516_25112# 0.08663f
C26881 a_9892_1256# VPWR 0.20536f
C26882 a_4068_7908# VPWR 0.2157f
C26883 a_39012_1256# a_39460_1256# 0.01328f
C26884 a_18044_2727# a_18492_2727# 0.0131f
C26885 a_53772_13703# a_54132_13800# 0.08707f
C26886 a_67660_13703# a_68108_13703# 0.0131f
C26887 a_1468_17272# a_1468_16839# 0.05841f
C26888 a_43580_27815# a_43008_26795# 0.00105f
C26889 a_40692_27912# a_40464_27165# 0.00186f
C26890 _304_.B _495_.I 0.14614f
C26891 a_54804_25156# a_54444_25112# 0.0869f
C26892 a_40556_16839# a_40916_16936# 0.08707f
C26893 a_62564_29032# a_63336_29480# 0.00647f
C26894 a_4940_23111# a_4964_22020# 0.0016f
C26895 _327_.A2 a_43400_18909# 0.08816f
C26896 _251_.A1 a_61860_26344# 0.00724f
C26897 a_35876_1636# VPWR 0.2085f
C26898 a_67884_16839# VPWR 0.33379f
C26899 a_47524_10664# a_47524_9476# 0.05841f
C26900 _311_.A2 a_37196_23544# 0.01581f
C26901 a_58948_26344# _251_.ZN 0.0184f
C26902 a_38808_27967# VPWR 0.00204f
C26903 a_4964_1636# a_4604_1592# 0.08707f
C26904 a_3172_29860# a_3620_29860# 0.01328f
C26905 a_45416_29885# a_45800_30345# 1.16391f
C26906 a_3172_17316# a_2812_17272# 0.08717f
C26907 _359_.B VPWR 2.87169f
C26908 _352_.A2 a_24636_25641# 0.01093f
C26909 a_58948_11044# a_59036_11000# 0.28563f
C26910 a_53908_16936# a_54356_16936# 0.01328f
C26911 _304_.A1 _327_.A2 0.0137f
C26912 a_48420_1636# a_48868_1636# 0.01328f
C26913 a_55004_11000# a_55452_11000# 0.01288f
C26914 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I 0.00329f
C26915 a_53996_25112# VPWR 0.30195f
C26916 a_58388_17316# a_58028_17272# 0.08674f
C26917 vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I 0.25349f
C26918 a_2276_20072# a_2276_18884# 0.05841f
C26919 a_38472_30169# uo_out[2] 0.0074f
C26920 _419_.A4 a_48084_18884# 0.00202f
C26921 a_20844_26680# _455_.D 0.06383f
C26922 _250_.A2 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN 0.00585f
C26923 a_46180_18504# a_46156_16839# 0.00144f
C26924 a_62980_18884# a_62620_18840# 0.08717f
C26925 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN VPWR 0.90143f
C26926 a_3620_25156# VPWR 0.22347f
C26927 _274_.A1 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN 0.12064f
C26928 a_23308_20408# VPWR 0.31143f
C26929 a_16588_27815# a_17036_27815# 0.0131f
C26930 a_2364_27815# a_2724_27912# 0.08717f
C26931 _350_.A1 uo_out[7] 0.11025f
C26932 a_36636_25112# _444_.D 0.01679f
C26933 a_61412_12612# VPWR 0.20595f
C26934 _383_.ZN _402_.A1 0.02477f
C26935 a_4068_15748# a_4156_15704# 0.28563f
C26936 _402_.A1 a_50068_27508# 0.03663f
C26937 _251_.A1 _267_.A1 0.01324f
C26938 a_18852_2824# a_19300_2824# 0.01328f
C26939 _399_.ZN a_49764_23588# 0.00505f
C26940 a_16700_29383# a_17060_29480# 0.08663f
C26941 a_16252_29383# _467_.D 0.00234f
C26942 a_53660_21543# a_52452_21236# 0.00491f
C26943 _371_.ZN a_28054_30196# 0.05384f
C26944 _311_.A2 a_34304_24029# 0.00152f
C26945 a_36188_25112# a_36212_23588# 0.00117f
C26946 a_53548_24679# clk 0.01875f
C26947 a_5388_8999# a_5300_9096# 0.28563f
C26948 a_61972_10664# VPWR 0.20641f
C26949 a_55004_15271# a_55364_15368# 0.08717f
C26950 a_65756_5863# a_65668_5960# 0.28563f
C26951 _304_.B a_40132_20072# 0.00143f
C26952 a_64860_7431# a_64772_7528# 0.28563f
C26953 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I 0.00225f
C26954 a_66652_4295# a_66564_4392# 0.28563f
C26955 a_36656_29123# VPWR 0.18592f
C26956 _251_.A1 a_62404_25156# 0.0051f
C26957 _474_.Q a_50280_19369# 0.00567f
C26958 a_35428_15368# VPWR 0.20736f
C26959 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN 0.77988f
C26960 a_38876_15271# VPWR 0.32938f
C26961 _441_.B a_39536_23588# 0.00571f
C26962 a_3172_14180# a_2812_14136# 0.08717f
C26963 _304_.B _424_.B1 0.50555f
C26964 a_62560_25112# vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN 0.00405f
C26965 a_63068_17272# VPWR 0.31389f
C26966 a_32292_1256# VPWR 0.20348f
C26967 a_67100_7431# VPWR 0.29679f
C26968 _251_.A1 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.00145f
C26969 _395_.A2 a_51332_24072# 0.00293f
C26970 _260_.ZN a_42784_22504# 0.0011f
C26971 a_37360_19325# a_37408_18504# 0.00139f
C26972 _284_.A2 _398_.C 0.00153f
C26973 a_64972_13703# a_64884_13800# 0.28563f
C26974 _234_.ZN a_39884_27815# 0.00354f
C26975 a_40038_28720# _436_.B 0.02225f
C26976 a_37444_17316# a_37420_16839# 0.00172f
C26977 a_33500_17272# a_33500_16839# 0.05841f
C26978 _495_.I VPWR 1.22814f
C26979 a_15460_31048# VPWR 0.37642f
C26980 a_51756_16839# a_51668_16936# 0.28563f
C26981 a_66004_18504# VPWR 0.27016f
C26982 a_42012_1592# VPWR 0.33609f
C26983 _268_.A2 a_51457_29861# 0.04165f
C26984 a_3620_23208# a_3620_22020# 0.05841f
C26985 a_10428_1159# a_10788_1256# 0.08717f
C26986 a_47412_16936# VPWR 0.20703f
C26987 a_1020_12135# a_1380_12232# 0.08717f
C26988 a_54668_12135# a_55116_12135# 0.01288f
C26989 a_11460_1636# a_11908_1636# 0.01328f
C26990 a_3620_29480# a_4068_29480# 0.01328f
C26991 _452_.CLK a_37532_26680# 0.0211f
C26992 a_25772_23544# a_25884_23111# 0.02634f
C26993 _411_.A2 a_50308_26476# 0.00588f
C26994 a_22636_25112# a_22748_24679# 0.02634f
C26995 a_25420_30345# _349_.A4 0.03037f
C26996 a_32964_17316# a_32604_17272# 0.08707f
C26997 a_22636_30951# uio_out[4] 0.00849f
C26998 _330_.A1 clkload0.Z 0.01798f
C26999 a_52540_11000# a_52428_10567# 0.02634f
C27000 a_55140_1636# a_55812_1636# 0.00347f
C27001 a_62308_11044# a_62396_11000# 0.28563f
C27002 _436_.B a_41028_26344# 0.04682f
C27003 a_12356_2824# VPWR 0.22423f
C27004 _294_.ZN a_32380_26247# 0.00435f
C27005 _337_.ZN _335_.ZN 0.0373f
C27006 _304_.B _386_.ZN 0.11912f
C27007 _393_.A3 a_49044_28292# 0.00156f
C27008 _416_.A1 _311_.A2 0.17864f
C27009 _404_.A1 _411_.A2 0.00887f
C27010 a_32144_26724# VPWR 0.01407f
C27011 a_17036_24679# a_17484_24679# 0.0131f
C27012 _459_.CLK a_17396_26344# 0.00641f
C27013 a_68020_20452# a_68108_20408# 0.28563f
C27014 a_60380_1159# a_60828_1159# 0.0131f
C27015 a_65892_15368# VPWR 0.23142f
C27016 _455_.Q a_21424_25987# 0.00123f
C27017 a_1468_18407# a_1916_18407# 0.0131f
C27018 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I VPWR 0.74919f
C27019 a_21964_25112# VPWR 0.34385f
C27020 _288_.ZN a_35818_29860# 0.02549f
C27021 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I 0.00125f
C27022 _255_.ZN _255_.I 0.49258f
C27023 _427_.ZN vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I 0.00885f
C27024 a_33860_15748# a_33948_15704# 0.28563f
C27025 a_37444_15748# a_37892_15748# 0.01328f
C27026 a_48060_12135# VPWR 0.29679f
C27027 a_47524_18504# a_47388_17272# 0.00154f
C27028 a_21852_2727# a_21988_1636# 0.00154f
C27029 a_51220_18504# a_51332_17316# 0.02666f
C27030 _281_.ZN a_51108_21640# 0.01788f
C27031 a_59260_23111# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I 0.0026f
C27032 a_1468_24679# VPWR 0.29679f
C27033 a_40132_20072# VPWR 0.20593f
C27034 _452_.CLK a_44812_16839# 0.00239f
C27035 a_31172_15748# VPWR 0.20348f
C27036 _293_.A2 a_38584_28292# 0.0242f
C27037 _324_.C a_56572_29383# 0.00292f
C27038 _424_.B1 a_52652_18407# 0.00273f
C27039 a_44752_18147# a_45820_18407# 0.00506f
C27040 a_27028_22020# a_27116_21976# 0.28563f
C27041 a_23084_21976# a_23532_21976# 0.01288f
C27042 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I clk 0.01145f
C27043 _324_.C a_45156_21236# 0.00487f
C27044 _424_.B1 VPWR 3.4092f
C27045 a_48844_16839# a_49292_16839# 0.01288f
C27046 a_47524_14180# a_47164_14136# 0.08707f
C27047 a_42572_16839# VPWR 0.36942f
C27048 a_48708_29816# a_49112_29885# 0.41635f
C27049 a_51956_26183# a_52360_26355# 0.41635f
C27050 a_61188_1256# a_61860_1256# 0.00347f
C27051 _371_.ZN _373_.A2 0.64265f
C27052 a_54692_1256# VPWR 0.20348f
C27053 a_40444_2727# a_40892_2727# 0.0131f
C27054 _416_.A3 a_45820_18840# 0.00166f
C27055 _397_.A4 _474_.Q 0.00808f
C27056 a_61524_13800# a_61972_13800# 0.01328f
C27057 _474_.CLK a_55788_25112# 0.01003f
C27058 a_44459_18559# a_44276_17316# 0.00123f
C27059 a_58687_31220# VPWR 0.58575f
C27060 a_33052_17272# VPWR 0.29736f
C27061 a_5300_10664# a_5388_8999# 0.0027f
C27062 a_35723_20569# a_35968_20937# 0.00232f
C27063 a_21316_23208# a_21428_22020# 0.02666f
C27064 _416_.A2 a_47259_20127# 0.09862f
C27065 a_55812_1636# VPWR 0.22925f
C27066 a_21852_1159# a_21764_1256# 0.28563f
C27067 a_51980_12135# a_51892_12232# 0.28563f
C27068 _402_.A1 a_44744_26355# 0.06719f
C27069 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I 0.00384f
C27070 a_63336_29480# _250_.B 0.00357f
C27071 _441_.ZN _441_.A2 0.18836f
C27072 a_9308_29816# a_9756_29816# 0.01288f
C27073 a_13252_29860# a_13340_29816# 0.28563f
C27074 _251_.A1 a_58276_25156# 0.00405f
C27075 a_9220_29860# uio_oe[5] 0.00193f
C27076 _336_.A1 a_28372_23588# 0.01864f
C27077 a_34532_2824# VPWR 0.21829f
C27078 a_59484_11000# a_59372_10567# 0.02634f
C27079 a_58500_1636# a_58588_1592# 0.28563f
C27080 a_62084_1636# a_62532_1636# 0.01328f
C27081 a_1916_10567# a_2364_10567# 0.0131f
C27082 _386_.ZN VPWR 0.39435f
C27083 _393_.ZN _416_.A1 0.05582f
C27084 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN a_57692_14136# 0.00328f
C27085 _424_.A1 _419_.Z 0.93237f
C27086 a_15692_23111# a_16052_23208# 0.08717f
C27087 a_27900_23111# a_28348_23111# 0.01288f
C27088 a_19612_24679# a_19972_24776# 0.08707f
C27089 _444_.D _439_.ZN 0.00276f
C27090 a_1916_9432# VPWR 0.297f
C27091 a_47612_14136# VPWR 0.29679f
C27092 a_52228_2824# a_52092_1592# 0.00154f
C27093 a_11684_2824# a_11772_1159# 0.0027f
C27094 a_1020_21543# a_1468_21543# 0.0131f
C27095 _400_.ZN a_44340_26183# 0.00221f
C27096 _442_.ZN a_39772_26247# 0.04763f
C27097 a_39536_26795# a_40220_26247# 0.00107f
C27098 a_32156_18407# a_32068_18504# 0.28563f
C27099 a_37108_23588# a_36748_23544# 0.0869f
C27100 _431_.A3 _260_.A2 0.15291f
C27101 a_17508_29860# uio_out[7] 0.00531f
C27102 a_56964_26724# a_58052_26724# 0.01618f
C27103 a_26916_31048# _349_.A4 0.00135f
C27104 a_54916_21640# a_54892_19975# 0.00131f
C27105 a_2276_12232# VPWR 0.20634f
C27106 a_50076_15704# a_50212_15368# 0.00168f
C27107 a_41252_2824# a_41700_2824# 0.01328f
C27108 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I a_61748_23588# 0.0029f
C27109 _363_.Z _287_.A1 0.12475f
C27110 _316_.ZN a_34732_19975# 0.00102f
C27111 a_15156_24776# VPWR 0.20348f
C27112 VPWR uio_out[4] 0.2719f
C27113 _290_.ZN _459_.CLK 0.02873f
C27114 _270_.A2 _237_.A1 0.37694f
C27115 a_1916_2727# a_1828_2824# 0.28563f
C27116 a_44836_15748# VPWR 0.20703f
C27117 a_3260_19975# a_3620_20072# 0.08717f
C27118 a_4604_18840# a_4516_17316# 0.0027f
C27119 a_47972_9476# a_48420_9476# 0.01328f
C27120 a_61836_25515# vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN 0.01164f
C27121 a_46628_9476# a_46268_9432# 0.08717f
C27122 _455_.Q _351_.ZN 0.00794f
C27123 _438_.A2 a_38628_25156# 0.00414f
C27124 a_54020_14180# a_54468_14180# 0.01328f
C27125 _257_.B a_59572_29076# 0.39851f
C27126 _304_.B a_53212_27815# 0.02218f
C27127 _223_.I a_30724_26020# 0.00618f
C27128 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I a_66764_20408# 0.00144f
C27129 a_2724_12612# a_2812_12568# 0.28563f
C27130 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_63180_26680# 0.00158f
C27131 a_37324_28776# uo_out[7] 0.00106f
C27132 a_35232_24029# a_34939_23705# 0.49319f
C27133 _416_.A3 a_47076_18504# 0.00774f
C27134 a_52652_18407# a_52676_17316# 0.0016f
C27135 a_50524_17272# a_50412_16839# 0.02634f
C27136 a_28260_23208# a_28372_22020# 0.02666f
C27137 _437_.A1 a_39587_24372# 0.00436f
C27138 a_52676_17316# VPWR 0.20672f
C27139 a_24452_23208# a_24428_21976# 0.0016f
C27140 a_29232_29931# a_30795_29977# 0.41635f
C27141 a_62508_12135# a_62868_12232# 0.08707f
C27142 a_65084_1592# VPWR 0.30253f
C27143 a_32828_1159# a_33188_1256# 0.08717f
C27144 a_59932_12568# a_59844_11044# 0.00151f
C27145 a_53212_29816# a_54000_30344# 0.00403f
C27146 a_48420_12232# a_49204_12232# 0.00276f
C27147 _229_.I a_61500_27815# 0.00722f
C27148 a_17596_1592# a_18044_1592# 0.01288f
C27149 a_21540_1636# a_21628_1592# 0.28563f
C27150 _362_.ZN _371_.A1 0.09484f
C27151 _424_.B1 a_50068_27508# 0.47376f
C27152 _419_.Z _416_.A2 0.03336f
C27153 _287_.A1 a_33812_29860# 0.0141f
C27154 a_17956_29860# _459_.CLK 0.01953f
C27155 a_25436_21543# VPWR 0.31768f
C27156 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I a_59260_23544# 0.01323f
C27157 a_51332_24072# _427_.A2 0.87003f
C27158 _398_.C a_52452_24072# 0.04987f
C27159 a_41924_1636# a_41788_1159# 0.00168f
C27160 a_56348_11000# a_56372_10664# 0.00172f
C27161 _384_.A3 _384_.A1 0.61798f
C27162 _455_.Q _337_.A3 3.24089f
C27163 a_56932_2824# VPWR 0.21171f
C27164 a_2724_2824# a_2724_1636# 0.05841f
C27165 _411_.A2 a_48384_26724# 0.07191f
C27166 a_27004_23111# a_26916_23208# 0.28563f
C27167 a_62732_26680# VPWR 0.32647f
C27168 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I 0.01436f
C27169 a_21764_24776# a_22212_24776# 0.01328f
C27170 _337_.ZN a_30596_28292# 0.01381f
C27171 a_56036_9476# VPWR 0.21311f
C27172 a_63204_14180# VPWR 0.20952f
C27173 _336_.A2 a_27452_23111# 0.00361f
C27174 _452_.CLK a_36172_24463# 0.00255f
C27175 _424_.B1 _424_.B2 0.38495f
C27176 a_13364_31048# a_13252_29860# 0.02666f
C27177 _397_.A4 _395_.A2 0.00277f
C27178 a_41160_29083# _265_.ZN 0.01087f
C27179 _218_.ZN VPWR 1.32972f
C27180 a_43580_15704# a_44028_15704# 0.01288f
C27181 a_63764_12232# VPWR 0.20622f
C27182 a_33312_28776# uo_out[6] 0.00144f
C27183 _473_.Q a_49604_22020# 0.02145f
C27184 a_35060_20569# VPWR 0.00388f
C27185 a_22064_27912# _454_.D 0.3043f
C27186 _359_.B _370_.B 0.22285f
C27187 a_62620_18840# a_62620_18407# 0.05841f
C27188 a_67012_18884# a_66988_18407# 0.00172f
C27189 _397_.A4 a_46984_23588# 0.23433f
C27190 a_1828_18884# VPWR 0.20348f
C27191 _459_.D a_30240_24776# 0.2496f
C27192 a_12892_2727# a_13252_2824# 0.08717f
C27193 _304_.B _386_.A4 0.47192f
C27194 _324_.C _324_.B 1.7325f
C27195 a_50972_15704# VPWR 0.33271f
C27196 _438_.A2 _302_.Z 0.02849f
C27197 a_64860_19975# a_65308_19975# 0.01222f
C27198 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I a_65668_27912# 0.02229f
C27199 _355_.C a_23868_26247# 0.01553f
C27200 a_43156_20452# _325_.B 0.00196f
C27201 _301_.A1 a_37532_21543# 0.0082f
C27202 _465_.D uio_out[7] 0.0127f
C27203 a_1380_20452# a_1020_20408# 0.08717f
C27204 _447_.Q a_39475_21236# 0.00122f
C27205 a_3172_20452# a_3620_20452# 0.01328f
C27206 a_47836_17272# a_47748_15748# 0.00151f
C27207 _355_.C a_19035_28409# 0.03457f
C27208 _319_.A3 a_38788_20072# 0.00188f
C27209 _336_.Z a_28460_23544# 0.00612f
C27210 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN 0.00304f
C27211 a_53212_27815# VPWR 0.3264f
C27212 a_62844_2727# a_63292_2727# 0.0131f
C27213 a_50660_12612# a_51108_12612# 0.01328f
C27214 a_47076_12612# a_47164_12568# 0.28563f
C27215 a_67996_18840# a_67908_17316# 0.00151f
C27216 _397_.A1 a_46356_24072# 0.08794f
C27217 a_40038_28720# a_40464_27165# 0.00132f
C27218 a_20060_1159# VPWR 0.33357f
C27219 a_31620_20072# a_32068_20072# 0.01328f
C27220 a_65220_9096# a_65220_7908# 0.05841f
C27221 a_44252_1159# a_44164_1256# 0.28563f
C27222 a_67012_5960# a_67012_4772# 0.05841f
C27223 a_63292_12568# a_63204_11044# 0.00151f
C27224 a_66116_7528# a_66116_6340# 0.05841f
C27225 a_24900_1636# a_24540_1592# 0.08707f
C27226 a_22660_21640# VPWR 0.20614f
C27227 a_36636_26247# a_37084_26247# 0.01222f
C27228 a_51420_17272# a_51868_17272# 0.01288f
C27229 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I a_56260_14180# 0.00137f
C27230 _435_.A3 a_40084_25156# 0.00174f
C27231 _350_.A1 _340_.A2 0.6619f
C27232 a_49740_10567# a_50100_10664# 0.08707f
C27233 a_43888_19204# a_44300_19001# 0.00275f
C27234 a_63404_10567# a_63852_10567# 0.01288f
C27235 _395_.A2 a_51956_26183# 0.00417f
C27236 a_4156_1159# a_4828_1159# 0.00544f
C27237 _325_.A2 a_36836_20072# 0.00396f
C27238 a_47476_28292# VPWR 0.01382f
C27239 _467_.D a_16588_26247# 0.00831f
C27240 _424_.B1 a_51240_23340# 0.18367f
C27241 a_61524_23208# VPWR 0.20915f
C27242 a_25348_23208# a_25796_23208# 0.01328f
C27243 _474_.CLK vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I 0.03522f
C27244 _304_.B a_42982_21730# 0.05723f
C27245 a_20084_23588# VPWR 0.20622f
C27246 a_67012_9476# VPWR 0.20677f
C27247 _304_.B _407_.A1 0.4587f
C27248 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN VPWR 0.782f
C27249 a_67908_2824# a_67772_1592# 0.00154f
C27250 _459_.CLK a_22620_27599# 0.02285f
C27251 a_50188_13703# VPWR 0.33011f
C27252 a_20060_21543# a_19972_21640# 0.28563f
C27253 a_31932_21543# a_32380_21543# 0.01288f
C27254 a_20003_29611# a_19328_28733# 0.02345f
C27255 a_65756_6296# VPWR 0.31505f
C27256 a_18628_26344# a_18716_24679# 0.00151f
C27257 _350_.A1 _459_.Q 1.44315f
C27258 a_67548_3160# VPWR 0.29679f
C27259 a_39236_26344# VPWR 0.12826f
C27260 _455_.Q a_21044_27508# 0.29732f
C27261 _290_.ZN uo_out[7] 0.02798f
C27262 a_27588_26724# a_28036_26724# 0.01328f
C27263 _287_.A1 uo_out[3] 0.00218f
C27264 a_50884_15748# a_50524_15704# 0.08707f
C27265 a_45372_11000# VPWR 0.30073f
C27266 a_13788_29816# a_13788_29383# 0.05841f
C27267 a_63652_2824# a_64100_2824# 0.01328f
C27268 a_48308_23588# a_49764_23588# 0.01731f
C27269 a_932_26724# VPWR 0.22176f
C27270 _250_.C a_60852_28292# 0.00126f
C27271 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_60964_27912# 0.00187f
C27272 _474_.CLK _419_.A4 0.0381f
C27273 a_60940_15704# a_61388_15704# 0.01222f
C27274 a_31284_20452# a_31260_19975# 0.00172f
C27275 _330_.A2 VPWR 1.05056f
C27276 a_44700_30951# vgaringosc.workerclkbuff_notouch_.I 0.00613f
C27277 a_3620_26344# VPWR 0.22347f
C27278 a_24316_2727# a_24228_2824# 0.28563f
C27279 _386_.A4 VPWR 1.10588f
C27280 _384_.ZN _395_.A3 0.00127f
C27281 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN VPWR 0.94837f
C27282 _460_.Q a_35140_26680# 0.26661f
C27283 _350_.A2 a_29788_30345# 0.01143f
C27284 a_57604_9476# a_57244_9432# 0.08717f
C27285 a_58948_9476# a_59396_9476# 0.01328f
C27286 a_4964_28292# VPWR 0.2136f
C27287 a_5636_31048# a_6084_31048# 0.01328f
C27288 _223_.I _337_.ZN 0.05011f
C27289 _436_.B a_39796_27912# 0.01422f
C27290 a_5188_1256# a_5636_1256# 0.01328f
C27291 _287_.A2 _371_.A1 0.32903f
C27292 a_1380_4772# a_1828_4772# 0.01328f
C27293 a_66340_14180# a_65980_14136# 0.08707f
C27294 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN a_55140_15748# 0.00254f
C27295 a_62396_14136# a_62844_14136# 0.01288f
C27296 a_2276_3204# a_2724_3204# 0.01328f
C27297 a_16948_20452# a_17036_20408# 0.28563f
C27298 a_35008_22461# a_34715_22137# 0.49319f
C27299 _355_.C uio_out[7] 0.0838f
C27300 _328_.A2 _325_.ZN 0.00666f
C27301 _350_.A1 _461_.D 0.00514f
C27302 a_22524_1592# a_22660_1256# 0.00168f
C27303 a_1828_1636# VPWR 0.20348f
C27304 a_52788_13800# a_52876_12135# 0.0027f
C27305 a_21740_29383# VPWR 0.31436f
C27306 _359_.B _360_.ZN 0.00105f
C27307 a_23108_29860# a_23196_29816# 0.28563f
C27308 a_5052_29816# a_5188_29480# 0.00168f
C27309 a_55228_1159# a_55588_1256# 0.08717f
C27310 a_53796_20452# VPWR 0.21208f
C27311 a_42236_1159# VPWR 0.36726f
C27312 a_63180_16839# a_63628_16839# 0.0131f
C27313 _397_.A2 _404_.A1 0.47485f
C27314 a_31260_1592# a_31708_1592# 0.012f
C27315 a_2724_11044# a_3172_11044# 0.01328f
C27316 a_42392_19243# _452_.D 0.00102f
C27317 a_47483_20569# a_47728_20937# 0.00232f
C27318 a_47776_20893# a_49068_20408# 0.00704f
C27319 a_40780_27815# a_41228_27815# 0.01222f
C27320 _229_.I a_61860_27912# 0.00521f
C27321 _252_.B a_59260_26680# 0.00803f
C27322 a_60716_10567# a_60628_10664# 0.28563f
C27323 a_3172_18504# a_3172_17316# 0.05841f
C27324 _281_.ZN _417_.A2 0.2663f
C27325 _452_.Q a_39536_23588# 0.00148f
C27326 a_67684_24776# vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN 0.00205f
C27327 a_39300_31048# uo_out[1] 0.00331f
C27328 _293_.A2 uo_out[3] 0.00645f
C27329 a_54020_21640# a_54468_21640# 0.01328f
C27330 a_20980_22020# VPWR 0.20622f
C27331 _246_.B2 ui_in[3] 0.0032f
C27332 a_42982_21730# VPWR 0.76716f
C27333 a_27564_23544# VPWR 0.32115f
C27334 _407_.A1 VPWR 0.94813f
C27335 a_3708_18840# a_4156_18840# 0.0131f
C27336 a_30588_21543# a_30948_21640# 0.08707f
C27337 a_22300_2727# VPWR 0.31143f
C27338 a_57020_23111# VPWR 0.33882f
C27339 a_4068_13800# VPWR 0.22146f
C27340 _459_.Q a_33396_26344# 0.00102f
C27341 a_22548_31048# a_22636_29383# 0.002f
C27342 a_58388_20452# a_58476_20408# 0.28563f
C27343 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN a_61388_16839# 0.00633f
C27344 a_7204_29860# VPWR 0.20641f
C27345 _238_.I _250_.C 0.00454f
C27346 a_41116_26247# a_41476_26344# 0.08674f
C27347 a_59036_11000# VPWR 0.31547f
C27348 a_19188_22020# a_19164_21543# 0.00172f
C27349 a_63964_15704# a_63964_15271# 0.05841f
C27350 a_15244_21976# a_15244_21543# 0.05841f
C27351 _267_.A1 a_55676_28248# 0.0246f
C27352 a_1020_23111# VPWR 0.30073f
C27353 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.00935f
C27354 a_1380_27912# VPWR 0.20348f
C27355 _431_.A3 _311_.A2 0.42009f
C27356 _437_.A1 _438_.A2 0.82041f
C27357 _296_.ZN a_37386_31048# 0.02604f
C27358 a_35292_2727# a_35652_2824# 0.08717f
C27359 a_56036_23208# a_56484_23208# 0.01328f
C27360 a_62508_23111# a_62868_23208# 0.08717f
C27361 _478_.D a_54040_22366# 0.01057f
C27362 a_49896_18909# a_50816_19369# 0.00306f
C27363 _334_.A1 a_35874_27937# 0.00102f
C27364 a_1468_4728# a_1468_4295# 0.05841f
C27365 a_64772_4772# a_64412_4728# 0.08717f
C27366 a_2364_3160# a_2364_2727# 0.05841f
C27367 a_65668_3204# a_65308_3160# 0.08717f
C27368 a_22324_20452# a_22772_20452# 0.01328f
C27369 _251_.A1 a_61948_26247# 0.01216f
C27370 a_8627_30644# a_8996_31048# 0.02397f
C27371 a_58588_26247# a_58500_26344# 0.28563f
C27372 _384_.ZN a_47525_29480# 0.08453f
C27373 _383_.ZN _386_.A4 0.03248f
C27374 _304_.B _304_.A1 0.02901f
C27375 _409_.ZN _408_.ZN 0.00191f
C27376 a_56796_12568# a_57244_12568# 0.01288f
C27377 a_15492_1636# VPWR 0.20348f
C27378 _460_.Q _460_.D 0.00586f
C27379 a_39772_26247# _441_.ZN 0.00221f
C27380 _459_.CLK a_25936_25597# 0.00906f
C27381 _459_.CLK uio_out[5] 0.00275f
C27382 a_66092_19975# a_66116_18884# 0.0016f
C27383 a_59708_23111# a_59620_23208# 0.28563f
C27384 _359_.B a_28556_29167# 0.05562f
C27385 a_4156_19975# VPWR 0.3269f
C27386 _330_.ZN a_38316_16839# 0.00543f
C27387 a_37408_18504# a_38764_16839# 0.00103f
C27388 a_64636_1159# VPWR 0.30056f
C27389 a_66652_1159# a_66564_1256# 0.28563f
C27390 a_38564_1636# a_38204_1592# 0.08707f
C27391 _435_.A3 _430_.ZN 0.15339f
C27392 a_1828_5960# VPWR 0.20348f
C27393 a_30812_18407# VPWR 0.30073f
C27394 _447_.Q _448_.Q 2.66708f
C27395 _384_.A3 clk 0.03556f
C27396 a_28000_29480# _371_.A2 0.00208f
C27397 a_57492_10664# a_57940_10664# 0.01328f
C27398 _325_.A2 a_44724_17316# 0.0013f
C27399 a_24228_26344# VPWR 0.2061f
C27400 a_63616_31128# a_64324_29860# 0.01792f
C27401 a_26556_1159# a_27004_1159# 0.0131f
C27402 _330_.ZN a_36548_17316# 0.00116f
C27403 a_45396_28292# VPWR 0.21523f
C27404 a_19524_24776# a_19612_23111# 0.00151f
C27405 _274_.A1 a_56036_28292# 0.03541f
C27406 a_54892_25112# a_54892_24679# 0.05841f
C27407 a_27116_21976# VPWR 0.36324f
C27408 a_1020_26680# a_1020_26247# 0.05841f
C27409 _229_.I _247_.ZN 0.22146f
C27410 a_29156_21640# a_29604_21640# 0.01328f
C27411 a_35504_18955# a_36060_19369# 0.8399f
C27412 a_13788_29816# uio_oe[2] 0.00697f
C27413 _433_.ZN a_41460_22020# 0.0018f
C27414 a_65780_13800# VPWR 0.22327f
C27415 a_56484_2824# a_56572_1159# 0.0027f
C27416 a_44700_2727# VPWR 0.31143f
C27417 a_4940_26247# a_4852_26344# 0.28563f
C27418 _441_.A2 a_41488_24072# 0.00215f
C27419 a_30724_15368# a_31172_15368# 0.01328f
C27420 a_59955_30600# ui_in[2] 0.02049f
C27421 _241_.Z _242_.Z 0.11544f
C27422 a_13340_29816# VPWR 0.29679f
C27423 a_67348_16936# a_67460_15748# 0.02666f
C27424 a_45820_10567# VPWR 0.29679f
C27425 vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN a_63316_23588# 0.03074f
C27426 a_32604_15271# a_32516_15368# 0.28563f
C27427 a_57020_2727# a_57156_1636# 0.00154f
C27428 _272_.A2 a_57220_29861# 0.0142f
C27429 a_31932_23111# VPWR 0.31555f
C27430 _419_.A4 _398_.C 0.02245f
C27431 _324_.B a_45396_22020# 0.01475f
C27432 _474_.D a_50384_19204# 0.23443f
C27433 a_33948_15271# a_34620_15271# 0.00544f
C27434 _407_.A1 a_50068_27508# 0.20119f
C27435 a_60828_26680# a_61748_26724# 0.00795f
C27436 a_1380_22020# a_1828_22020# 0.01328f
C27437 a_46716_2727# a_46628_2824# 0.28563f
C27438 vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN a_64772_26344# 0.00591f
C27439 a_43400_18909# VPWR 1.10301f
C27440 a_31920_29480# a_32848_29123# 1.16391f
C27441 a_66564_17316# a_67012_17316# 0.01328f
C27442 _399_.ZN _399_.A2 0.9209f
C27443 a_48956_30951# uio_in[1] 0.00318f
C27444 a_62980_17316# a_62620_17272# 0.08717f
C27445 a_50084_24328# a_51332_24372# 0.02129f
C27446 a_27588_1256# a_28036_1256# 0.01328f
C27447 a_66316_20408# a_66452_20072# 0.00168f
C27448 a_67100_7864# a_67100_7431# 0.05841f
C27449 _474_.CLK vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I 0.02269f
C27450 a_2812_8999# a_3260_8999# 0.0131f
C27451 a_3708_7431# a_4156_7431# 0.0131f
C27452 a_18828_23544# a_19276_23544# 0.01288f
C27453 a_33508_31048# VPWR 0.01455f
C27454 a_64412_4295# a_64860_4295# 0.0131f
C27455 a_4940_5863# a_5388_5863# 0.01222f
C27456 a_6620_2727# a_7068_2727# 0.0131f
C27457 a_56460_13703# a_57132_13703# 0.00544f
C27458 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN a_59652_25640# 0.084f
C27459 a_2812_13703# a_3172_13800# 0.08717f
C27460 _223_.I a_30795_29977# 0.00894f
C27461 a_27924_20452# a_28012_20408# 0.28563f
C27462 a_38676_16936# a_38876_15271# 0.00119f
C27463 a_4156_16839# a_4852_16936# 0.01227f
C27464 _304_.A1 VPWR 2.93167f
C27465 a_21628_1592# VPWR 0.3289f
C27466 _427_.B1 a_53908_24776# 0.00112f
C27467 a_64100_12612# a_64188_12568# 0.28563f
C27468 a_10092_30951# a_10540_30951# 0.01222f
C27469 a_1916_23544# a_1916_23111# 0.05841f
C27470 _404_.A1 _330_.A1 0.00811f
C27471 a_67324_15271# a_67236_15368# 0.28563f
C27472 _267_.A2 _246_.B2 0.0389f
C27473 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I 0.02277f
C27474 a_51644_11000# a_52092_11000# 0.01288f
C27475 _359_.B a_41056_30669# 0.00263f
C27476 _264_.B a_41642_25156# 0.0014f
C27477 a_42932_16936# a_43380_16936# 0.01328f
C27478 a_41476_1636# a_41564_1592# 0.28563f
C27479 a_45060_1636# a_45508_1636# 0.01328f
C27480 _397_.A2 a_48384_26724# 0.11369f
C27481 a_2812_26680# a_3260_26680# 0.0131f
C27482 _245_.I1 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I 0.00237f
C27483 a_22548_29480# VPWR 0.20348f
C27484 a_4852_21640# a_4940_19975# 0.00151f
C27485 a_2812_20408# VPWR 0.30213f
C27486 _452_.CLK a_31844_23208# 0.0036f
C27487 a_67100_2727# VPWR 0.29679f
C27488 a_47164_12568# VPWR 0.29679f
C27489 _452_.Q a_42610_21812# 0.00122f
C27490 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.00379f
C27491 hold2.Z _451_.Q 0.27317f
C27492 a_7516_2727# a_7652_1636# 0.00154f
C27493 a_7428_2824# a_7876_2824# 0.01328f
C27494 _267_.ZN a_52316_27815# 0.00243f
C27495 a_5276_29383# a_5636_29480# 0.08717f
C27496 _251_.A1 a_60656_29612# 0.00126f
C27497 _416_.A3 _421_.B 0.4452f
C27498 _448_.D VPWR 0.41936f
C27499 _324_.C _403_.ZN 0.74188f
C27500 a_1916_28248# a_1916_27815# 0.05841f
C27501 a_67660_10567# VPWR 0.31389f
C27502 a_31820_21976# a_31932_21543# 0.02634f
C27503 _274_.A1 a_53616_29480# 0.00171f
C27504 a_43580_15271# a_43940_15368# 0.08717f
C27505 a_29604_23208# VPWR 0.20595f
C27506 _390_.ZN a_52316_27815# 0.02258f
C27507 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I 0.00272f
C27508 _324_.C a_56124_28248# 0.00977f
C27509 a_16052_28292# a_16500_28292# 0.01328f
C27510 a_15156_28292# a_15244_28248# 0.28563f
C27511 a_57468_2727# a_58052_2824# 0.01675f
C27512 _459_.Q a_31732_23588# 0.002f
C27513 _328_.A2 a_41572_20072# 0.00395f
C27514 a_65220_15748# VPWR 0.21168f
C27515 _327_.Z _450_.D 0.03997f
C27516 a_14372_31048# uio_oe[2] 0.01582f
C27517 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN a_65756_23111# 0.00184f
C27518 _245_.I1 a_60212_25156# 0.0014f
C27519 a_56684_23544# clk 0.00613f
C27520 a_61188_15368# a_61636_15368# 0.01328f
C27521 a_32476_29167# uo_out[6] 0.00207f
C27522 a_53460_18504# a_53908_18504# 0.01328f
C27523 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I VPWR 0.94317f
C27524 a_9444_1256# VPWR 0.20348f
C27525 a_3620_7908# VPWR 0.22347f
C27526 a_26580_23588# a_26668_23544# 0.28563f
C27527 a_13364_31048# VPWR 0.20843f
C27528 a_17484_25112# a_17932_25112# 0.01288f
C27529 a_21428_25156# a_21516_25112# 0.28563f
C27530 a_1020_4728# VPWR 0.30073f
C27531 a_53772_13703# a_53684_13800# 0.28563f
C27532 a_31260_18840# a_31260_18407# 0.05841f
C27533 a_49652_16936# a_49852_15271# 0.00119f
C27534 a_27004_30951# a_27668_31048# 0.00401f
C27535 a_54356_25156# a_54444_25112# 0.28563f
C27536 a_40556_16839# a_40468_16936# 0.28563f
C27537 a_41056_30669# _495_.I 0.02868f
C27538 _251_.A1 a_61412_26344# 0.00725f
C27539 _311_.A2 a_36748_23544# 0.01311f
C27540 a_67436_16839# VPWR 0.31389f
C27541 a_35428_1636# VPWR 0.21238f
C27542 a_58500_26344# _251_.ZN 0.00573f
C27543 a_4516_1636# a_4604_1592# 0.28563f
C27544 a_37860_27967# VPWR 0.00246f
C27545 a_3708_12135# a_4156_12135# 0.0131f
C27546 a_17932_23544# a_17932_23111# 0.05841f
C27547 a_21876_23588# a_21852_23111# 0.00172f
C27548 _474_.CLK _381_.A2 0.15395f
C27549 vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN clk 0.00202f
C27550 a_2724_17316# a_2812_17272# 0.28563f
C27551 a_45012_29816# _393_.ZN 0.00115f
C27552 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I VPWR 0.78284f
C27553 a_61524_12232# a_61612_10567# 0.00151f
C27554 a_58948_11044# a_58588_11000# 0.08707f
C27555 a_20644_1636# a_20508_1159# 0.00168f
C27556 a_16700_1592# a_16700_1159# 0.05841f
C27557 _352_.A2 a_25008_25597# 0.02039f
C27558 a_46794_25156# VPWR 0.01473f
C27559 a_57940_17316# a_58028_17272# 0.28563f
C27560 a_20396_26680# _455_.D 0.01204f
C27561 a_53436_18840# a_53548_18407# 0.02634f
C27562 a_48956_1159# a_49404_1159# 0.0131f
C27563 a_37892_2824# a_37756_1592# 0.00154f
C27564 a_14708_27912# a_14708_26724# 0.05841f
C27565 a_54692_18884# VPWR 0.20834f
C27566 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I 0.01956f
C27567 a_62532_18884# a_62620_18840# 0.28563f
C27568 a_66564_18884# a_67012_18884# 0.01328f
C27569 a_3172_25156# VPWR 0.20993f
C27570 a_2364_27815# a_2276_27912# 0.28563f
C27571 _250_.C VPWR 0.8066f
C27572 a_22860_20408# VPWR 0.31143f
C27573 a_36188_25112# _444_.D 0.02051f
C27574 _459_.Q _290_.ZN 0.031f
C27575 _435_.A3 _441_.A3 0.01594f
C27576 a_4068_15748# a_3708_15704# 0.08717f
C27577 a_60964_12612# VPWR 0.2267f
C27578 a_1468_15704# a_1916_15704# 0.0131f
C27579 a_35740_15704# a_35876_15368# 0.00168f
C27580 a_16700_29383# a_16612_29480# 0.28563f
C27581 _399_.ZN a_49316_23588# 0.00343f
C27582 a_52900_15368# a_53572_15368# 0.00347f
C27583 _371_.ZN a_26427_29977# 0.00108f
C27584 a_28124_30600# a_28054_30196# 0.01746f
C27585 a_64412_7431# a_64772_7528# 0.08717f
C27586 a_61524_10664# VPWR 0.20641f
C27587 a_30476_21976# a_30500_21640# 0.00172f
C27588 a_4940_8999# a_5300_9096# 0.08674f
C27589 a_55004_15271# a_54916_15368# 0.28563f
C27590 a_66204_4295# a_66564_4392# 0.08717f
C27591 a_65308_5863# a_65668_5960# 0.08717f
C27592 _474_.Q a_50384_19204# 0.00744f
C27593 a_35728_29480# VPWR 1.10134f
C27594 a_34980_15368# VPWR 0.2406f
C27595 a_56348_15271# a_56796_15271# 0.0131f
C27596 _251_.A1 a_60416_25156# 0.00389f
C27597 _284_.A2 a_50176_26724# 0.003f
C27598 a_19724_21976# a_20172_21976# 0.01288f
C27599 a_38428_15271# VPWR 0.33333f
C27600 _441_.B a_39332_23588# 0.00259f
C27601 a_2724_14180# a_2812_14136# 0.28563f
C27602 a_37868_16839# a_38316_16839# 0.01288f
C27603 a_27116_23544# a_27028_22020# 0.00151f
C27604 a_41812_16936# a_41700_15748# 0.02666f
C27605 a_62620_17272# VPWR 0.31389f
C27606 a_31372_23544# a_31820_23544# 0.01255f
C27607 a_66652_7431# VPWR 0.29679f
C27608 a_49764_1256# a_50436_1256# 0.00347f
C27609 _424_.A2 hold2.I 0.05484f
C27610 a_31844_1256# VPWR 0.20348f
C27611 _395_.A2 a_50940_24072# 0.00222f
C27612 a_65220_3204# a_65084_2727# 0.00168f
C27613 a_29020_2727# a_29468_2727# 0.0131f
C27614 a_64300_13703# a_64884_13800# 0.01675f
C27615 _245_.I1 VPWR 1.14292f
C27616 a_51048_26680# _398_.C 0.38838f
C27617 a_50548_13800# a_50996_13800# 0.01328f
C27618 a_40038_28720# a_39884_27815# 0.00866f
C27619 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN 0.0121f
C27620 a_14908_30951# VPWR 0.32203f
C27621 a_40644_31048# VPWR 0.01492f
C27622 input9.Z ui_in[5] 0.00228f
C27623 a_51308_16839# a_51668_16936# 0.08717f
C27624 a_65220_18504# VPWR 0.21513f
C27625 _244_.Z a_60276_26724# 0.00129f
C27626 _287_.A1 _294_.ZN 2.09735f
C27627 _334_.A1 _288_.ZN 0.01298f
C27628 _352_.ZN _457_.D 0.63602f
C27629 a_41564_1592# VPWR 0.33368f
C27630 a_10428_1159# a_10340_1256# 0.28563f
C27631 a_50748_1592# a_50884_1256# 0.00168f
C27632 a_46964_16936# VPWR 0.20703f
C27633 a_54580_10664# a_54692_9476# 0.02666f
C27634 a_1020_12135# a_932_12232# 0.28563f
C27635 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I a_57940_18884# 0.00106f
C27636 _452_.CLK a_37084_26680# 0.0211f
C27637 a_58028_20408# a_57940_18884# 0.0027f
C27638 a_48516_24080# _399_.A2 0.00133f
C27639 a_5948_29816# a_6396_29816# 0.01288f
C27640 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I clk 0.06018f
C27641 a_25792_30301# _349_.A4 0.01974f
C27642 a_32516_17316# a_32604_17272# 0.28563f
C27643 a_36100_17316# a_36548_17316# 0.01328f
C27644 a_22188_30951# uio_out[4] 0.00877f
C27645 a_65444_11044# a_65892_11044# 0.01328f
C27646 a_62308_11044# a_61948_11000# 0.08707f
C27647 _330_.A1 a_48384_26724# 0.02829f
C27648 a_48196_15368# a_48060_14136# 0.00154f
C27649 a_52004_15368# a_52004_14180# 0.05841f
C27650 _436_.B a_40580_26344# 0.01491f
C27651 a_11684_2824# VPWR 0.24925f
C27652 a_55140_1636# a_55228_1592# 0.28563f
C27653 a_51196_1592# a_51644_1592# 0.01288f
C27654 _304_.A1 a_36636_21543# 0.03208f
C27655 _393_.A3 a_48820_28292# 0.00234f
C27656 _416_.A1 a_37532_25112# 0.00294f
C27657 a_16588_23111# a_17036_23111# 0.0131f
C27658 _459_.CLK a_16948_26344# 0.00641f
C27659 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN a_54804_18504# 0.05177f
C27660 _421_.A1 _473_.Q 0.21892f
C27661 a_67212_20408# a_68108_20408# 0.00373f
C27662 a_65444_15368# VPWR 0.21032f
C27663 a_5052_4728# a_4964_3204# 0.00151f
C27664 a_58164_18504# VPWR 0.26753f
C27665 a_21516_25112# VPWR 0.31547f
C27666 a_16948_27912# a_17396_27912# 0.01328f
C27667 _452_.CLK _450_.D 0.66995f
C27668 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN a_56708_15368# 0.00126f
C27669 _427_.ZN a_55140_20452# 0.00336f
C27670 a_47612_12135# VPWR 0.29679f
C27671 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN a_62084_18884# 0.00204f
C27672 a_33860_15748# a_33500_15704# 0.08707f
C27673 _251_.A1 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I 0.59218f
C27674 a_29828_2824# a_30276_2824# 0.01328f
C27675 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN 0.00287f
C27676 _397_.A1 _412_.B2 0.36007f
C27677 a_55140_28292# a_55588_28292# 0.01328f
C27678 a_1020_24679# VPWR 0.30073f
C27679 a_44476_15704# a_44476_15271# 0.05841f
C27680 _416_.A3 a_47524_22021# 0.13242f
C27681 a_39684_20072# VPWR 0.20734f
C27682 a_20420_21640# a_20396_20408# 0.0016f
C27683 _452_.CLK a_44364_16839# 0.00239f
C27684 a_30724_15748# VPWR 0.22176f
C27685 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I VPWR 0.81379f
C27686 a_1828_9476# a_2276_9476# 0.01328f
C27687 _260_.ZN a_42982_21730# 0.01724f
C27688 _435_.ZN a_39985_24372# 0.00422f
C27689 a_27028_22020# a_26668_21976# 0.08707f
C27690 a_56148_24776# clk 0.0155f
C27691 a_47600_27912# VPWR 0.01356f
C27692 _304_.B _424_.A2 0.91292f
C27693 a_47076_14180# a_47164_14136# 0.28563f
C27694 a_50660_14180# a_51108_14180# 0.01328f
C27695 a_35652_31048# _288_.ZN 0.00419f
C27696 a_48756_16936# a_48644_15748# 0.02666f
C27697 vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN 0.10099f
C27698 a_47524_31048# _386_.ZN 0.00187f
C27699 a_41900_16839# VPWR 0.33242f
C27700 a_54244_1256# VPWR 0.22423f
C27701 _371_.ZN a_28672_31048# 0.00898f
C27702 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN VPWR 0.73465f
C27703 a_65084_14136# a_64996_12612# 0.00151f
C27704 a_45284_13800# a_45284_12612# 0.05841f
C27705 _474_.CLK a_55340_25112# 0.02464f
C27706 _362_.B a_35204_26344# 0.00214f
C27707 _421_.A1 _475_.D 0.39068f
C27708 a_58519_31220# VPWR 0.00474f
C27709 a_29244_23111# a_29268_22020# 0.0016f
C27710 a_32604_17272# VPWR 0.29679f
C27711 a_21404_1159# a_21764_1256# 0.08717f
C27712 a_61972_10664# a_61860_9476# 0.02666f
C27713 a_55228_1592# VPWR 0.32517f
C27714 a_65420_12135# a_65868_12135# 0.0131f
C27715 a_14596_29480# a_15044_29480# 0.01328f
C27716 a_51532_12135# a_51892_12232# 0.08707f
C27717 a_14236_1592# a_14684_1592# 0.01288f
C27718 a_24428_23544# a_24452_23208# 0.00172f
C27719 a_63336_29480# a_63952_29480# 0.00329f
C27720 a_59348_29076# a_59572_29076# 0.01436f
C27721 a_13252_29860# a_12892_29816# 0.08707f
C27722 _398_.C _381_.A2 0.08831f
C27723 a_40040_17675# a_40644_17272# 0.49241f
C27724 _317_.A2 _319_.A3 0.32538f
C27725 _336_.A1 a_27924_23588# 0.00354f
C27726 a_58500_1636# a_58140_1592# 0.08707f
C27727 a_34084_2824# VPWR 0.20902f
C27728 _335_.ZN _452_.CLK 0.00464f
C27729 a_15692_23111# a_15604_23208# 0.28563f
C27730 a_19612_24679# a_19524_24776# 0.28563f
C27731 a_1380_24776# a_1828_24776# 0.01328f
C27732 a_1468_9432# VPWR 0.29679f
C27733 a_65220_9096# a_65668_9096# 0.01328f
C27734 a_66116_7528# a_66564_7528# 0.01328f
C27735 a_47164_14136# VPWR 0.29679f
C27736 a_67012_5960# a_67460_5960# 0.01328f
C27737 _231_.ZN vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN 0.00702f
C27738 _442_.ZN a_39324_26247# 0.00957f
C27739 a_39536_26795# a_39772_26247# 0.00984f
C27740 a_31708_18407# a_32068_18504# 0.08717f
C27741 a_932_18504# a_1380_18504# 0.01328f
C27742 _250_.A2 a_63721_28776# 0.00106f
C27743 a_36660_23588# a_36748_23544# 0.28563f
C27744 a_17060_29860# uio_out[7] 0.00288f
C27745 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN 0.14745f
C27746 a_40356_15748# a_40804_15748# 0.01328f
C27747 a_26468_31048# _349_.A4 0.00133f
C27748 a_1828_12232# VPWR 0.20348f
C27749 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN a_63336_29480# 0.01618f
C27750 _330_.A1 _435_.A3 0.00335f
C27751 _251_.A1 _324_.C 2.21575f
C27752 a_14708_24776# VPWR 0.22176f
C27753 a_11460_31048# uio_oe[4] 0.00345f
C27754 a_1468_2727# a_1828_2824# 0.08717f
C27755 _251_.A1 a_64996_31048# 0.04255f
C27756 a_3260_19975# a_3172_20072# 0.28563f
C27757 a_44388_15748# VPWR 0.20703f
C27758 _451_.Q _448_.Q 0.50068f
C27759 a_38472_30169# uo_out[1] 0.04952f
C27760 _424_.A2 a_52652_18407# 0.00747f
C27761 a_44864_27165# a_44571_26841# 0.49319f
C27762 _459_.CLK a_21868_27208# 0.00124f
C27763 a_46180_9476# a_46268_9432# 0.28563f
C27764 a_31372_21976# a_31820_21976# 0.01255f
C27765 _427_.B2 _427_.ZN 0.00363f
C27766 _455_.Q a_24304_26795# 0.01744f
C27767 _399_.A2 a_48308_23588# 0.48718f
C27768 _424_.A2 VPWR 2.39778f
C27769 _294_.A2 a_39300_29480# 0.0019f
C27770 _304_.B a_52764_27815# 0.04459f
C27771 hold2.Z a_42161_24776# 0.02747f
C27772 a_2724_12612# a_2364_12568# 0.08717f
C27773 a_4516_12612# a_4964_12612# 0.01328f
C27774 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I a_66316_20408# 0.02066f
C27775 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN a_62732_26680# 0.00115f
C27776 a_51420_2727# a_51868_2727# 0.0131f
C27777 a_36828_28776# uo_out[7] 0.00106f
C27778 _459_.D VPWR 0.53921f
C27779 _251_.A1 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN 0.00483f
C27780 a_28891_25273# a_29136_25641# 0.00232f
C27781 _447_.Q a_41664_22020# 0.00446f
C27782 a_52228_17316# VPWR 0.20672f
C27783 _370_.ZN a_29788_30345# 0.21711f
C27784 a_64636_1592# VPWR 0.30056f
C27785 a_29232_29931# a_31088_30301# 0.02307f
C27786 a_32828_1159# a_32740_1256# 0.28563f
C27787 a_66428_1592# a_66564_1256# 0.00168f
C27788 a_53212_29816# a_53796_30344# 0.00629f
C27789 _362_.ZN a_30388_28776# 0.01646f
C27790 a_22996_31048# uio_out[4] 0.0063f
C27791 a_62508_12135# a_62420_12232# 0.28563f
C27792 a_21540_1636# a_21180_1592# 0.08707f
C27793 _313_.ZN _312_.ZN 0.26544f
C27794 _229_.I a_61052_27815# 0.00711f
C27795 a_17508_29860# _459_.CLK 0.02271f
C27796 _287_.A1 a_33140_29860# 0.00167f
C27797 a_16948_26344# a_16948_25156# 0.05841f
C27798 a_24988_21543# VPWR 0.31547f
C27799 _457_.D a_26746_26344# 0.02561f
C27800 a_48196_17316# a_48644_17316# 0.01328f
C27801 _319_.ZN a_34396_18840# 0.00123f
C27802 _460_.D a_33164_24679# 0.00176f
C27803 _478_.D a_52920_22760# 0.03939f
C27804 _398_.C a_51988_24072# 0.00142f
C27805 _454_.Q _345_.A2 0.59943f
C27806 a_56484_2824# VPWR 0.20955f
C27807 a_66428_11000# a_66316_10567# 0.02634f
C27808 a_64996_1636# a_65444_1636# 0.01328f
C27809 a_52428_10567# a_52876_10567# 0.01288f
C27810 a_55140_27912# a_55588_27912# 0.01328f
C27811 a_62284_26680# VPWR 0.31389f
C27812 _337_.ZN a_29575_28293# 0.0026f
C27813 a_26556_23111# a_26916_23208# 0.08707f
C27814 a_55588_9476# VPWR 0.20692f
C27815 _230_.I vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN 0.02099f
C27816 a_22660_2824# a_22748_1159# 0.0027f
C27817 a_62756_14180# VPWR 0.20952f
C27818 a_20956_21543# a_21404_21543# 0.01288f
C27819 _231_.ZN a_59652_25640# 0.03616f
C27820 _336_.A2 a_27004_23111# 0.00215f
C27821 _358_.A2 a_31116_26020# 0.00127f
C27822 _452_.CLK a_36544_24419# 0.00167f
C27823 _256_.A2 _246_.B2 0.33262f
C27824 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I a_65756_27815# 0.03496f
C27825 a_41160_29083# a_41440_28363# 0.00267f
C27826 a_63316_12232# VPWR 0.20622f
C27827 a_35740_2727# a_35876_1636# 0.00154f
C27828 a_52228_2824# a_52676_2824# 0.01328f
C27829 _473_.Q a_48921_22020# 0.00337f
C27830 a_6172_30951# a_6308_29860# 0.00154f
C27831 _287_.A1 a_34404_31048# 0.00873f
C27832 a_33524_24776# VPWR 0.21278f
C27833 _452_.Q _438_.ZN 0.72915f
C27834 a_1380_18884# VPWR 0.20348f
C27835 a_12892_2727# a_12804_2824# 0.28563f
C27836 a_50524_15704# VPWR 0.37088f
C27837 _355_.C a_23420_26247# 0.01997f
C27838 a_52639_30644# a_52891_30644# 0.00184f
C27839 _274_.ZN _267_.A2 0.13201f
C27840 a_51420_9432# a_51868_9432# 0.0131f
C27841 a_19076_31048# uio_out[7] 0.00371f
C27842 _258_.I _238_.I 0.17853f
C27843 _325_.A1 a_42252_20936# 0.00155f
C27844 a_64324_15368# a_64300_13703# 0.00131f
C27845 a_932_20452# a_1020_20408# 0.28563f
C27846 _473_.Q a_48172_18840# 0.00252f
C27847 _459_.CLK _373_.ZN 0.76394f
C27848 _319_.A3 a_38304_20072# 0.00908f
C27849 a_52764_27815# VPWR 0.31487f
C27850 _336_.Z a_28012_23544# 0.00234f
C27851 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN 0.01179f
C27852 a_47076_12612# a_46716_12568# 0.08707f
C27853 _274_.ZN a_53212_29816# 0.01181f
C27854 vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I a_63316_20452# 0.00255f
C27855 a_21852_24679# a_21876_23588# 0.0016f
C27856 _312_.ZN _316_.ZN 0.00303f
C27857 _323_.A3 a_38876_19975# 0.00108f
C27858 a_43804_1159# a_44164_1256# 0.08717f
C27859 a_59284_12232# a_59732_12232# 0.01328f
C27860 a_19388_1159# VPWR 0.36593f
C27861 a_24452_1636# a_24540_1592# 0.28563f
C27862 a_28036_1636# a_28484_1636# 0.01328f
C27863 _393_.A1 _404_.A1 0.00842f
C27864 a_22212_21640# VPWR 0.20614f
C27865 _435_.A3 a_39860_25156# 0.00246f
C27866 _350_.A1 a_31484_30951# 0.01205f
C27867 _305_.A2 a_42168_22504# 0.1211f
C27868 a_63292_11000# a_63316_10664# 0.00172f
C27869 a_49740_10567# a_49652_10664# 0.28563f
C27870 _427_.A2 a_53572_21640# 0.00692f
C27871 a_46804_28292# VPWR 0.00667f
C27872 _325_.A2 a_36612_20072# 0.01232f
C27873 a_61076_23208# VPWR 0.19865f
C27874 a_31803_24831# a_32088_24831# 0.00277f
C27875 a_34396_24679# a_34844_24679# 0.01222f
C27876 _304_.B a_42778_21812# 0.03268f
C27877 a_66564_9476# VPWR 0.20959f
C27878 a_58476_20408# VPWR 0.34455f
C27879 _350_.A1 a_29804_30951# 0.01602f
C27880 a_65308_6296# VPWR 0.30378f
C27881 a_19636_23588# VPWR 0.21659f
C27882 _252_.B _243_.ZN 0.04956f
C27883 a_19612_21543# a_19972_21640# 0.08707f
C27884 a_64772_20072# a_65220_20072# 0.01328f
C27885 a_18760_29032# a_19328_28733# 0.00118f
C27886 a_67100_3160# VPWR 0.29679f
C27887 a_49740_13703# VPWR 0.32115f
C27888 _459_.CLK a_22992_27555# 0.01586f
C27889 a_19372_30345# uio_out[7] 0.00224f
C27890 _424_.A2 _424_.B2 0.00274f
C27891 _465_.D _459_.CLK 0.00528f
C27892 a_40004_22020# VPWR 0.00407f
C27893 _459_.CLK a_28124_26680# 0.00715f
C27894 a_50436_15748# a_50524_15704# 0.28563f
C27895 a_46492_15704# a_46940_15704# 0.01288f
C27896 a_52452_11044# VPWR 0.21241f
C27897 a_57168_26724# vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN 0.00157f
C27898 a_48308_23588# a_49316_23588# 0.01836f
C27899 a_59172_26724# a_59260_26680# 0.28563f
C27900 a_9532_29383# uio_oe[5] 0.00106f
C27901 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I VPWR 0.84175f
C27902 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN 0.25032f
C27903 a_3172_26344# VPWR 0.20993f
C27904 a_38644_19368# VPWR 0.00417f
C27905 a_44252_30951# vgaringosc.workerclkbuff_notouch_.I 0.00352f
C27906 a_23868_2727# a_24228_2824# 0.08717f
C27907 a_55228_20408# VPWR 0.32282f
C27908 VPWR uio_in[5] 0.00114f
C27909 _345_.A2 a_23284_26724# 0.00414f
C27910 _355_.C _346_.ZN 0.01091f
C27911 _459_.CLK _369_.ZN 0.00103f
C27912 _409_.ZN _381_.Z 0.02835f
C27913 _473_.Q a_49034_21640# 0.0063f
C27914 _350_.A2 a_30160_30301# 0.00376f
C27915 _324_.C a_58020_27508# 0.00145f
C27916 a_57156_9476# a_57244_9432# 0.28563f
C27917 _287_.A2 a_30388_28776# 0.02118f
C27918 a_4516_28292# VPWR 0.20812f
C27919 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I a_58836_18884# 0.00141f
C27920 a_45416_29885# a_44795_29535# 0.00705f
C27921 a_39884_27815# a_39796_27912# 0.28563f
C27922 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN a_54692_15748# 0.00135f
C27923 a_65892_14180# a_65980_14136# 0.28563f
C27924 a_14796_20408# a_15244_20408# 0.0131f
C27925 a_16948_20452# a_16588_20408# 0.08717f
C27926 a_19164_30951# uio_out[7] 0.00257f
C27927 _267_.A1 _267_.ZN 0.37871f
C27928 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 1.07398f
C27929 a_61860_30736# a_62532_30736# 0.00219f
C27930 a_1380_1636# VPWR 0.20348f
C27931 _397_.A2 a_49212_26369# 0.00708f
C27932 _416_.A1 _284_.B 0.73468f
C27933 _251_.A1 _252_.ZN 0.45434f
C27934 a_53572_12612# a_54020_12612# 0.01328f
C27935 a_36748_23544# a_36860_23111# 0.02634f
C27936 a_22560_30288# a_23196_29816# 0.0057f
C27937 a_41788_1159# VPWR 0.33478f
C27938 _267_.A1 _390_.ZN 0.01118f
C27939 a_55228_1159# a_55140_1256# 0.28563f
C27940 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I 0.64644f
C27941 _467_.D a_16796_27209# 0.21478f
C27942 _304_.A1 _311_.Z 0.53033f
C27943 _229_.I a_61412_27912# 0.00546f
C27944 a_55812_1636# a_55676_1159# 0.00168f
C27945 a_15132_1159# a_15580_1159# 0.0131f
C27946 a_60268_10567# a_60628_10664# 0.08707f
C27947 a_46180_10664# a_46628_10664# 0.01328f
C27948 a_37968_31048# uo_out[3] 0.00254f
C27949 a_16612_2824# a_16612_1636# 0.05841f
C27950 a_54356_23588# a_54804_23588# 0.01328f
C27951 a_20532_22020# VPWR 0.20622f
C27952 _424_.A2 a_51240_23340# 0.07467f
C27953 a_42778_21812# VPWR 0.61363f
C27954 _390_.ZN _408_.ZN 0.02522f
C27955 a_27116_23544# VPWR 0.36266f
C27956 a_56572_23111# VPWR 0.31699f
C27957 a_3620_13800# VPWR 0.22347f
C27958 a_47860_21640# _416_.A2 0.0889f
C27959 a_30588_21543# a_30500_21640# 0.28563f
C27960 a_21852_2727# VPWR 0.31143f
C27961 a_17844_21640# a_18628_21640# 0.00276f
C27962 a_58388_20452# a_58028_20408# 0.08674f
C27963 a_61724_15271# a_62172_15271# 0.0131f
C27964 a_8996_31048# uio_oe[6] 0.00329f
C27965 a_6756_29860# VPWR 0.20648f
C27966 a_53660_21543# a_53796_20452# 0.00154f
C27967 a_67012_15748# a_66876_15271# 0.00168f
C27968 a_58588_11000# VPWR 0.32371f
C27969 a_41116_26247# a_41028_26344# 0.28563f
C27970 _287_.A1 _362_.B 0.03041f
C27971 a_59172_22020# vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.00278f
C27972 _355_.C _459_.CLK 2.47416f
C27973 _267_.A1 a_55228_28248# 0.0054f
C27974 a_65308_15704# a_65756_15704# 0.01255f
C27975 _325_.A1 a_42154_21236# 0.01722f
C27976 a_932_27912# VPWR 0.22176f
C27977 _437_.A1 a_37980_26247# 0.04814f
C27978 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I 0.03595f
C27979 _373_.ZN uo_out[7] 0.00142f
C27980 a_62508_23111# a_62420_23208# 0.28563f
C27981 _424_.A2 a_44744_26355# 0.00179f
C27982 a_35292_2727# a_35204_2824# 0.28563f
C27983 _371_.A3 a_28124_26680# 0.00195f
C27984 a_62396_9432# a_62844_9432# 0.0131f
C27985 a_15604_23588# a_16052_23588# 0.01328f
C27986 _407_.A1 _407_.ZN 0.35752f
C27987 a_64324_7908# a_64772_7908# 0.01328f
C27988 a_16164_1256# a_16612_1256# 0.01328f
C27989 a_65220_6340# a_65668_6340# 0.01328f
C27990 a_64324_4772# a_64412_4728# 0.28563f
C27991 a_66116_4772# a_66564_4772# 0.01328f
C27992 a_65220_3204# a_65308_3160# 0.28563f
C27993 a_67012_3204# a_67460_3204# 0.01328f
C27994 _251_.A1 a_61500_26247# 0.00628f
C27995 a_45372_13703# a_45820_13703# 0.0131f
C27996 hold2.I hold1.Z 0.1921f
C27997 a_58364_25112# vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN 0.0024f
C27998 a_8627_30644# a_7540_31048# 0.00182f
C27999 a_7628_30951# a_8996_31048# 0.00266f
C28000 a_6620_29383# a_7068_29383# 0.0131f
C28001 a_47776_20893# a_47552_19715# 0.0015f
C28002 _452_.CLK _443_.D 0.08297f
C28003 a_15044_1636# VPWR 0.20348f
C28004 _459_.CLK a_24636_25641# 0.00171f
C28005 _369_.ZN _371_.A3 0.42255f
C28006 a_60292_12612# a_60964_12612# 0.00347f
C28007 a_63316_13800# a_63404_12135# 0.00151f
C28008 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN 0.78579f
C28009 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62503_28293# 0.02098f
C28010 _336_.A1 a_28596_26725# 0.03274f
C28011 a_59260_23111# a_59620_23208# 0.08674f
C28012 _359_.B a_28928_29123# 0.05667f
C28013 _330_.ZN a_37868_16839# 0.00667f
C28014 a_66204_1159# a_66564_1256# 0.0869f
C28015 a_1380_5960# VPWR 0.20348f
C28016 a_3708_19975# VPWR 0.33374f
C28017 a_64188_1159# VPWR 0.2977f
C28018 _435_.A3 a_38616_24328# 0.00497f
C28019 a_36188_25112# a_36636_25112# 0.01255f
C28020 a_31620_16936# a_32068_16936# 0.01328f
C28021 a_38116_1636# a_38204_1592# 0.28563f
C28022 a_34172_1592# a_34620_1592# 0.01288f
C28023 a_2364_1592# a_2364_1159# 0.05841f
C28024 a_6308_1636# a_6172_1159# 0.00168f
C28025 a_48420_11044# a_48868_11044# 0.01328f
C28026 a_5388_18407# VPWR 0.35526f
C28027 a_23780_26344# VPWR 0.20674f
C28028 _325_.A2 a_44276_17316# 0.08637f
C28029 a_44948_28292# VPWR 0.14344f
C28030 _255_.ZN _238_.I 0.00227f
C28031 _459_.CLK a_27908_27912# 0.00135f
C28032 _274_.A1 a_55588_28292# 0.03795f
C28033 _436_.B _438_.ZN 0.00155f
C28034 a_40580_26344# _433_.ZN 0.00166f
C28035 _397_.A2 _411_.A2 0.52839f
C28036 a_26668_21976# VPWR 0.32418f
C28037 _390_.ZN _412_.A1 0.12786f
C28038 _324_.C _421_.A1 0.02778f
C28039 _452_.CLK a_33724_23111# 0.00815f
C28040 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I 0.68102f
C28041 a_42908_30951# a_43356_30951# 0.0131f
C28042 a_35504_18955# a_36432_19325# 1.16391f
C28043 a_44252_2727# VPWR 0.31143f
C28044 a_65332_13800# VPWR 0.21224f
C28045 a_40264_30320# VPWR 0.47878f
C28046 a_18716_26247# a_19164_26247# 0.01222f
C28047 a_4156_26247# a_4852_26344# 0.01227f
C28048 a_57244_27815# _242_.Z 0.00217f
C28049 a_12892_29816# VPWR 0.29679f
C28050 a_58911_30644# ui_in[2] 0.00123f
C28051 a_63988_16936# a_63964_15704# 0.0016f
C28052 a_45372_10567# VPWR 0.30073f
C28053 _272_.A2 a_56596_29861# 0.15334f
C28054 _369_.ZN uo_out[7] 0.01158f
C28055 a_32156_15271# a_32516_15368# 0.08717f
C28056 a_31484_23111# VPWR 0.31572f
C28057 _379_.A2 a_20672_30301# 0.08558f
C28058 a_61836_23544# a_61972_23208# 0.00168f
C28059 _324_.B a_44948_22020# 0.03038f
C28060 _474_.D a_49896_18909# 0.3019f
C28061 a_46624_19715# a_47259_20127# 0.02112f
C28062 _258_.I VPWR 0.97398f
C28063 _424_.B2 a_52136_20936# 0.00757f
C28064 a_46044_2727# a_46628_2824# 0.01675f
C28065 a_48508_30951# uio_in[1] 0.00118f
C28066 a_62532_17316# a_62620_17272# 0.28563f
C28067 a_52852_24372# _427_.A2 0.00101f
C28068 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I 0.01926f
C28069 a_932_16936# a_932_15748# 0.05841f
C28070 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN VPWR 0.71673f
C28071 a_65756_9432# a_65756_8999# 0.05841f
C28072 a_59260_26680# a_59397_26344# 0.00109f
C28073 a_66540_18407# a_66988_18407# 0.01255f
C28074 _474_.CLK a_55140_20452# 0.04193f
C28075 _304_.B hold1.Z 0.61923f
C28076 _223_.I a_31088_30301# 0.19672f
C28077 a_33060_31048# VPWR 0.01457f
C28078 a_2812_13703# a_2724_13800# 0.28563f
C28079 a_27924_20452# a_27564_20408# 0.08717f
C28080 a_63876_18504# a_63876_17316# 0.05841f
C28081 _416_.A1 a_45088_29123# 0.01589f
C28082 _457_.D a_25348_24776# 0.00467f
C28083 a_54432_31128# input9.Z 0.05393f
C28084 a_4156_16839# a_4068_16936# 0.28563f
C28085 a_36412_1592# a_36548_1256# 0.00168f
C28086 _419_.Z a_47483_20569# 0.01058f
C28087 a_21180_1592# VPWR 0.3289f
C28088 a_67236_12612# a_67684_12612# 0.01328f
C28089 _427_.B1 a_53460_24776# 0.01111f
C28090 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN 0.63963f
C28091 a_64100_12612# a_63740_12568# 0.08707f
C28092 _390_.ZN a_51968_26724# 0.02369f
C28093 _276_.A2 uio_in[0] 0.02098f
C28094 a_66876_15271# a_67236_15368# 0.08674f
C28095 _304_.A1 a_39780_22805# 0.00148f
C28096 a_64212_12232# a_64188_11000# 0.0016f
C28097 a_41476_1636# a_41116_1592# 0.08707f
C28098 _264_.B a_40468_25157# 0.12726f
C28099 a_50548_12232# a_50636_10567# 0.00151f
C28100 _260_.A1 _324_.B 0.17596f
C28101 a_4964_26724# a_5052_26680# 0.28563f
C28102 _245_.I1 a_62796_25640# 0.00157f
C28103 _242_.Z a_58500_26344# 0.0026f
C28104 a_22100_29480# VPWR 0.2094f
C28105 a_37532_1159# a_37980_1159# 0.0131f
C28106 _324_.B a_47047_21640# 0.00108f
C28107 _397_.A2 _399_.ZN 0.02145f
C28108 _336_.A2 a_28012_24679# 0.01777f
C28109 a_2364_20408# VPWR 0.30029f
C28110 a_66652_2727# VPWR 0.29679f
C28111 a_67460_2824# a_67548_1159# 0.0027f
C28112 _452_.CLK a_31396_23208# 0.00187f
C28113 a_46716_12568# VPWR 0.29679f
C28114 a_62196_16936# a_62644_16936# 0.01328f
C28115 _452_.Q a_40692_21640# 0.00519f
C28116 a_41476_26344# _451_.Q 0.00259f
C28117 a_5276_29383# a_5188_29480# 0.28563f
C28118 a_35716_20072# VPWR 0.00673f
C28119 a_41476_15368# a_42148_15368# 0.00347f
C28120 _371_.A3 a_27908_27912# 0.02028f
C28121 a_67212_10567# VPWR 0.31389f
C28122 a_61076_20452# vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I 0.07122f
C28123 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN a_61164_20408# 0.00678f
C28124 a_64324_29860# vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I 0.11153f
C28125 _274_.A1 a_53412_29480# 0.00307f
C28126 a_43580_15271# a_43492_15368# 0.28563f
C28127 a_29156_23208# VPWR 0.20595f
C28128 _430_.ZN _441_.A3 0.02314f
C28129 a_44924_15271# a_45372_15271# 0.0131f
C28130 _304_.B _478_.D 0.01281f
C28131 _247_.B a_60156_27815# 0.0303f
C28132 a_54892_19975# a_55340_19975# 0.012f
C28133 a_15156_28292# a_14796_28248# 0.0869f
C28134 _272_.B1 _255_.ZN 0.13658f
C28135 _448_.Q _319_.A2 0.06307f
C28136 a_57468_2727# a_57380_2824# 0.28563f
C28137 a_16500_22020# a_16948_22020# 0.01328f
C28138 _336_.A2 a_29184_25597# 0.00773f
C28139 a_40668_19975# _450_.D 0.00818f
C28140 a_1468_16839# a_1916_16839# 0.0131f
C28141 a_13364_31048# uio_oe[2] 0.00726f
C28142 a_56236_23544# clk 0.00613f
C28143 a_64772_15748# VPWR 0.20973f
C28144 _459_.Q a_31284_23588# 0.002f
C28145 _358_.A3 a_36100_26724# 0.00241f
C28146 a_32848_29123# uo_out[6] 0.02912f
C28147 a_59260_21976# VPWR 0.32419f
C28148 a_34644_16936# a_34756_15748# 0.02666f
C28149 _332_.Z a_40644_17272# 0.00238f
C28150 _409_.ZN _324_.C 0.19871f
C28151 hold1.Z VPWR 0.6628f
C28152 a_23108_23208# a_23196_21543# 0.00151f
C28153 a_3172_7908# VPWR 0.20993f
C28154 a_23084_23544# a_23532_23544# 0.0131f
C28155 a_38340_1256# a_39012_1256# 0.00347f
C28156 a_26580_23588# a_26220_23544# 0.0869f
C28157 a_8996_1256# VPWR 0.20348f
C28158 a_12916_31048# VPWR 0.20809f
C28159 a_21428_25156# a_21068_25112# 0.08707f
C28160 a_4964_4772# VPWR 0.21167f
C28161 a_67212_13703# a_67660_13703# 0.0131f
C28162 a_17596_2727# a_18044_2727# 0.0131f
C28163 _251_.A1 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN 0.02792f
C28164 a_53324_13703# a_53684_13800# 0.08707f
C28165 _369_.ZN a_30128_27508# 0.00101f
C28166 _424_.A2 a_52434_22504# 0.00571f
C28167 a_40580_26344# _261_.ZN 0.00329f
C28168 a_1020_17272# a_1020_16839# 0.05841f
C28169 a_40108_16839# a_40468_16936# 0.08707f
C28170 a_54356_25156# a_53996_25112# 0.0869f
C28171 _251_.A1 a_60964_26344# 0.00569f
C28172 _311_.A2 a_36300_23544# 0.01311f
C28173 a_47076_10664# a_47076_9476# 0.05841f
C28174 a_66988_16839# VPWR 0.31389f
C28175 a_34980_1636# VPWR 0.24722f
C28176 a_4516_1636# a_4156_1592# 0.08707f
C28177 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN _250_.C 0.006f
C28178 a_2724_29860# a_3172_29860# 0.01328f
C28179 a_45012_29816# a_45800_30345# 0.02112f
C28180 a_45416_29885# a_45904_30180# 0.8399f
C28181 a_49988_21236# VPWR 0.8484f
C28182 a_2724_17316# a_2364_17272# 0.08717f
C28183 a_4516_17316# a_4964_17316# 0.01328f
C28184 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN clk 0.00914f
C28185 a_54556_11000# a_55004_11000# 0.01288f
C28186 _352_.A2 a_24080_25227# 0.04958f
C28187 a_58500_11044# a_58588_11000# 0.28563f
C28188 a_47972_1636# a_48420_1636# 0.01328f
C28189 a_53460_16936# a_53908_16936# 0.01328f
C28190 a_45396_25156# VPWR 0.02076f
C28191 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN a_61412_17316# 0.07117f
C28192 a_1828_20072# a_1828_18884# 0.05841f
C28193 a_57940_17316# a_57580_17272# 0.0869f
C28194 a_19948_26680# _455_.D 0.00296f
C28195 a_20396_26680# a_20844_26680# 0.012f
C28196 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I 0.00128f
C28197 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN a_57380_16936# 0.00902f
C28198 _330_.A1 _411_.A2 0.04151f
C28199 a_54244_18884# VPWR 0.22779f
C28200 _359_.ZN VPWR 0.40941f
C28201 a_2724_25156# VPWR 0.20782f
C28202 a_62532_18884# a_62172_18840# 0.08717f
C28203 a_62148_29505# VPWR 0.01105f
C28204 a_1916_27815# a_2276_27912# 0.08717f
C28205 a_16140_27815# a_16588_27815# 0.0131f
C28206 a_22412_20408# VPWR 0.31605f
C28207 a_35740_25112# _444_.D 0.00449f
C28208 a_3620_15748# a_3708_15704# 0.28563f
C28209 a_60380_12568# VPWR 0.34385f
C28210 _417_.A2 _475_.Q 0.1714f
C28211 a_18404_2824# a_18852_2824# 0.01328f
C28212 a_16252_29383# a_16612_29480# 0.08674f
C28213 _399_.ZN a_48308_23588# 0.05112f
C28214 _371_.ZN a_26720_30301# 0.00257f
C28215 _395_.A1 _281_.ZN 0.0512f
C28216 a_61076_10664# VPWR 0.20641f
C28217 a_4940_8999# a_4852_9096# 0.28563f
C28218 a_64412_7431# a_64324_7528# 0.28563f
C28219 a_54556_15271# a_54916_15368# 0.08717f
C28220 a_65308_5863# a_65220_5960# 0.28563f
C28221 a_66204_4295# a_66116_4392# 0.28563f
C28222 _474_.Q a_49896_18909# 0.00893f
C28223 a_34532_15368# VPWR 0.23243f
C28224 _478_.D VPWR 0.35929f
C28225 _249_.A2 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN 0.00928f
C28226 _284_.A2 a_49952_26724# 0.00126f
C28227 _304_.B a_47376_27912# 0.01247f
C28228 a_37756_15271# VPWR 0.3577f
C28229 a_21740_29383# _378_.I 0.00717f
C28230 a_4516_14180# a_4964_14180# 0.01328f
C28231 a_2724_14180# a_2364_14136# 0.08717f
C28232 a_33768_29535# VPWR 0.0022f
C28233 a_62172_17272# VPWR 0.3185f
C28234 a_14908_30951# uio_oe[2] 0.00333f
C28235 a_31396_1256# VPWR 0.22423f
C28236 a_66204_7431# VPWR 0.31657f
C28237 a_932_4392# VPWR 0.22176f
C28238 a_62308_26344# VPWR 0.20566f
C28239 a_64300_13703# a_64212_13800# 0.28563f
C28240 _284_.A2 _384_.A3 0.02023f
C28241 a_14460_30951# VPWR 0.31184f
C28242 a_33052_17272# a_33052_16839# 0.05841f
C28243 a_36996_17316# a_36972_16839# 0.00172f
C28244 a_51308_16839# a_51220_16936# 0.28563f
C28245 a_40196_31048# VPWR 0.01455f
C28246 a_3172_23208# a_3172_22020# 0.05841f
C28247 a_64772_18504# VPWR 0.20727f
C28248 a_9980_1159# a_10340_1256# 0.08717f
C28249 a_54220_12135# a_54668_12135# 0.01288f
C28250 _251_.A1 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN 0.01061f
C28251 a_41116_1592# VPWR 0.33204f
C28252 a_24316_26247# _457_.D 0.00299f
C28253 a_46516_16936# VPWR 0.20703f
C28254 a_25324_23544# a_25436_23111# 0.02634f
C28255 a_48104_30219# _392_.A2 0.00556f
C28256 a_3172_29480# a_3620_29480# 0.01328f
C28257 _452_.CLK a_36636_26680# 0.04136f
C28258 a_11012_1636# a_11460_1636# 0.01328f
C28259 hold2.I clkbuf_1_0__f_clk.I 0.08575f
C28260 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I a_57492_18884# 0.0082f
C28261 _325_.A1 a_43664_17317# 0.10741f
C28262 a_32516_17316# a_32156_17272# 0.08707f
C28263 a_21740_30951# uio_out[4] 0.00619f
C28264 a_52092_11000# a_51980_10567# 0.02634f
C28265 _436_.B a_40132_26344# 0.00554f
C28266 a_61860_11044# a_61948_11000# 0.28563f
C28267 a_11236_2824# VPWR 0.21654f
C28268 _255_.ZN VPWR 1.06482f
C28269 a_55140_1636# a_54780_1592# 0.08663f
C28270 _393_.A3 a_48596_28292# 0.00426f
C28271 _474_.CLK _400_.ZN 0.07145f
C28272 _359_.B a_35204_26344# 0.05046f
C28273 _459_.CLK a_16500_26344# 0.00641f
C28274 _416_.A2 a_47483_20569# 0.049f
C28275 a_16588_24679# a_17036_24679# 0.0131f
C28276 a_59932_1159# a_60380_1159# 0.0131f
C28277 a_67212_20408# a_68020_20452# 0.00965f
C28278 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN a_54356_18504# 0.00876f
C28279 a_54892_18407# a_54804_18504# 0.28563f
C28280 a_64996_15368# VPWR 0.22891f
C28281 a_21068_25112# VPWR 0.31547f
C28282 a_1020_18407# a_1468_18407# 0.0131f
C28283 _427_.ZN a_54692_20452# 0.00422f
C28284 a_33412_15748# a_33500_15704# 0.28563f
C28285 a_47164_12135# VPWR 0.29679f
C28286 _340_.A2 _373_.ZN 0.00594f
C28287 a_36996_15748# a_37444_15748# 0.01328f
C28288 a_21404_2727# a_21540_1636# 0.00154f
C28289 _260_.A2 _324_.B 0.18917f
C28290 a_50772_18504# a_50884_17316# 0.02666f
C28291 a_47076_18504# a_46940_17272# 0.00154f
C28292 _397_.A1 a_50792_26344# 0.02759f
C28293 _301_.A1 VPWR 1.69251f
C28294 a_44160_29123# a_44795_29535# 0.02112f
C28295 a_61412_26344# vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN 0.00164f
C28296 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN a_59260_23544# 0.00382f
C28297 a_62864_25156# VPWR 0.00645f
C28298 a_39236_20072# VPWR 0.20753f
C28299 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN a_55228_15704# 0.00189f
C28300 _452_.CLK a_43916_16839# 0.00239f
C28301 a_5052_15704# VPWR 0.33516f
C28302 a_56708_15368# VPWR 0.21257f
C28303 _260_.ZN a_42778_21812# 0.01274f
C28304 a_44459_18559# a_44752_18147# 0.49319f
C28305 _424_.B1 _279_.Z 0.01375f
C28306 a_55700_24776# clk 0.01113f
C28307 a_22636_21976# a_23084_21976# 0.01288f
C28308 a_26580_22020# a_26668_21976# 0.28563f
C28309 _330_.A1 _430_.ZN 0.41112f
C28310 a_47376_27912# VPWR 0.01379f
C28311 a_47076_14180# a_46716_14136# 0.08707f
C28312 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN a_54804_16936# 0.00615f
C28313 a_48396_16839# a_48844_16839# 0.01288f
C28314 _304_.B a_46198_27060# 0.00228f
C28315 a_41452_16839# VPWR 0.30108f
C28316 a_53572_1256# VPWR 0.20968f
C28317 a_37644_23544# _439_.ZN 0.01615f
C28318 a_60740_1256# a_61188_1256# 0.01328f
C28319 _435_.A3 _264_.B 0.1424f
C28320 a_58836_17316# VPWR 0.20981f
C28321 a_61076_13800# a_61524_13800# 0.01328f
C28322 a_50176_26724# _381_.A2 0.00109f
C28323 a_39996_2727# a_40444_2727# 0.0131f
C28324 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I VPWR 0.74623f
C28325 _474_.CLK a_54892_25112# 0.02247f
C28326 _421_.A1 a_47271_21640# 0.09058f
C28327 _284_.ZN uo_out[0] 1.50447f
C28328 _346_.B _346_.A2 0.0101f
C28329 a_20868_23208# a_20980_22020# 0.02666f
C28330 a_32156_17272# VPWR 0.29679f
C28331 a_4852_10664# a_4940_8999# 0.00151f
C28332 _416_.A2 a_46624_19715# 0.01138f
C28333 a_54780_1592# VPWR 0.29679f
C28334 a_21404_1159# a_21316_1256# 0.28563f
C28335 _304_.B clkbuf_1_0__f_clk.I 0.02986f
C28336 a_51532_12135# a_51444_12232# 0.28563f
C28337 _402_.A1 a_44340_26183# 0.00541f
C28338 a_8860_29816# a_9308_29816# 0.01288f
C28339 a_12804_29860# a_12892_29816# 0.28563f
C28340 a_40040_17675# a_39324_17272# 0.00367f
C28341 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN 0.04219f
C28342 _317_.A2 a_37532_21543# 0.00235f
C28343 _336_.A2 a_28372_23588# 0.00292f
C28344 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN 0.65475f
C28345 _336_.A1 a_27476_23588# 0.00173f
C28346 a_1468_10567# a_1916_10567# 0.0131f
C28347 a_59036_11000# a_58924_10567# 0.02634f
C28348 a_58052_1636# a_58140_1592# 0.28563f
C28349 a_61636_1636# a_62084_1636# 0.01328f
C28350 a_33636_2824# VPWR 0.20713f
C28351 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I 0.0012f
C28352 _424_.B1 a_50704_27912# 0.00367f
C28353 a_15244_23111# a_15604_23208# 0.08717f
C28354 a_27452_23111# a_27900_23111# 0.01288f
C28355 a_19164_24679# a_19524_24776# 0.08707f
C28356 _402_.ZN _417_.A2 0.00223f
C28357 _444_.D a_37196_23544# 0.00277f
C28358 a_1020_9432# VPWR 0.30073f
C28359 a_51780_2824# a_51644_1592# 0.00154f
C28360 a_11236_2824# a_11324_1159# 0.0027f
C28361 a_46716_14136# VPWR 0.29679f
C28362 _397_.A1 _281_.ZN 0.33459f
C28363 a_31708_18407# a_31620_18504# 0.28563f
C28364 _250_.A2 a_63313_28776# 0.00102f
C28365 a_36660_23588# a_36300_23544# 0.0869f
C28366 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN 0.05473f
C28367 a_16612_29860# uio_out[7] 0.00178f
C28368 a_4068_31048# a_4068_29860# 0.05841f
C28369 a_1380_12232# VPWR 0.20348f
C28370 a_54088_22895# a_54040_22366# 0.00173f
C28371 a_49628_15704# a_49764_15368# 0.00168f
C28372 a_40804_2824# a_41252_2824# 0.01328f
C28373 a_54468_21640# a_54444_19975# 0.00131f
C28374 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN 0.01477f
C28375 _304_.B a_42252_20936# 0.21519f
C28376 _355_.C a_31820_25112# 0.00136f
C28377 _375_.Z uio_out[5] 0.00584f
C28378 a_5300_24776# VPWR 0.21406f
C28379 a_10452_31048# uio_oe[4] 0.00409f
C28380 a_29156_21640# a_29268_20452# 0.02666f
C28381 a_1468_2727# a_1380_2824# 0.28563f
C28382 _350_.A2 _352_.A2 2.09747f
C28383 a_43940_15748# VPWR 0.20692f
C28384 a_2812_19975# a_3172_20072# 0.08717f
C28385 a_43008_26795# a_43888_27209# 0.00306f
C28386 _301_.A1 a_40452_22504# 0.00167f
C28387 a_46180_9476# a_45820_9432# 0.08717f
C28388 a_47524_9476# a_47972_9476# 0.01328f
C28389 _455_.Q a_21600_26725# 0.10815f
C28390 _334_.A1 a_37516_27599# 0.00547f
C28391 a_46198_27060# VPWR 0.67733f
C28392 _459_.CLK uio_out[3] 0.03153f
C28393 a_53572_14180# a_54020_14180# 0.01328f
C28394 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN a_57828_25156# 0.02061f
C28395 _267_.A2 a_53592_30344# 0.00127f
C28396 _304_.B a_52316_27815# 0.03198f
C28397 a_31732_25156# VPWR 0.19114f
C28398 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I a_67124_20452# 0.00177f
C28399 a_2276_12612# a_2364_12568# 0.28563f
C28400 a_52204_18407# a_52228_17316# 0.0016f
C28401 a_36420_28776# uo_out[7] 0.00106f
C28402 a_34304_24029# a_34939_23705# 0.02112f
C28403 _447_.Q a_41460_22020# 0.00135f
C28404 a_24004_23208# a_23980_21976# 0.0016f
C28405 _370_.ZN a_30160_30301# 0.0072f
C28406 a_51780_17316# VPWR 0.20651f
C28407 a_29232_29931# a_29788_30345# 0.8399f
C28408 a_27812_23208# a_27924_22020# 0.02666f
C28409 a_32380_1159# a_32740_1256# 0.08717f
C28410 clkbuf_1_0__f_clk.I VPWR 5.83508f
C28411 a_53212_29816# a_53592_30344# 0.00736f
C28412 a_64188_1592# VPWR 0.2977f
C28413 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I clk 0.009f
C28414 a_47972_12232# a_48420_12232# 0.01328f
C28415 a_59484_12568# a_59396_11044# 0.00151f
C28416 a_62060_12135# a_62420_12232# 0.08707f
C28417 _294_.ZN _337_.ZN 0.00343f
C28418 a_22548_31048# uio_out[4] 0.01302f
C28419 a_21092_1636# a_21180_1592# 0.28563f
C28420 a_17148_1592# a_17596_1592# 0.01288f
C28421 _243_.B2 _243_.ZN 0.09222f
C28422 _242_.Z a_58656_27912# 0.0036f
C28423 _313_.ZN a_33636_23208# 0.00586f
C28424 _287_.A1 a_32916_29860# 0.00991f
C28425 _296_.ZN _288_.ZN 0.00291f
C28426 _229_.I a_60604_27815# 0.00553f
C28427 _379_.A2 a_19140_29612# 0.00647f
C28428 a_24540_21543# VPWR 0.31547f
C28429 a_17060_29860# _459_.CLK 0.0156f
C28430 _355_.C _340_.A2 0.04336f
C28431 a_49092_15368# a_49292_13703# 0.00119f
C28432 a_55900_11000# a_55924_10664# 0.00172f
C28433 a_23084_28248# _345_.A2 0.02082f
C28434 a_56036_2824# VPWR 0.20815f
C28435 _324_.C _305_.A2 0.00168f
C28436 a_41476_1636# a_41340_1159# 0.00168f
C28437 _284_.ZN hold2.Z 0.05548f
C28438 a_2276_2824# a_2276_1636# 0.05841f
C28439 _246_.B2 _238_.ZN 0.00386f
C28440 _350_.A1 uo_out[4] 0.09864f
C28441 _400_.ZN _398_.C 0.00122f
C28442 a_61836_26680# VPWR 0.32058f
C28443 a_26556_23111# a_26468_23208# 0.28563f
C28444 a_21316_24776# a_21764_24776# 0.01328f
C28445 a_41476_24776# _304_.A1 0.01277f
C28446 a_55140_9476# VPWR 0.20692f
C28447 _355_.C _459_.Q 0.10856f
C28448 a_62308_14180# VPWR 0.20952f
C28449 a_37408_18504# _330_.ZN 0.28969f
C28450 _441_.ZN a_39781_24372# 0.00543f
C28451 _452_.CLK a_35616_24776# 0.0183f
C28452 _433_.ZN _438_.ZN 0.09346f
C28453 a_12916_31048# a_12804_29860# 0.02666f
C28454 _462_.D _459_.CLK 0.01199f
C28455 a_62868_12232# VPWR 0.20622f
C28456 _258_.ZN ui_in[4] 0.00132f
C28457 a_43132_15704# a_43580_15704# 0.01288f
C28458 a_42252_20936# VPWR 0.01013f
C28459 _416_.A1 _444_.D 0.54235f
C28460 a_62172_18840# a_62172_18407# 0.05841f
C28461 a_66564_18884# a_66540_18407# 0.00172f
C28462 a_33076_24776# VPWR 0.13249f
C28463 a_932_18884# VPWR 0.22176f
C28464 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN 0.42606f
C28465 a_30476_25112# a_30240_24776# 0.00984f
C28466 a_12444_2727# a_12804_2824# 0.08717f
C28467 _255_.I _324_.C 0.24944f
C28468 a_50076_15704# VPWR 0.33936f
C28469 _350_.A2 a_30912_27508# 0.00394f
C28470 a_64412_19975# a_64860_19975# 0.01222f
C28471 _243_.ZN a_59172_26724# 0.03529f
C28472 _355_.C a_22352_25987# 0.05571f
C28473 _301_.A1 a_36636_21543# 0.00344f
C28474 _325_.A1 a_40668_20408# 0.00191f
C28475 a_18628_31048# uio_out[7] 0.01212f
C28476 a_47388_17272# a_47300_15748# 0.00151f
C28477 a_23084_25112# a_22996_23588# 0.00151f
C28478 a_2724_20452# a_3172_20452# 0.01328f
C28479 _459_.CLK a_25962_29480# 0.00269f
C28480 a_52316_27815# VPWR 0.32775f
C28481 _336_.Z a_27564_23544# 0.00118f
C28482 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I 0.00271f
C28483 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN 0.01067f
C28484 _324_.B a_44276_20072# 0.01227f
C28485 _243_.B2 a_58140_26680# 0.03466f
C28486 a_46628_12612# a_46716_12568# 0.28563f
C28487 a_62396_2727# a_62844_2727# 0.0131f
C28488 a_50212_12612# a_50660_12612# 0.01328f
C28489 _312_.ZN a_33152_22091# 0.00341f
C28490 a_33636_23208# _316_.ZN 0.0046f
C28491 _268_.A1 _275_.ZN 0.0015f
C28492 _276_.A2 _274_.ZN 0.46354f
C28493 _370_.B a_32308_29167# 0.00129f
C28494 a_67548_18840# a_67460_17316# 0.00151f
C28495 a_18940_1159# VPWR 0.30585f
C28496 a_31172_20072# a_31620_20072# 0.01328f
C28497 a_43804_1159# a_43716_1256# 0.28563f
C28498 _323_.A3 a_37384_19624# 0.03686f
C28499 a_64772_9096# a_64772_7908# 0.05841f
C28500 a_23868_1592# a_24540_1592# 0.00544f
C28501 a_65668_7528# a_65668_6340# 0.05841f
C28502 a_62844_12568# a_62756_11044# 0.00151f
C28503 a_66564_5960# a_66564_4772# 0.05841f
C28504 _390_.ZN _381_.Z 0.03759f
C28505 a_49764_26724# clkload0.Z 0.01045f
C28506 a_67460_4392# a_67460_3204# 0.05841f
C28507 a_21764_21640# VPWR 0.20641f
C28508 a_36188_26247# a_36636_26247# 0.01255f
C28509 a_50972_17272# a_51420_17272# 0.01288f
C28510 _397_.A2 _330_.A1 0.0312f
C28511 a_62956_10567# a_63404_10567# 0.01288f
C28512 _452_.CLK a_40580_26344# 0.00546f
C28513 a_49292_10567# a_49652_10664# 0.08707f
C28514 a_3708_1159# a_4156_1159# 0.0131f
C28515 _260_.ZN hold1.Z 0.94357f
C28516 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN a_65668_27912# 0.00617f
C28517 a_46580_28292# VPWR 0.01385f
C28518 a_24900_23208# a_25348_23208# 0.01328f
C28519 a_59620_23208# VPWR 0.21096f
C28520 _304_.B a_42154_21236# 0.01923f
C28521 a_66116_9476# VPWR 0.24066f
C28522 a_31484_21543# a_31932_21543# 0.01288f
C28523 a_58028_20408# VPWR 0.35366f
C28524 a_64860_6296# VPWR 0.30145f
C28525 a_19188_23588# VPWR 0.22891f
C28526 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I VPWR 0.76632f
C28527 a_19612_21543# a_19524_21640# 0.28563f
C28528 a_66652_3160# VPWR 0.29679f
C28529 a_19744_30301# uio_out[7] 0.0017f
C28530 a_67460_2824# a_67324_1592# 0.00154f
C28531 a_5188_29480# a_5052_28248# 0.00154f
C28532 a_49292_13703# VPWR 0.32411f
C28533 _470_.Q _403_.ZN 0.00735f
C28534 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN 0.63788f
C28535 _395_.A2 a_51332_24372# 0.00546f
C28536 _427_.ZN a_52452_21236# 0.44225f
C28537 a_27140_26724# a_27588_26724# 0.01328f
C28538 _459_.CLK a_27676_26680# 0.01765f
C28539 a_52004_11044# VPWR 0.20622f
C28540 a_37296_22020# VPWR 0.01421f
C28541 a_50436_15748# a_50076_15704# 0.08707f
C28542 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN 0.1729f
C28543 a_13340_29816# a_13340_29383# 0.05841f
C28544 a_35108_28776# VPWR 0.00228f
C28545 a_63204_2824# a_63652_2824# 0.01328f
C28546 a_62756_27912# a_62732_26680# 0.0016f
C28547 a_62508_21976# VPWR 0.3396f
C28548 a_30836_20452# a_30812_19975# 0.00172f
C28549 a_39268_18840# VPWR 0.49542f
C28550 a_2724_26344# VPWR 0.20782f
C28551 a_43804_30951# vgaringosc.workerclkbuff_notouch_.I 0.00352f
C28552 a_23868_2727# a_23780_2824# 0.28563f
C28553 a_53260_26399# VPWR 0.00246f
C28554 _355_.C a_20308_27912# 0.00515f
C28555 _345_.A2 a_23060_26724# 0.01232f
C28556 _293_.A2 _402_.A1 0.00617f
C28557 _267_.A2 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I 0.03471f
C28558 a_54780_20408# VPWR 0.31389f
C28559 _327_.A2 a_40668_20408# 0.00545f
C28560 _325_.A1 a_42168_22504# 0.00524f
C28561 _330_.A2 a_38842_17316# 0.00898f
C28562 _474_.CLK a_53572_17316# 0.00204f
C28563 a_57156_9476# a_56796_9432# 0.08717f
C28564 a_58500_9476# a_58948_9476# 0.01328f
C28565 a_4740_1256# a_5188_1256# 0.01328f
C28566 a_4068_28292# VPWR 0.2157f
C28567 _334_.A1 _284_.ZN 0.01748f
C28568 a_45012_29816# a_45088_29123# 0.00103f
C28569 a_5188_31048# a_5636_31048# 0.01328f
C28570 a_38816_27555# a_39796_27912# 0.00702f
C28571 _287_.A1 _359_.B 0.6784f
C28572 a_61948_14136# a_62396_14136# 0.01288f
C28573 a_1828_3204# a_2276_3204# 0.01328f
C28574 a_65892_14180# a_65532_14136# 0.08707f
C28575 a_16500_20452# a_16588_20408# 0.28563f
C28576 _448_.Q _441_.A2 0.19486f
C28577 a_34080_22461# a_34715_22137# 0.02112f
C28578 a_52640_29860# _267_.ZN 0.00175f
C28579 a_18716_30951# uio_out[7] 0.00872f
C28580 a_22076_1592# a_22212_1256# 0.00168f
C28581 a_52340_13800# a_52428_12135# 0.00151f
C28582 _397_.A2 a_48988_26369# 0.01082f
C28583 _350_.A2 _223_.ZN 0.55779f
C28584 _251_.A1 a_60276_29032# 0.00975f
C28585 _352_.A2 _457_.D 0.21776f
C28586 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN 0.63655f
C28587 a_41340_1159# VPWR 0.33277f
C28588 a_4604_29816# a_4740_29480# 0.00168f
C28589 a_54780_1159# a_55140_1256# 0.08717f
C28590 _261_.ZN _438_.ZN 0.12309f
C28591 a_2276_11044# a_2724_11044# 0.01328f
C28592 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN a_62796_25640# 0.00126f
C28593 a_62732_16839# a_63180_16839# 0.0131f
C28594 a_30812_1592# a_31260_1592# 0.01288f
C28595 _467_.D a_17168_27165# 0.00732f
C28596 _242_.Z vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I 0.03695f
C28597 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN a_55140_20452# 0.00467f
C28598 a_34155_25273# a_34756_24776# 0.00172f
C28599 _229_.I a_60964_27912# 0.00546f
C28600 _304_.A1 a_34980_22895# 0.41924f
C28601 _360_.ZN _359_.ZN 0.0013f
C28602 a_2724_18504# a_2724_17316# 0.05841f
C28603 a_60268_10567# a_60180_10664# 0.28563f
C28604 _462_.D uo_out[7] 0.0032f
C28605 a_37386_31048# uo_out[3] 0.00254f
C28606 a_53572_21640# a_54020_21640# 0.01328f
C28607 a_20084_22020# VPWR 0.20622f
C28608 _287_.A1 a_36656_29123# 0.00121f
C28609 a_38616_24328# _430_.ZN 0.03085f
C28610 a_42154_21236# VPWR 0.8211f
C28611 a_26668_23544# VPWR 0.32414f
C28612 a_3260_18840# a_3708_18840# 0.0131f
C28613 a_30140_21543# a_30500_21640# 0.08707f
C28614 a_21404_2727# VPWR 0.31143f
C28615 a_3172_13800# VPWR 0.20993f
C28616 a_56124_23111# VPWR 0.31627f
C28617 a_22100_31048# a_22188_29383# 0.00248f
C28618 a_18760_29032# uio_out[7] 0.41806f
C28619 a_57940_20452# a_58028_20408# 0.28563f
C28620 a_7540_31048# uio_oe[6] 0.00129f
C28621 _274_.A3 _267_.ZN 0.00103f
C28622 a_6308_29860# VPWR 0.2085f
C28623 a_58140_11000# VPWR 0.35527f
C28624 a_40668_26247# a_41028_26344# 0.08674f
C28625 _245_.Z a_61836_25515# 0.22862f
C28626 a_14796_21976# a_14796_21543# 0.05841f
C28627 a_63516_15704# a_63516_15271# 0.05841f
C28628 a_18740_22020# a_18716_21543# 0.00172f
C28629 _325_.A1 a_40780_21543# 0.00291f
C28630 _223_.ZN a_31516_28292# 0.00476f
C28631 _441_.A3 _300_.ZN 0.59111f
C28632 _359_.B _293_.A2 0.05281f
C28633 _363_.Z _452_.CLK 0.01467f
C28634 _437_.A1 a_37532_26247# 0.00599f
C28635 a_46198_27060# a_44744_26355# 0.00562f
C28636 a_932_2824# a_1380_2824# 0.01328f
C28637 a_34620_2727# a_35204_2824# 0.01675f
C28638 a_62060_23111# a_62420_23208# 0.08717f
C28639 _256_.A2 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN 1.86223f
C28640 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN a_59172_23588# 0.00112f
C28641 a_39796_22504# a_40004_22020# 0.01751f
C28642 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN 0.23414f
C28643 a_65108_23588# a_65556_23588# 0.01328f
C28644 a_50384_19204# a_50280_19369# 0.10745f
C28645 _419_.A4 _421_.B 0.12982f
C28646 _448_.Q a_39772_19975# 0.0012f
C28647 _407_.A1 a_50704_27912# 0.0061f
C28648 a_65220_3204# a_64860_3160# 0.08717f
C28649 a_1916_3160# a_1916_2727# 0.05841f
C28650 a_1020_4728# a_1020_4295# 0.05841f
C28651 _251_.A1 a_61052_26247# 0.00599f
C28652 a_21740_20408# a_22324_20452# 0.01675f
C28653 a_47776_20893# a_47259_20127# 0.00602f
C28654 _452_.CLK a_36960_27912# 0.02496f
C28655 a_7628_30951# a_7540_31048# 0.28563f
C28656 _383_.A2 _390_.ZN 0.14722f
C28657 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I 0.00631f
C28658 a_14596_1636# VPWR 0.20348f
C28659 a_60292_12612# a_60380_12568# 0.28563f
C28660 a_63404_23111# vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I 0.00147f
C28661 a_56348_12568# a_56796_12568# 0.01288f
C28662 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I a_62279_28293# 0.00176f
C28663 _359_.B a_28000_29480# 0.04439f
C28664 a_59260_23111# a_59172_23208# 0.28563f
C28665 a_11548_29816# a_11684_29480# 0.00168f
C28666 a_63740_1159# VPWR 0.29679f
C28667 a_66204_1159# a_66116_1256# 0.28563f
C28668 a_3260_19975# VPWR 0.30487f
C28669 a_4940_18407# VPWR 0.31945f
C28670 a_38116_1636# a_37756_1592# 0.08707f
C28671 _305_.A2 a_45396_22020# 0.01347f
C28672 a_23332_26344# VPWR 0.13442f
C28673 a_36436_18504# a_36548_17316# 0.02666f
C28674 a_26108_1159# a_26556_1159# 0.0131f
C28675 a_57044_10664# a_57492_10664# 0.01328f
C28676 a_43003_28409# VPWR 0.35986f
C28677 a_19076_24776# a_19164_23111# 0.00151f
C28678 _459_.CLK a_26916_27912# 0.0098f
C28679 a_26220_21976# VPWR 0.33593f
C28680 _384_.ZN _417_.A2 0.00582f
C28681 a_54444_25112# a_54444_24679# 0.05841f
C28682 _324_.C a_45128_26031# 0.00755f
C28683 _452_.CLK a_33276_23111# 0.02566f
C28684 _304_.ZN a_42982_21730# 0.08451f
C28685 a_43804_2727# VPWR 0.31143f
C28686 a_64884_13800# VPWR 0.23091f
C28687 a_44632_30206# VPWR 0.5052f
C28688 a_56036_2824# a_56124_1159# 0.0027f
C28689 a_28708_21640# a_29156_21640# 0.01328f
C28690 a_4156_26247# a_4068_26344# 0.28563f
C28691 _284_.ZN _448_.Q 0.00128f
C28692 a_58687_31220# ui_in[2] 0.0012f
C28693 a_12444_29816# VPWR 0.29679f
C28694 _346_.A2 _351_.A2 0.25466f
C28695 a_66900_16936# a_67012_15748# 0.02666f
C28696 a_5388_10567# VPWR 0.35526f
C28697 a_32156_15271# a_32068_15368# 0.28563f
C28698 a_31036_23111# VPWR 0.31557f
C28699 _452_.CLK _325_.ZN 0.05501f
C28700 a_56572_2727# a_56708_1636# 0.00154f
C28701 _327_.A2 a_40780_21543# 0.02226f
C28702 _447_.Q a_38576_22504# 0.16042f
C28703 _379_.A2 a_20379_29977# 0.05694f
C28704 _324_.B a_44500_22020# 0.02127f
C28705 a_33500_15271# a_33948_15271# 0.0131f
C28706 _229_.I a_63105_28293# 0.15453f
C28707 a_46624_19715# a_46252_19759# 0.10745f
C28708 a_59620_27208# a_60828_26680# 0.00445f
C28709 a_932_22020# a_1380_22020# 0.01328f
C28710 a_46044_2727# a_45956_2824# 0.28563f
C28711 a_62532_17316# a_62172_17272# 0.08717f
C28712 a_52512_19715# a_52924_20127# 0.00275f
C28713 a_54444_19975# a_54356_20072# 0.28563f
C28714 a_45732_18884# VPWR 0.13565f
C28715 a_66116_17316# a_66564_17316# 0.01328f
C28716 a_62396_26247# VPWR 0.31983f
C28717 _251_.A1 _249_.A2 0.09505f
C28718 a_18380_23544# a_18828_23544# 0.01288f
C28719 a_3260_7431# a_3708_7431# 0.0131f
C28720 a_2364_8999# a_2812_8999# 0.0131f
C28721 _355_.C a_27004_27815# 0.00162f
C28722 a_26916_1256# a_27588_1256# 0.00347f
C28723 a_66652_7864# a_66652_7431# 0.05841f
C28724 a_4156_5863# a_4940_5863# 0.00443f
C28725 a_67548_6296# a_67548_5863# 0.05841f
C28726 _474_.CLK a_54692_20452# 0.01403f
C28727 a_2364_13703# a_2724_13800# 0.08717f
C28728 a_6172_2727# a_6620_2727# 0.0131f
C28729 a_31396_31048# a_31088_30301# 0.0022f
C28730 a_56012_13703# a_56460_13703# 0.012f
C28731 a_38228_16936# a_38428_15271# 0.00119f
C28732 a_27476_20452# a_27564_20408# 0.28563f
C28733 _416_.A1 a_44795_29535# 0.01126f
C28734 a_3708_16839# a_4068_16936# 0.08717f
C28735 _457_.D a_24900_24776# 0.00467f
C28736 a_20732_1592# VPWR 0.3289f
C28737 _427_.B1 a_53076_24776# 0.00175f
C28738 _419_.Z a_47776_20893# 0.01752f
C28739 a_9635_30644# a_10092_30951# 0.00916f
C28740 a_63652_12612# a_63740_12568# 0.28563f
C28741 _324_.C _267_.ZN 0.03608f
C28742 a_1468_23544# a_1468_23111# 0.05841f
C28743 _325_.A1 a_42996_18840# 0.05514f
C28744 _417_.A2 a_49068_20408# 0.08463f
C28745 _334_.A1 _223_.ZN 0.0096f
C28746 a_67572_12232# a_67684_11044# 0.02666f
C28747 a_66876_15271# a_66788_15368# 0.28563f
C28748 a_51196_11000# a_51644_11000# 0.01288f
C28749 a_41028_1636# a_41116_1592# 0.28563f
C28750 a_44612_1636# a_45060_1636# 0.01328f
C28751 a_42484_16936# a_42932_16936# 0.01328f
C28752 _402_.A1 a_47297_25596# 0.00222f
C28753 _304_.A1 a_38529_22804# 0.00456f
C28754 _324_.C _390_.ZN 0.23123f
C28755 a_4964_26724# a_4604_26680# 0.08674f
C28756 a_2364_26680# a_2812_26680# 0.0131f
C28757 _474_.CLK _275_.ZN 0.04267f
C28758 _346_.B _455_.D 0.0109f
C28759 _336_.A2 a_28756_25940# 0.00384f
C28760 a_21652_29480# VPWR 0.12127f
C28761 _290_.ZN uo_out[4] 0.14719f
C28762 _355_.B _355_.ZN 0.08485f
C28763 _336_.A2 a_27172_24328# 0.39666f
C28764 a_1916_20408# VPWR 0.297f
C28765 _388_.B a_45956_31048# 0.00151f
C28766 _452_.Q a_40244_21640# 0.04634f
C28767 a_46268_12568# VPWR 0.29679f
C28768 a_66204_2727# VPWR 0.31654f
C28769 a_7068_2727# a_7204_1636# 0.00154f
C28770 a_6980_2824# a_7428_2824# 0.01328f
C28771 a_19076_26344# a_19524_26344# 0.01328f
C28772 a_41028_26344# _451_.Q 0.00459f
C28773 _251_.A1 a_62564_29032# 0.05895f
C28774 a_4828_29383# a_5188_29480# 0.08717f
C28775 a_35492_20072# VPWR 0.01469f
C28776 a_1468_28248# a_1468_27815# 0.05841f
C28777 _416_.A1 a_44571_26841# 0.06645f
C28778 a_5052_15704# a_4940_15271# 0.02634f
C28779 _371_.A3 a_26916_27912# 0.00566f
C28780 a_66764_10567# VPWR 0.31389f
C28781 a_61524_20452# a_61972_20452# 0.01328f
C28782 a_43132_15271# a_43492_15368# 0.08717f
C28783 a_31372_21976# a_31484_21543# 0.02634f
C28784 a_28708_23208# VPWR 0.20595f
C28785 _334_.A1 a_32592_25227# 0.00126f
C28786 a_38616_24328# _441_.A3 0.00619f
C28787 a_34396_24679# a_33932_24073# 0.00104f
C28788 a_14708_28292# a_14796_28248# 0.28563f
C28789 a_15604_28292# a_16052_28292# 0.01328f
C28790 _395_.A1 a_47636_25940# 0.00729f
C28791 _336_.A2 a_27884_25641# 0.02572f
C28792 a_64324_15748# VPWR 0.20801f
C28793 a_12916_31048# uio_oe[2] 0.00354f
C28794 a_57020_2727# a_57380_2824# 0.08717f
C28795 _327_.Z a_41572_20072# 0.01909f
C28796 a_55788_23544# clk 0.00613f
C28797 _358_.A3 a_35140_26680# 0.50927f
C28798 _311_.Z _301_.A1 0.65302f
C28799 a_49764_26724# a_50120_26476# 0.00215f
C28800 a_31920_29480# uo_out[6] 0.05861f
C28801 a_53012_18504# a_53460_18504# 0.01328f
C28802 _452_.CLK a_35660_27508# 0.00518f
C28803 a_26132_23588# a_26220_23544# 0.28563f
C28804 a_17036_25112# a_17484_25112# 0.01288f
C28805 a_4516_4772# VPWR 0.20862f
C28806 a_20980_25156# a_21068_25112# 0.28563f
C28807 a_11460_31048# VPWR 0.2534f
C28808 a_8548_1256# VPWR 0.22423f
C28809 _417_.A2 a_48776_20204# 0.40283f
C28810 a_2724_7908# VPWR 0.20782f
C28811 _251_.A1 a_63092_26724# 0.00875f
C28812 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.02585f
C28813 a_30812_18840# a_30812_18407# 0.05841f
C28814 _419_.A4 a_47524_22021# 0.04006f
C28815 _260_.ZN a_42252_20936# 0.04547f
C28816 a_53324_13703# a_53236_13800# 0.28563f
C28817 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_56684_23544# 0.00174f
C28818 _424_.A2 a_52240_22504# 0.00443f
C28819 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN 0.72599f
C28820 a_32716_20408# a_33164_20408# 0.0131f
C28821 a_26556_30951# a_27004_30951# 0.012f
C28822 _400_.ZN a_45577_27509# 0.00788f
C28823 _285_.Z VPWR 1.16046f
C28824 a_40132_26344# _261_.ZN 0.00262f
C28825 _431_.A3 _444_.D 0.04204f
C28826 a_53908_25156# a_53996_25112# 0.28563f
C28827 a_40108_16839# a_40020_16936# 0.28563f
C28828 _304_.A1 _304_.ZN 0.62455f
C28829 _327_.A2 a_42996_18840# 0.00121f
C28830 a_66540_16839# VPWR 0.3163f
C28831 a_34532_1636# VPWR 0.21168f
C28832 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I 0.00596f
C28833 _251_.A1 a_60516_26344# 0.00466f
C28834 a_3260_12135# a_3708_12135# 0.0131f
C28835 a_44476_27815# VPWR 0.32095f
C28836 a_21428_23588# a_21404_23111# 0.00172f
C28837 a_17484_23544# a_17484_23111# 0.05841f
C28838 a_7652_1636# a_8100_1636# 0.01328f
C28839 a_4068_1636# a_4156_1592# 0.28563f
C28840 _330_.A1 a_35723_20569# 0.00469f
C28841 a_2276_17316# a_2364_17272# 0.28563f
C28842 a_58500_11044# a_58140_11000# 0.08707f
C28843 a_20196_1636# a_20060_1159# 0.00168f
C28844 a_61076_12232# a_61164_10567# 0.00151f
C28845 a_44948_25156# VPWR 0.0086f
C28846 a_57492_17316# a_57580_17272# 0.28563f
C28847 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_54692_26344# 0.00425f
C28848 a_48508_1159# a_48956_1159# 0.0131f
C28849 a_37444_2824# a_37308_1592# 0.00154f
C28850 a_53436_18840# VPWR 0.33579f
C28851 _304_.B _267_.A1 0.17808f
C28852 a_62084_18884# a_62172_18840# 0.28563f
C28853 a_66116_18884# a_66564_18884# 0.01328f
C28854 a_2276_25156# VPWR 0.20634f
C28855 a_60916_29612# VPWR 0.00502f
C28856 a_1916_27815# a_1828_27912# 0.28563f
C28857 a_25460_20452# VPWR 0.21526f
C28858 a_1020_15704# a_1468_15704# 0.0131f
C28859 a_59932_12568# VPWR 0.31547f
C28860 a_3620_15748# a_3260_15704# 0.08717f
C28861 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I 0.16719f
C28862 a_35292_15704# a_35428_15368# 0.00168f
C28863 a_52452_15368# a_52900_15368# 0.01328f
C28864 a_16252_29383# a_16164_29480# 0.28563f
C28865 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN 0.00586f
C28866 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I a_55364_21640# 0.0059f
C28867 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN 0.02382f
C28868 a_932_7528# a_1380_7528# 0.01328f
C28869 a_4156_8999# a_4852_9096# 0.01227f
C28870 a_60628_10664# VPWR 0.20641f
C28871 _304_.B _408_.ZN 0.09597f
C28872 a_54556_15271# a_54468_15368# 0.28563f
C28873 a_64860_5863# a_65220_5960# 0.08717f
C28874 _255_.I a_59796_29480# 0.00219f
C28875 _294_.A2 a_37844_29860# 0.00299f
C28876 a_65756_4295# a_66116_4392# 0.08717f
C28877 _476_.Q a_52024_20083# 0.00589f
C28878 a_55900_15271# a_56348_15271# 0.0131f
C28879 _251_.A1 a_59226_25156# 0.00253f
C28880 a_51988_24776# VPWR 0.00419f
C28881 a_33860_15368# VPWR 0.21418f
C28882 a_19276_21976# a_19724_21976# 0.01288f
C28883 _395_.A3 _424_.A1 0.08918f
C28884 a_932_2824# a_932_1636# 0.05841f
C28885 _371_.A1 a_31396_26724# 0.00116f
C28886 a_37308_15271# VPWR 0.32932f
C28887 a_2276_14180# a_2364_14136# 0.28563f
C28888 a_37420_16839# a_37868_16839# 0.01288f
C28889 _304_.B a_47172_27912# 0.00391f
C28890 a_41364_16936# a_41252_15748# 0.02666f
C28891 a_26668_23544# a_26580_22020# 0.00151f
C28892 a_43664_17317# VPWR 0.59274f
C28893 vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN a_64884_26724# 0.00591f
C28894 a_32820_29535# VPWR 0.00246f
C28895 a_14460_30951# uio_oe[2] 0.00741f
C28896 a_30924_23544# a_31372_23544# 0.01255f
C28897 a_32180_23588# a_32268_23544# 0.28563f
C28898 a_33636_23208# a_33724_21543# 0.00227f
C28899 a_30724_1256# VPWR 0.20968f
C28900 a_65756_7431# VPWR 0.31505f
C28901 a_49316_1256# a_49764_1256# 0.01328f
C28902 a_67548_4295# VPWR 0.32135f
C28903 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN 0.88258f
C28904 a_51048_26680# _384_.A3 0.4942f
C28905 a_50100_13800# a_50548_13800# 0.01328f
C28906 a_64772_3204# a_64636_2727# 0.00168f
C28907 a_28572_2727# a_29020_2727# 0.0131f
C28908 a_63852_13703# a_64212_13800# 0.08663f
C28909 a_61860_26344# VPWR 0.20348f
C28910 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN 0.6226f
C28911 _370_.ZN _352_.A2 0.40897f
C28912 a_39748_31048# VPWR 0.01438f
C28913 a_14004_31048# VPWR 0.36263f
C28914 a_50860_16839# a_51220_16936# 0.08717f
C28915 a_64324_18504# VPWR 0.20554f
C28916 a_54132_10664# a_54244_9476# 0.02666f
C28917 _358_.A3 _460_.D 0.05405f
C28918 a_40668_1592# VPWR 0.3289f
C28919 a_54432_31128# _274_.A1 0.00208f
C28920 a_21852_23111# a_21876_22020# 0.0016f
C28921 a_50300_1592# a_50436_1256# 0.00168f
C28922 a_9980_1159# a_9892_1256# 0.28563f
C28923 a_46068_16936# VPWR 0.20944f
C28924 _416_.A1 _436_.ZN 0.16087f
C28925 a_46984_23588# a_47636_23588# 0.00195f
C28926 _452_.CLK a_36188_26680# 0.02294f
C28927 a_28372_23588# a_28348_23111# 0.00172f
C28928 a_5500_29816# a_5948_29816# 0.01288f
C28929 a_32068_17316# a_32156_17272# 0.28563f
C28930 a_35652_17316# a_36100_17316# 0.01328f
C28931 _416_.ZN a_47724_18840# 0.00303f
C28932 a_51556_15368# a_51556_14180# 0.05841f
C28933 _459_.CLK a_31964_28292# 0.00458f
C28934 a_21292_30951# uio_out[4] 0.00366f
C28935 a_47748_15368# a_47612_14136# 0.00154f
C28936 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I 0.09388f
C28937 a_27140_1636# a_27004_1159# 0.00168f
C28938 a_50748_1592# a_51196_1592# 0.01288f
C28939 a_54692_1636# a_54780_1592# 0.28563f
C28940 a_64996_11044# a_65444_11044# 0.01328f
C28941 a_61860_11044# a_61500_11000# 0.08707f
C28942 a_10788_2824# VPWR 0.21382f
C28943 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN 0.7848f
C28944 _393_.A3 a_47924_28292# 0.00142f
C28945 _397_.A2 _393_.A1 0.03524f
C28946 a_37444_26724# VPWR 0.21366f
C28947 _359_.B a_34308_26344# 0.05658f
C28948 a_16140_23111# a_16588_23111# 0.0131f
C28949 _459_.CLK a_16052_26344# 0.0063f
C28950 _416_.A2 a_47776_20893# 0.03473f
C28951 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN a_53908_18504# 0.00345f
C28952 a_54444_18407# a_54804_18504# 0.08663f
C28953 a_64324_15368# VPWR 0.21723f
C28954 _412_.B2 clk 0.01046f
C28955 _267_.A1 VPWR 0.50956f
C28956 a_4604_4728# a_4516_3204# 0.0027f
C28957 a_20620_25112# VPWR 0.31547f
C28958 a_16500_27912# a_16948_27912# 0.01328f
C28959 _255_.ZN a_58116_30344# 0.41672f
C28960 _427_.ZN a_54244_20452# 0.00422f
C28961 a_46716_12135# VPWR 0.29679f
C28962 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN 0.01254f
C28963 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I _250_.A2 0.00662f
C28964 a_33412_15748# a_33052_15704# 0.08707f
C28965 _336_.Z _459_.D 0.0119f
C28966 _340_.A2 a_25962_29480# 0.01244f
C28967 a_29380_2824# a_29828_2824# 0.01328f
C28968 _397_.A1 a_47636_25940# 0.21088f
C28969 _388_.B _474_.CLK 0.10625f
C28970 a_44160_29123# a_43788_29167# 0.10745f
C28971 a_37408_23208# VPWR 0.01436f
C28972 a_62404_25156# VPWR 0.00966f
C28973 _251_.A1 _250_.B 0.24096f
C28974 a_44028_15704# a_44028_15271# 0.05841f
C28975 a_38788_20072# VPWR 0.12664f
C28976 _408_.ZN VPWR 0.76204f
C28977 a_19972_21640# a_19948_20408# 0.0016f
C28978 a_57940_17316# vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN 0.00117f
C28979 a_21764_21640# a_21652_20452# 0.02666f
C28980 _304_.B _412_.A1 0.10684f
C28981 a_4604_15704# VPWR 0.33016f
C28982 a_56260_15368# VPWR 0.20348f
C28983 _301_.A1 a_39780_22805# 0.00143f
C28984 _275_.A2 _324_.C 0.16727f
C28985 a_1380_9476# a_1828_9476# 0.01328f
C28986 a_55252_24776# clk 0.0155f
C28987 a_26580_22020# a_26220_21976# 0.08707f
C28988 _330_.A1 a_38616_24328# 0.03185f
C28989 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN VPWR 0.81904f
C28990 a_46628_14180# a_46716_14136# 0.28563f
C28991 a_50212_14180# a_50660_14180# 0.01328f
C28992 a_37980_17272# a_37892_15748# 0.00151f
C28993 a_47172_27912# VPWR 0.00677f
C28994 _247_.B a_60068_27912# 0.10199f
C28995 a_5052_21976# a_4964_20452# 0.00151f
C28996 _343_.A2 _345_.A2 0.39489f
C28997 a_32268_23544# a_32180_22020# 0.00151f
C28998 a_41004_16839# VPWR 0.32214f
C28999 a_48308_16936# a_48196_15748# 0.02666f
C29000 _450_.D _325_.B 0.09939f
C29001 a_53124_1256# VPWR 0.20348f
C29002 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I a_56148_24776# 0.00702f
C29003 a_64636_14136# a_64548_12612# 0.0027f
C29004 a_58388_17316# VPWR 0.23733f
C29005 a_42896_18504# a_44276_17316# 0.00999f
C29006 _474_.CLK a_54444_25112# 0.03044f
C29007 _421_.A1 a_47047_21640# 0.0082f
C29008 a_31708_17272# VPWR 0.29679f
C29009 a_61524_10664# a_61412_9476# 0.02666f
C29010 a_28796_23111# a_28820_22020# 0.0016f
C29011 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I 0.01017f
C29012 a_54332_1592# VPWR 0.29679f
C29013 a_20956_1159# a_21316_1256# 0.08717f
C29014 a_57244_1592# a_57380_1256# 0.00168f
C29015 a_64972_12135# a_65420_12135# 0.0131f
C29016 a_51084_12135# a_51444_12232# 0.08707f
C29017 a_23980_23544# a_24004_23208# 0.00172f
C29018 a_13788_1592# a_14236_1592# 0.01288f
C29019 a_14148_29480# a_14596_29480# 0.01328f
C29020 a_24080_25227# a_24452_24776# 0.00113f
C29021 a_12804_29860# a_12444_29816# 0.08707f
C29022 _355_.C _375_.Z 0.00812f
C29023 a_39236_17316# a_39324_17272# 0.28563f
C29024 _317_.A2 a_37084_21543# 0.00184f
C29025 a_33188_2824# VPWR 0.2051f
C29026 a_58052_1636# a_57692_1592# 0.08707f
C29027 _371_.A1 VPWR 2.02221f
C29028 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN a_59172_22020# 0.00618f
C29029 a_932_24776# a_1380_24776# 0.01328f
C29030 a_19164_24679# a_19076_24776# 0.28563f
C29031 a_15244_23111# a_15156_23208# 0.28563f
C29032 _444_.D a_36748_23544# 0.00277f
C29033 a_4964_9476# VPWR 0.21167f
C29034 a_64772_9096# a_65220_9096# 0.01328f
C29035 a_67996_7864# a_67908_6340# 0.0027f
C29036 a_65668_7528# a_66116_7528# 0.01328f
C29037 a_66564_5960# a_67012_5960# 0.01328f
C29038 a_46268_14136# VPWR 0.29679f
C29039 a_31260_18407# a_31620_18504# 0.08717f
C29040 _442_.ZN _438_.A2 0.00413f
C29041 a_36212_23588# a_36300_23544# 0.28563f
C29042 a_39908_15748# a_40356_15748# 0.01328f
C29043 a_932_12232# VPWR 0.22176f
C29044 _304_.B a_40668_20408# 0.00717f
C29045 a_4852_24776# VPWR 0.22733f
C29046 _412_.A1 VPWR 1.00302f
C29047 a_1020_2727# a_1380_2824# 0.08717f
C29048 a_43492_15748# VPWR 0.20692f
C29049 a_2812_19975# a_2724_20072# 0.28563f
C29050 _231_.I vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN 0.03048f
C29051 a_43008_26795# a_43396_27209# 0.00393f
C29052 a_43936_27165# a_44571_26841# 0.02112f
C29053 _311_.Z a_37296_22020# 0.00869f
C29054 a_45732_9476# a_45820_9432# 0.28563f
C29055 _301_.A1 a_39796_22504# 0.07233f
C29056 a_30924_21976# a_31372_21976# 0.01255f
C29057 a_32180_22020# a_32268_21976# 0.28563f
C29058 _417_.A2 a_51540_23588# 0.00327f
C29059 a_41384_26841# VPWR 0.00219f
C29060 _334_.A1 a_37888_27555# 0.00284f
C29061 a_36960_27912# a_38816_27555# 0.02307f
C29062 _408_.ZN a_50068_27508# 0.37644f
C29063 a_7740_1592# a_7876_1256# 0.00168f
C29064 a_4068_12612# a_4516_12612# 0.01328f
C29065 a_30476_25112# VPWR 0.33084f
C29066 a_2276_12612# a_1916_12568# 0.08717f
C29067 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I a_66676_20452# 0.00476f
C29068 a_50972_2727# a_51420_2727# 0.0131f
C29069 _284_.ZN _234_.ZN 0.02145f
C29070 a_49628_17272# a_49740_16839# 0.02634f
C29071 a_53572_17316# a_53548_16839# 0.00172f
C29072 _447_.Q a_43600_22504# 0.00132f
C29073 _424_.B1 _412_.ZN 0.08028f
C29074 a_58276_25156# VPWR 0.25255f
C29075 a_29232_29931# a_30160_30301# 1.16391f
C29076 a_51332_17316# VPWR 0.20694f
C29077 a_62060_12135# a_61972_12232# 0.28563f
C29078 a_63740_1592# VPWR 0.30141f
C29079 a_32380_1159# a_32292_1256# 0.28563f
C29080 a_65980_1592# a_66116_1256# 0.00168f
C29081 _378_.I a_22100_29480# 0.00157f
C29082 a_22100_31048# uio_out[4] 0.00733f
C29083 a_21092_1636# a_20732_1592# 0.08707f
C29084 _313_.ZN a_33188_23208# 0.00101f
C29085 _229_.I a_60156_27815# 0.00633f
C29086 _427_.B1 _419_.Z 0.00958f
C29087 a_17596_29816# a_18044_29816# 0.01255f
C29088 a_16612_29860# _459_.CLK 0.00208f
C29089 _276_.A2 a_53592_30344# 0.00159f
C29090 a_24092_21543# VPWR 0.31547f
C29091 _379_.A2 a_18264_29480# 0.10235f
C29092 a_16500_26344# a_16500_25156# 0.05841f
C29093 _451_.Q a_38576_22504# 0.00122f
C29094 _282_.ZN _284_.B 0.65817f
C29095 a_47748_17316# a_48196_17316# 0.01328f
C29096 a_51980_10567# a_52428_10567# 0.01288f
C29097 a_64548_1636# a_64996_1636# 0.01328f
C29098 _384_.A3 a_51988_24072# 0.00376f
C29099 a_55588_2824# VPWR 0.20812f
C29100 a_65980_11000# a_65868_10567# 0.02634f
C29101 a_51968_26724# VPWR 0.01428f
C29102 a_4852_23208# a_5300_23208# 0.01328f
C29103 a_25884_23111# a_26468_23208# 0.01675f
C29104 _281_.A1 a_54040_22366# 0.18293f
C29105 uio_in[7] uio_in[6] 0.01021f
C29106 a_54692_9476# VPWR 0.20692f
C29107 a_22212_2824# a_22300_1159# 0.0027f
C29108 a_61860_14180# VPWR 0.20948f
C29109 a_20508_21543# a_20956_21543# 0.01288f
C29110 _441_.ZN a_39587_24372# 0.00122f
C29111 a_36436_18504# _330_.ZN 0.00159f
C29112 _452_.CLK a_34756_24776# 0.01994f
C29113 _324_.C _399_.A1 0.00101f
C29114 _304_.B a_42168_22504# 0.087f
C29115 a_62420_12232# VPWR 0.20622f
C29116 a_51780_2824# a_52228_2824# 0.01328f
C29117 a_35292_2727# a_35428_1636# 0.00154f
C29118 a_40668_20408# VPWR 0.32114f
C29119 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I VPWR 1.03976f
C29120 a_5724_30951# a_5860_29860# 0.00154f
C29121 _288_.ZN a_37584_29123# 0.0012f
C29122 a_67796_20072# VPWR 0.2115f
C29123 a_12444_2727# a_12356_2824# 0.28563f
C29124 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN a_63404_20408# 0.00969f
C29125 _350_.A2 a_30520_27508# 0.00164f
C29126 a_60401_30300# _324_.C 0.0179f
C29127 _342_.ZN _340_.ZN 0.50813f
C29128 a_49628_15704# VPWR 0.33528f
C29129 _452_.Q a_40132_20072# 0.08362f
C29130 _355_.C a_22059_26399# 0.00987f
C29131 _243_.ZN a_58052_26724# 0.00485f
C29132 _324_.C _325_.A1 0.06285f
C29133 a_48508_30951# a_48708_29816# 0.00159f
C29134 a_50972_9432# a_51420_9432# 0.0131f
C29135 a_35504_18955# a_35652_17316# 0.0013f
C29136 a_18180_31048# uio_out[7] 0.01794f
C29137 _301_.A1 a_35816_21192# 0.00161f
C29138 a_57244_14136# a_57692_14136# 0.012f
C29139 a_63876_15368# a_63852_13703# 0.00131f
C29140 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I 0.20189f
C29141 _284_.ZN _284_.A2 1.3203f
C29142 a_5052_11000# a_4964_9476# 0.00151f
C29143 _402_.A1 _436_.B 0.06012f
C29144 _274_.ZN a_51665_30344# 0.0039f
C29145 a_46628_12612# a_46268_12568# 0.08707f
C29146 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN 0.08247f
C29147 a_33636_23208# a_33152_22091# 0.00263f
C29148 a_21404_24679# a_21428_23588# 0.0016f
C29149 a_18492_1159# VPWR 0.30281f
C29150 _323_.A3 a_36836_20072# 0.01909f
C29151 a_43356_1159# a_43716_1256# 0.08717f
C29152 a_27588_1636# a_28036_1636# 0.01328f
C29153 a_58836_12232# a_59284_12232# 0.01328f
C29154 a_49764_26724# a_48384_26724# 0.00295f
C29155 _427_.A2 a_54420_21976# 0.00218f
C29156 a_21316_21640# VPWR 0.20641f
C29157 _350_.A1 _294_.A2 0.08377f
C29158 _452_.CLK a_40132_26344# 0.00546f
C29159 a_62844_11000# a_62868_10664# 0.00172f
C29160 a_49292_10567# a_49204_10664# 0.28563f
C29161 _419_.A4 _402_.B 0.02475f
C29162 a_59172_23208# VPWR 0.14647f
C29163 a_33612_24679# a_34396_24679# 0.00443f
C29164 _304_.B a_40780_21543# 0.00786f
C29165 a_30796_24463# a_31140_24831# 0.00275f
C29166 a_18740_23588# VPWR 0.21276f
C29167 a_65668_9476# VPWR 0.21537f
C29168 a_51912_20452# VPWR 0.61603f
C29169 a_64412_6296# VPWR 0.3038f
C29170 a_48508_13703# VPWR 0.31817f
C29171 a_55252_20072# VPWR 0.20922f
C29172 a_19164_21543# a_19524_21640# 0.08707f
C29173 _438_.A2 _435_.ZN 0.6492f
C29174 a_64324_20072# a_64772_20072# 0.01328f
C29175 _407_.ZN a_52316_27815# 0.01027f
C29176 a_66204_3160# VPWR 0.31657f
C29177 a_18816_29931# uio_out[7] 0.02196f
C29178 _349_.A4 uio_out[2] 0.00316f
C29179 _258_.I _274_.A2 0.39955f
C29180 a_42168_22504# VPWR 0.03623f
C29181 _459_.CLK a_27228_26680# 0.0477f
C29182 a_49988_15748# a_50076_15704# 0.28563f
C29183 a_51556_11044# VPWR 0.20622f
C29184 a_42236_2727# a_42372_1636# 0.00154f
C29185 vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I 0.00303f
C29186 _337_.A3 _355_.B 0.01818f
C29187 _304_.A1 _441_.B 0.15442f
C29188 a_58052_26724# a_58140_26680# 0.28563f
C29189 _427_.B1 _424_.A1 0.03256f
C29190 a_67908_22020# VPWR 0.15788f
C29191 a_2276_26344# VPWR 0.20634f
C29192 a_52304_26399# VPWR 0.00204f
C29193 a_43356_30951# vgaringosc.workerclkbuff_notouch_.I 0.00225f
C29194 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN 0.70783f
C29195 a_23196_2727# a_23780_2824# 0.01675f
C29196 _324_.C _327_.A2 0.7387f
C29197 a_54332_20408# VPWR 0.31389f
C29198 _355_.C a_19860_27912# 0.00467f
C29199 _384_.A1 a_55340_23544# 0.0022f
C29200 a_3620_28292# VPWR 0.22347f
C29201 _474_.CLK a_53124_17316# 0.00202f
C29202 a_56708_9476# a_56796_9432# 0.28563f
C29203 a_65444_14180# a_65532_14136# 0.28563f
C29204 a_16500_20452# a_16140_20408# 0.08717f
C29205 a_18268_30951# uio_out[7] 0.01566f
C29206 _231_.ZN vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I 0.0023f
C29207 a_60909_30600# a_61860_30736# 0.01935f
C29208 a_53124_12612# a_53572_12612# 0.01328f
C29209 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I a_64324_20072# 0.00108f
C29210 _397_.A2 a_48560_26369# 0.00909f
C29211 a_6396_29816# uio_oe[7] 0.00276f
C29212 a_54780_1159# a_54692_1256# 0.28563f
C29213 _346_.A2 a_24860_27209# 0.00145f
C29214 _304_.A1 _328_.A2 0.00553f
C29215 a_40892_1159# VPWR 0.33008f
C29216 _397_.Z _324_.B 0.03955f
C29217 _467_.D a_16240_26795# 0.2786f
C29218 vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN clk 0.08001f
C29219 a_54420_21976# a_54468_21640# 0.00148f
C29220 _229_.I a_60516_27912# 0.00468f
C29221 a_45732_10664# a_46180_10664# 0.01328f
C29222 _419_.Z _422_.ZN 0.05642f
C29223 a_59820_10567# a_60180_10664# 0.08707f
C29224 a_14684_1159# a_15132_1159# 0.0131f
C29225 a_55228_1592# a_55228_1159# 0.05841f
C29226 a_16164_2824# a_16028_1592# 0.00154f
C29227 a_19636_22020# VPWR 0.21659f
C29228 _287_.A1 a_35728_29480# 0.00883f
C29229 a_40780_21543# VPWR 0.34068f
C29230 a_26220_23544# VPWR 0.33593f
C29231 a_43288_28409# VPWR 0.00214f
C29232 a_17396_21640# a_17844_21640# 0.01328f
C29233 a_30140_21543# a_30052_21640# 0.28563f
C29234 a_20956_2727# VPWR 0.31143f
C29235 a_54088_22895# VPWR 0.18737f
C29236 a_2724_13800# VPWR 0.20782f
C29237 a_61276_15271# a_61724_15271# 0.0131f
C29238 a_5860_29860# VPWR 0.2085f
C29239 a_40668_26247# a_40580_26344# 0.28563f
C29240 a_57692_11000# VPWR 0.32364f
C29241 _267_.A2 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN 0.1678f
C29242 a_66564_15748# a_66428_15271# 0.00168f
C29243 a_64860_15704# a_65308_15704# 0.0131f
C29244 _363_.Z a_35874_27937# 0.01236f
C29245 a_20396_27815# VPWR 0.31549f
C29246 _324_.C vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN 0.0316f
C29247 _370_.B _371_.A1 0.40814f
C29248 _437_.A1 a_37084_26247# 0.00284f
C29249 _474_.CLK a_53660_27815# 0.03324f
C29250 a_34620_2727# a_34532_2824# 0.28563f
C29251 a_53212_29816# vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN 0.29476f
C29252 _409_.ZN a_50468_29977# 0.00242f
C29253 a_62060_23111# a_61972_23208# 0.28563f
C29254 a_49896_18909# a_50280_19369# 1.16391f
C29255 _251_.A1 _245_.Z 0.16108f
C29256 a_63652_9476# a_64324_9476# 0.00347f
C29257 a_61948_9432# a_62396_9432# 0.0131f
C29258 a_15156_23588# a_15604_23588# 0.01328f
C29259 a_15492_1256# a_16164_1256# 0.00347f
C29260 _448_.Q a_39324_19975# 0.00348f
C29261 _330_.A1 _332_.Z 0.02975f
C29262 a_64772_6340# a_65220_6340# 0.01328f
C29263 a_65668_4772# a_66116_4772# 0.01328f
C29264 a_64772_3204# a_64860_3160# 0.28563f
C29265 a_66564_3204# a_67012_3204# 0.01328f
C29266 a_7180_30951# a_7540_31048# 0.08674f
C29267 a_6172_29383# a_6620_29383# 0.0131f
C29268 _383_.A2 a_48141_29480# 0.00103f
C29269 a_60292_12612# a_59932_12568# 0.08663f
C29270 a_62868_13800# a_62956_12135# 0.00151f
C29271 a_14148_1636# VPWR 0.20348f
C29272 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I a_54780_26247# 0.00755f
C29273 _424_.B2 a_51912_20452# 0.33438f
C29274 _459_.CLK a_24080_25227# 0.0116f
C29275 _438_.A2 _441_.ZN 0.53563f
C29276 a_38228_20452# _323_.A3 0.00303f
C29277 a_22560_30288# uio_out[5] 0.00138f
C29278 _336_.A2 a_28596_26725# 0.13359f
C29279 a_63292_1159# VPWR 0.32982f
C29280 a_65756_1159# a_66116_1256# 0.0869f
C29281 a_2812_19975# VPWR 0.30213f
C29282 a_61636_18504# a_61836_16839# 0.00119f
C29283 a_4156_18407# VPWR 0.3269f
C29284 a_5860_1636# a_5724_1159# 0.00168f
C29285 a_1916_1592# a_1916_1159# 0.05841f
C29286 a_33724_1592# a_34172_1592# 0.01288f
C29287 a_37668_1636# a_37756_1592# 0.28563f
C29288 a_35740_25112# a_36188_25112# 0.01255f
C29289 _255_.I a_60276_29032# 0.00479f
C29290 a_47972_11044# a_48420_11044# 0.01328f
C29291 _282_.ZN _474_.Q 0.01469f
C29292 _336_.Z a_29156_23208# 0.00803f
C29293 _424_.B1 _427_.ZN 0.00287f
C29294 a_31172_16936# a_31620_16936# 0.01328f
C29295 _305_.A2 a_44948_22020# 0.00653f
C29296 a_44388_27912# _330_.A1 0.0077f
C29297 hold2.I a_44500_25156# 0.00152f
C29298 a_22344_26399# VPWR 0.00204f
C29299 a_23108_2824# a_22972_1592# 0.00154f
C29300 a_43296_28733# VPWR 0.5136f
C29301 a_25772_21976# VPWR 0.31815f
C29302 a_18028_28777# VPWR 0.40352f
C29303 _324_.C a_45232_25987# 0.05001f
C29304 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN VPWR 0.84714f
C29305 _251_.A1 _252_.B 0.1402f
C29306 _452_.CLK a_32828_23111# 0.05291f
C29307 _304_.ZN a_42778_21812# 0.05032f
C29308 a_64212_13800# VPWR 0.21343f
C29309 a_43828_29860# VPWR 0.14466f
C29310 a_43356_2727# VPWR 0.31143f
C29311 _473_.Q VPWR 1.83277f
C29312 a_17932_26247# a_18716_26247# 0.00443f
C29313 a_3708_26247# a_4068_26344# 0.08717f
C29314 a_61748_16936# a_61724_15271# 0.00144f
C29315 _438_.A2 a_39873_21236# 0.00824f
C29316 a_11996_29816# VPWR 0.33603f
C29317 _346_.A2 a_24900_27912# 0.10906f
C29318 a_63540_16936# a_63516_15704# 0.0016f
C29319 a_4940_10567# VPWR 0.31945f
C29320 a_31708_15271# a_32068_15368# 0.08717f
C29321 _452_.CLK a_43784_19369# 0.00262f
C29322 _452_.Q a_42376_22504# 0.00285f
C29323 a_30588_23111# VPWR 0.31547f
C29324 _324_.B a_44028_22020# 0.02456f
C29325 _229_.I a_62503_28293# 0.0048f
C29326 _424_.A1 _422_.ZN 0.20933f
C29327 _260_.A1 _305_.A2 0.00223f
C29328 a_45596_2727# a_45956_2824# 0.08717f
C29329 _452_.Q _330_.A2 0.03227f
C29330 a_42996_18840# VPWR 0.38073f
C29331 a_28000_29480# a_28880_29167# 0.00306f
C29332 a_62084_17316# a_62172_17272# 0.28563f
C29333 a_67884_16839# a_67796_16936# 0.28563f
C29334 a_61948_26247# VPWR 0.31547f
C29335 a_66092_18407# a_66540_18407# 0.01255f
C29336 a_4604_25112# a_5052_25112# 0.01222f
C29337 a_21876_23588# a_22548_23588# 0.00347f
C29338 _474_.CLK a_54244_20452# 0.00906f
C29339 a_65308_9432# a_65308_8999# 0.05841f
C29340 _355_.C a_26556_27815# 0.04805f
C29341 a_1020_4295# a_932_4392# 0.28563f
C29342 _424_.B1 a_51618_22504# 0.0021f
C29343 a_2364_13703# a_2276_13800# 0.28563f
C29344 _319_.A3 a_37067_19001# 0.01204f
C29345 a_28820_20452# a_29268_20452# 0.01328f
C29346 a_27476_20452# a_27116_20408# 0.08717f
C29347 _274_.A2 _255_.ZN 0.00682f
C29348 a_63428_18504# a_63428_17316# 0.05841f
C29349 a_3708_16839# a_3620_16936# 0.28563f
C29350 _457_.D a_24452_24776# 0.0023f
C29351 _296_.ZN _284_.ZN 1.84274f
C29352 _419_.Z a_46476_20937# 0.00102f
C29353 a_20284_1592# VPWR 0.3289f
C29354 a_35964_1592# a_36100_1256# 0.00168f
C29355 a_63652_12612# a_63292_12568# 0.08707f
C29356 a_66788_12612# a_67236_12612# 0.01328f
C29357 _324_.C a_49740_29383# 0.01666f
C29358 _437_.A1 _435_.A3 0.48107f
C29359 _475_.D VPWR 0.22379f
C29360 a_66428_15271# a_66788_15368# 0.08674f
C29361 a_50100_12232# a_50188_10567# 0.00151f
C29362 _304_.A1 a_38325_22804# 0.00597f
C29363 a_63764_12232# a_63740_11000# 0.0016f
C29364 a_41028_1636# a_40668_1592# 0.08707f
C29365 _304_.B a_44500_25156# 0.00258f
C29366 _281_.ZN _384_.A1 0.03932f
C29367 ui_in[5] VGND 0.04589f
C29368 ui_in[6] VGND 0.04633f
C29369 uio_in[2] VGND 0.04602f
C29370 uio_in[3] VGND 0.04598f
C29371 uio_in[4] VGND 0.04619f
C29372 uio_in[5] VGND 0.0462f
C29373 uio_in[6] VGND 0.04304f
C29374 uio_in[7] VGND 0.04658f
C29375 clk VGND 12.05168f
C29376 uo_out[6] VGND 1.78871f
C29377 uo_out[7] VGND 2.59555f
C29378 uo_out[3] VGND 1.81285f
C29379 uo_out[1] VGND 2.34677f
C29380 uio_out[7] VGND 1.69421f
C29381 rst_n VGND 0.80411f
C29382 uo_out[2] VGND 1.69239f
C29383 uo_out[4] VGND 1.6289f
C29384 uio_out[4] VGND 0.52525f
C29385 ena VGND 0.87945f
C29386 ui_in[0] VGND 0.70478f
C29387 ui_in[1] VGND 0.68751f
C29388 ui_in[2] VGND 0.78272f
C29389 ui_in[3] VGND 1.16701f
C29390 ui_in[4] VGND 0.8807f
C29391 ui_in[7] VGND 0.77509f
C29392 uo_out[0] VGND 1.58799f
C29393 uo_out[5] VGND 1.54476f
C29394 uio_in[0] VGND 0.88184f
C29395 uio_in[1] VGND 0.67151f
C29396 uio_out[0] VGND 0.48365f
C29397 uio_out[1] VGND 0.4564f
C29398 uio_out[2] VGND 0.37292f
C29399 uio_out[3] VGND 0.41884f
C29400 uio_oe[0] VGND 0.41849f
C29401 uio_out[6] VGND 1.78903f
C29402 uio_oe[1] VGND 0.41336f
C29403 uio_oe[2] VGND 0.4453f
C29404 uio_oe[3] VGND 0.58755f
C29405 uio_oe[4] VGND 0.23781f
C29406 uio_oe[5] VGND 0.23032f
C29407 uio_oe[6] VGND 0.34027f
C29408 uio_oe[7] VGND 0.31045f
C29409 uio_out[5] VGND 2.68711f
C29410 VPWR VGND 2.38637p
C29411 a_67908_1256# VGND 0.49509f
C29412 a_67460_1256# VGND 0.49004f
C29413 a_67012_1256# VGND 0.48947f
C29414 a_66564_1256# VGND 0.51466f
C29415 a_66116_1256# VGND 0.48299f
C29416 a_65668_1256# VGND 0.49231f
C29417 a_64996_1256# VGND 0.47896f
C29418 a_64548_1256# VGND 0.47513f
C29419 a_64100_1256# VGND 0.47513f
C29420 a_63652_1256# VGND 0.47513f
C29421 a_63204_1256# VGND 0.47513f
C29422 a_62756_1256# VGND 0.47513f
C29423 a_62308_1256# VGND 0.47513f
C29424 a_61860_1256# VGND 0.48718f
C29425 a_61188_1256# VGND 0.47896f
C29426 a_60740_1256# VGND 0.47547f
C29427 a_60292_1256# VGND 0.47833f
C29428 a_59844_1256# VGND 0.48007f
C29429 a_59396_1256# VGND 0.48274f
C29430 a_58948_1256# VGND 0.51179f
C29431 a_58500_1256# VGND 0.48297f
C29432 a_58052_1256# VGND 0.48718f
C29433 a_57380_1256# VGND 0.47896f
C29434 a_56932_1256# VGND 0.47513f
C29435 a_56484_1256# VGND 0.47513f
C29436 a_56036_1256# VGND 0.47513f
C29437 a_55588_1256# VGND 0.47513f
C29438 a_55140_1256# VGND 0.47513f
C29439 a_54692_1256# VGND 0.47513f
C29440 a_54244_1256# VGND 0.48718f
C29441 a_53572_1256# VGND 0.47896f
C29442 a_53124_1256# VGND 0.47513f
C29443 a_52676_1256# VGND 0.47789f
C29444 a_52228_1256# VGND 0.47937f
C29445 a_51780_1256# VGND 0.48155f
C29446 a_51332_1256# VGND 0.49357f
C29447 a_50884_1256# VGND 0.49313f
C29448 a_50436_1256# VGND 0.48718f
C29449 a_49764_1256# VGND 0.47896f
C29450 a_49316_1256# VGND 0.47513f
C29451 a_48868_1256# VGND 0.47513f
C29452 a_48420_1256# VGND 0.47513f
C29453 a_47972_1256# VGND 0.47513f
C29454 a_47524_1256# VGND 0.47513f
C29455 a_47076_1256# VGND 0.47513f
C29456 a_46628_1256# VGND 0.48718f
C29457 a_45956_1256# VGND 0.47896f
C29458 a_45508_1256# VGND 0.47513f
C29459 a_45060_1256# VGND 0.47668f
C29460 a_44612_1256# VGND 0.47876f
C29461 a_44164_1256# VGND 0.48072f
C29462 a_43716_1256# VGND 0.4837f
C29463 a_43268_1256# VGND 0.51289f
C29464 a_42820_1256# VGND 0.49029f
C29465 a_42148_1256# VGND 0.47896f
C29466 a_41700_1256# VGND 0.47513f
C29467 a_41252_1256# VGND 0.47513f
C29468 a_40804_1256# VGND 0.47513f
C29469 a_40356_1256# VGND 0.47513f
C29470 a_39908_1256# VGND 0.47513f
C29471 a_39460_1256# VGND 0.47513f
C29472 a_39012_1256# VGND 0.48718f
C29473 a_38340_1256# VGND 0.47896f
C29474 a_37892_1256# VGND 0.47513f
C29475 a_37444_1256# VGND 0.47519f
C29476 a_36996_1256# VGND 0.47826f
C29477 a_36548_1256# VGND 0.47995f
C29478 a_36100_1256# VGND 0.48255f
C29479 a_35652_1256# VGND 0.50895f
C29480 a_35204_1256# VGND 0.49545f
C29481 a_34532_1256# VGND 0.47896f
C29482 a_34084_1256# VGND 0.47513f
C29483 a_33636_1256# VGND 0.47513f
C29484 a_33188_1256# VGND 0.47513f
C29485 a_32740_1256# VGND 0.47513f
C29486 a_32292_1256# VGND 0.47513f
C29487 a_31844_1256# VGND 0.47513f
C29488 a_31396_1256# VGND 0.48718f
C29489 a_30724_1256# VGND 0.47896f
C29490 a_30276_1256# VGND 0.47513f
C29491 a_29828_1256# VGND 0.47513f
C29492 a_29380_1256# VGND 0.47783f
C29493 a_28932_1256# VGND 0.47926f
C29494 a_28484_1256# VGND 0.4814f
C29495 a_28036_1256# VGND 0.48952f
C29496 a_27588_1256# VGND 0.50812f
C29497 a_26916_1256# VGND 0.47896f
C29498 a_26468_1256# VGND 0.47513f
C29499 a_26020_1256# VGND 0.47513f
C29500 a_25572_1256# VGND 0.47513f
C29501 a_25124_1256# VGND 0.47513f
C29502 a_24676_1256# VGND 0.47513f
C29503 a_24228_1256# VGND 0.47513f
C29504 a_23780_1256# VGND 0.48718f
C29505 a_23108_1256# VGND 0.47896f
C29506 a_22660_1256# VGND 0.47513f
C29507 a_22212_1256# VGND 0.47513f
C29508 a_21764_1256# VGND 0.47646f
C29509 a_21316_1256# VGND 0.47868f
C29510 a_20868_1256# VGND 0.48059f
C29511 a_20420_1256# VGND 0.48353f
C29512 a_19972_1256# VGND 0.52905f
C29513 a_19300_1256# VGND 0.47902f
C29514 a_18852_1256# VGND 0.47513f
C29515 a_18404_1256# VGND 0.47513f
C29516 a_17956_1256# VGND 0.47513f
C29517 a_17508_1256# VGND 0.47513f
C29518 a_17060_1256# VGND 0.47513f
C29519 a_16612_1256# VGND 0.47513f
C29520 a_16164_1256# VGND 0.48718f
C29521 a_15492_1256# VGND 0.47896f
C29522 a_15044_1256# VGND 0.47513f
C29523 a_14596_1256# VGND 0.47513f
C29524 a_14148_1256# VGND 0.47513f
C29525 a_13700_1256# VGND 0.47818f
C29526 a_13252_1256# VGND 0.47983f
C29527 a_12804_1256# VGND 0.48236f
C29528 a_12356_1256# VGND 0.51868f
C29529 a_11684_1256# VGND 0.48152f
C29530 a_11236_1256# VGND 0.47513f
C29531 a_10788_1256# VGND 0.47513f
C29532 a_10340_1256# VGND 0.47513f
C29533 a_9892_1256# VGND 0.47513f
C29534 a_9444_1256# VGND 0.47513f
C29535 a_8996_1256# VGND 0.47513f
C29536 a_8548_1256# VGND 0.48718f
C29537 a_7876_1256# VGND 0.47896f
C29538 a_7428_1256# VGND 0.47513f
C29539 a_6980_1256# VGND 0.47513f
C29540 a_6532_1256# VGND 0.47513f
C29541 a_6084_1256# VGND 0.47765f
C29542 a_5636_1256# VGND 0.47916f
C29543 a_5188_1256# VGND 0.48126f
C29544 a_4740_1256# VGND 0.49929f
C29545 a_4068_1256# VGND 0.48653f
C29546 a_3620_1256# VGND 0.47513f
C29547 a_3172_1256# VGND 0.47513f
C29548 a_2724_1256# VGND 0.47513f
C29549 a_2276_1256# VGND 0.47513f
C29550 a_1828_1256# VGND 0.47513f
C29551 a_1380_1256# VGND 0.47513f
C29552 a_932_1256# VGND 0.50325f
C29553 a_67996_1159# VGND 0.2929f
C29554 a_67548_1159# VGND 0.29477f
C29555 a_67100_1159# VGND 0.29674f
C29556 a_66652_1159# VGND 0.3353f
C29557 a_66204_1159# VGND 0.29388f
C29558 a_65756_1159# VGND 0.29054f
C29559 a_65084_1159# VGND 0.28628f
C29560 a_64636_1159# VGND 0.2812f
C29561 a_64188_1159# VGND 0.2812f
C29562 a_63740_1159# VGND 0.2812f
C29563 a_63292_1159# VGND 0.2844f
C29564 a_62844_1159# VGND 0.28448f
C29565 a_62396_1159# VGND 0.28447f
C29566 a_61948_1159# VGND 0.28818f
C29567 a_61276_1159# VGND 0.28628f
C29568 a_60828_1159# VGND 0.2812f
C29569 a_60380_1159# VGND 0.28446f
C29570 a_59932_1159# VGND 0.28611f
C29571 a_59484_1159# VGND 0.28836f
C29572 a_59036_1159# VGND 0.30606f
C29573 a_58588_1159# VGND 0.29305f
C29574 a_58140_1159# VGND 0.28492f
C29575 a_57468_1159# VGND 0.28954f
C29576 a_57020_1159# VGND 0.28447f
C29577 a_56572_1159# VGND 0.28447f
C29578 a_56124_1159# VGND 0.28447f
C29579 a_55676_1159# VGND 0.28456f
C29580 a_55228_1159# VGND 0.2812f
C29581 a_54780_1159# VGND 0.2812f
C29582 a_54332_1159# VGND 0.28492f
C29583 a_53660_1159# VGND 0.28954f
C29584 a_53212_1159# VGND 0.28447f
C29585 a_52764_1159# VGND 0.28687f
C29586 a_52316_1159# VGND 0.28871f
C29587 a_51868_1159# VGND 0.2908f
C29588 a_51420_1159# VGND 0.29362f
C29589 a_50972_1159# VGND 0.31953f
C29590 a_50524_1159# VGND 0.29064f
C29591 a_49852_1159# VGND 0.28628f
C29592 a_49404_1159# VGND 0.2812f
C29593 a_48956_1159# VGND 0.2812f
C29594 a_48508_1159# VGND 0.2812f
C29595 a_48060_1159# VGND 0.2812f
C29596 a_47612_1159# VGND 0.2844f
C29597 a_47164_1159# VGND 0.28448f
C29598 a_46716_1159# VGND 0.28818f
C29599 a_46044_1159# VGND 0.28628f
C29600 a_45596_1159# VGND 0.2812f
C29601 a_45148_1159# VGND 0.28198f
C29602 a_44700_1159# VGND 0.28487f
C29603 a_44252_1159# VGND 0.28673f
C29604 a_43804_1159# VGND 0.28905f
C29605 a_43356_1159# VGND 0.32338f
C29606 a_42908_1159# VGND 0.29236f
C29607 a_42236_1159# VGND 0.28954f
C29608 a_41788_1159# VGND 0.28447f
C29609 a_41340_1159# VGND 0.28447f
C29610 a_40892_1159# VGND 0.28447f
C29611 a_40444_1159# VGND 0.28447f
C29612 a_39996_1159# VGND 0.28456f
C29613 a_39548_1159# VGND 0.2812f
C29614 a_39100_1159# VGND 0.28492f
C29615 a_38428_1159# VGND 0.28954f
C29616 a_37980_1159# VGND 0.28447f
C29617 a_37532_1159# VGND 0.28447f
C29618 a_37084_1159# VGND 0.28765f
C29619 a_36636_1159# VGND 0.28926f
C29620 a_36188_1159# VGND 0.29149f
C29621 a_35740_1159# VGND 0.30728f
C29622 a_35292_1159# VGND 0.30392f
C29623 a_34620_1159# VGND 0.28628f
C29624 a_34172_1159# VGND 0.2812f
C29625 a_33724_1159# VGND 0.2812f
C29626 a_33276_1159# VGND 0.2812f
C29627 a_32828_1159# VGND 0.2812f
C29628 a_32380_1159# VGND 0.2812f
C29629 a_31932_1159# VGND 0.2844f
C29630 a_31484_1159# VGND 0.28819f
C29631 a_30812_1159# VGND 0.28628f
C29632 a_30364_1159# VGND 0.2812f
C29633 a_29916_1159# VGND 0.2812f
C29634 a_29468_1159# VGND 0.28338f
C29635 a_29020_1159# VGND 0.28534f
C29636 a_28572_1159# VGND 0.2874f
C29637 a_28124_1159# VGND 0.29011f
C29638 a_27676_1159# VGND 0.3222f
C29639 a_27004_1159# VGND 0.28969f
C29640 a_26556_1159# VGND 0.28447f
C29641 a_26108_1159# VGND 0.28447f
C29642 a_25660_1159# VGND 0.28447f
C29643 a_25212_1159# VGND 0.28447f
C29644 a_24764_1159# VGND 0.28447f
C29645 a_24316_1159# VGND 0.28456f
C29646 a_23868_1159# VGND 0.28492f
C29647 a_23196_1159# VGND 0.28954f
C29648 a_22748_1159# VGND 0.28447f
C29649 a_22300_1159# VGND 0.28447f
C29650 a_21852_1159# VGND 0.28498f
C29651 a_21404_1159# VGND 0.28805f
C29652 a_20956_1159# VGND 0.28987f
C29653 a_20508_1159# VGND 0.29218f
C29654 a_20060_1159# VGND 0.32748f
C29655 a_19388_1159# VGND 0.28756f
C29656 a_18940_1159# VGND 0.2812f
C29657 a_18492_1159# VGND 0.2812f
C29658 a_18044_1159# VGND 0.2812f
C29659 a_17596_1159# VGND 0.2812f
C29660 a_17148_1159# VGND 0.2812f
C29661 a_16700_1159# VGND 0.2812f
C29662 a_16252_1159# VGND 0.28811f
C29663 a_15580_1159# VGND 0.28628f
C29664 a_15132_1159# VGND 0.2812f
C29665 a_14684_1159# VGND 0.2812f
C29666 a_14236_1159# VGND 0.2812f
C29667 a_13788_1159# VGND 0.28431f
C29668 a_13340_1159# VGND 0.28588f
C29669 a_12892_1159# VGND 0.28809f
C29670 a_12444_1159# VGND 0.30384f
C29671 a_11772_1159# VGND 0.29666f
C29672 a_11324_1159# VGND 0.28447f
C29673 a_10876_1159# VGND 0.28447f
C29674 a_10428_1159# VGND 0.28447f
C29675 a_9980_1159# VGND 0.28447f
C29676 a_9532_1159# VGND 0.28447f
C29677 a_9084_1159# VGND 0.28447f
C29678 a_8636_1159# VGND 0.28827f
C29679 a_7964_1159# VGND 0.28955f
C29680 a_7516_1159# VGND 0.28447f
C29681 a_7068_1159# VGND 0.28447f
C29682 a_6620_1159# VGND 0.28447f
C29683 a_6172_1159# VGND 0.28639f
C29684 a_5724_1159# VGND 0.28851f
C29685 a_5276_1159# VGND 0.29053f
C29686 a_4828_1159# VGND 0.29748f
C29687 a_4156_1159# VGND 0.2987f
C29688 a_3708_1159# VGND 0.2812f
C29689 a_3260_1159# VGND 0.2812f
C29690 a_2812_1159# VGND 0.2812f
C29691 a_2364_1159# VGND 0.2812f
C29692 a_1916_1159# VGND 0.2812f
C29693 a_1468_1159# VGND 0.2812f
C29694 a_1020_1159# VGND 0.29134f
C29695 a_67772_1592# VGND 0.28907f
C29696 a_67324_1592# VGND 0.29953f
C29697 a_66876_1592# VGND 0.30917f
C29698 a_66428_1592# VGND 0.31142f
C29699 a_65980_1592# VGND 0.28814f
C29700 a_65532_1592# VGND 0.28816f
C29701 a_65084_1592# VGND 0.2812f
C29702 a_64636_1592# VGND 0.2812f
C29703 a_64188_1592# VGND 0.2812f
C29704 a_63740_1592# VGND 0.28492f
C29705 a_67684_1636# VGND 0.49163f
C29706 a_67236_1636# VGND 0.48755f
C29707 a_66788_1636# VGND 0.50141f
C29708 a_66340_1636# VGND 0.48002f
C29709 a_65892_1636# VGND 0.47122f
C29710 a_65444_1636# VGND 0.47187f
C29711 a_64996_1636# VGND 0.43828f
C29712 a_64548_1636# VGND 0.43828f
C29713 a_64100_1636# VGND 0.43828f
C29714 a_63652_1636# VGND 0.45034f
C29715 a_63068_1592# VGND 0.29459f
C29716 a_62620_1592# VGND 0.2927f
C29717 a_62172_1592# VGND 0.28922f
C29718 a_61724_1592# VGND 0.28932f
C29719 a_61276_1592# VGND 0.28236f
C29720 a_60828_1592# VGND 0.28236f
C29721 a_60380_1592# VGND 0.28562f
C29722 a_59932_1592# VGND 0.28727f
C29723 a_59484_1592# VGND 0.28952f
C29724 a_59036_1592# VGND 0.30721f
C29725 a_58588_1592# VGND 0.29418f
C29726 a_58140_1592# VGND 0.28236f
C29727 a_57692_1592# VGND 0.28916f
C29728 a_57244_1592# VGND 0.28922f
C29729 a_56796_1592# VGND 0.28922f
C29730 a_56348_1592# VGND 0.28922f
C29731 a_55900_1592# VGND 0.29272f
C29732 a_62980_1636# VGND 0.48791f
C29733 a_62532_1636# VGND 0.474f
C29734 a_62084_1636# VGND 0.474f
C29735 a_61636_1636# VGND 0.47466f
C29736 a_61188_1636# VGND 0.44029f
C29737 a_60740_1636# VGND 0.44063f
C29738 a_60292_1636# VGND 0.44349f
C29739 a_59844_1636# VGND 0.44523f
C29740 a_59396_1636# VGND 0.4479f
C29741 a_58948_1636# VGND 0.47694f
C29742 a_58500_1636# VGND 0.44813f
C29743 a_58052_1636# VGND 0.44029f
C29744 a_57604_1636# VGND 0.47343f
C29745 a_57156_1636# VGND 0.474f
C29746 a_56708_1636# VGND 0.474f
C29747 a_56260_1636# VGND 0.474f
C29748 a_55812_1636# VGND 0.48596f
C29749 a_55228_1592# VGND 0.28772f
C29750 a_54780_1592# VGND 0.28584f
C29751 a_54332_1592# VGND 0.28236f
C29752 a_53884_1592# VGND 0.28916f
C29753 a_53436_1592# VGND 0.28922f
C29754 a_52988_1592# VGND 0.28934f
C29755 a_52540_1592# VGND 0.29268f
C29756 a_52092_1592# VGND 0.29444f
C29757 a_51644_1592# VGND 0.29671f
C29758 a_51196_1592# VGND 0.32395f
C29759 a_50748_1592# VGND 0.29908f
C29760 a_50300_1592# VGND 0.28932f
C29761 a_49852_1592# VGND 0.28236f
C29762 a_49404_1592# VGND 0.28236f
C29763 a_48956_1592# VGND 0.28236f
C29764 a_48508_1592# VGND 0.28236f
C29765 a_48060_1592# VGND 0.28586f
C29766 a_55140_1636# VGND 0.4542f
C29767 a_54692_1636# VGND 0.44029f
C29768 a_54244_1636# VGND 0.44029f
C29769 a_53796_1636# VGND 0.47343f
C29770 a_53348_1636# VGND 0.474f
C29771 a_52900_1636# VGND 0.475f
C29772 a_52452_1636# VGND 0.47742f
C29773 a_52004_1636# VGND 0.47926f
C29774 a_51556_1636# VGND 0.48208f
C29775 a_51108_1636# VGND 0.52042f
C29776 a_50660_1636# VGND 0.47882f
C29777 a_50212_1636# VGND 0.47466f
C29778 a_49764_1636# VGND 0.44029f
C29779 a_49316_1636# VGND 0.44029f
C29780 a_48868_1636# VGND 0.44029f
C29781 a_48420_1636# VGND 0.44029f
C29782 a_47972_1636# VGND 0.45225f
C29783 a_47388_1592# VGND 0.29459f
C29784 a_46940_1592# VGND 0.2927f
C29785 a_46492_1592# VGND 0.28932f
C29786 a_46044_1592# VGND 0.28236f
C29787 a_45596_1592# VGND 0.28236f
C29788 a_45148_1592# VGND 0.28314f
C29789 a_44700_1592# VGND 0.28603f
C29790 a_44252_1592# VGND 0.28789f
C29791 a_43804_1592# VGND 0.29021f
C29792 a_43356_1592# VGND 0.32454f
C29793 a_42908_1592# VGND 0.28978f
C29794 a_42460_1592# VGND 0.28916f
C29795 a_42012_1592# VGND 0.28922f
C29796 a_41564_1592# VGND 0.28922f
C29797 a_41116_1592# VGND 0.28922f
C29798 a_40668_1592# VGND 0.28922f
C29799 a_40220_1592# VGND 0.29272f
C29800 a_47300_1636# VGND 0.48791f
C29801 a_46852_1636# VGND 0.474f
C29802 a_46404_1636# VGND 0.47466f
C29803 a_45956_1636# VGND 0.44029f
C29804 a_45508_1636# VGND 0.44029f
C29805 a_45060_1636# VGND 0.44184f
C29806 a_44612_1636# VGND 0.44392f
C29807 a_44164_1636# VGND 0.44588f
C29808 a_43716_1636# VGND 0.44886f
C29809 a_43268_1636# VGND 0.47805f
C29810 a_42820_1636# VGND 0.44339f
C29811 a_42372_1636# VGND 0.47343f
C29812 a_41924_1636# VGND 0.474f
C29813 a_41476_1636# VGND 0.474f
C29814 a_41028_1636# VGND 0.474f
C29815 a_40580_1636# VGND 0.474f
C29816 a_40132_1636# VGND 0.48596f
C29817 a_39548_1592# VGND 0.28772f
C29818 a_39100_1592# VGND 0.28584f
C29819 a_38652_1592# VGND 0.28916f
C29820 a_38204_1592# VGND 0.28922f
C29821 a_37756_1592# VGND 0.28922f
C29822 a_37308_1592# VGND 0.2907f
C29823 a_36860_1592# VGND 0.29312f
C29824 a_36412_1592# VGND 0.29508f
C29825 a_35964_1592# VGND 0.29764f
C29826 a_35516_1592# VGND 0.33528f
C29827 a_35068_1592# VGND 0.29451f
C29828 a_34620_1592# VGND 0.28236f
C29829 a_34172_1592# VGND 0.28236f
C29830 a_33724_1592# VGND 0.28236f
C29831 a_33276_1592# VGND 0.28236f
C29832 a_32828_1592# VGND 0.28236f
C29833 a_32380_1592# VGND 0.28586f
C29834 a_39460_1636# VGND 0.4542f
C29835 a_39012_1636# VGND 0.44029f
C29836 a_38564_1636# VGND 0.47343f
C29837 a_38116_1636# VGND 0.474f
C29838 a_37668_1636# VGND 0.474f
C29839 a_37220_1636# VGND 0.47615f
C29840 a_36772_1636# VGND 0.47788f
C29841 a_36324_1636# VGND 0.47993f
C29842 a_35876_1636# VGND 0.48363f
C29843 a_35428_1636# VGND 0.50558f
C29844 a_34980_1636# VGND 0.47626f
C29845 a_34532_1636# VGND 0.44029f
C29846 a_34084_1636# VGND 0.44029f
C29847 a_33636_1636# VGND 0.44029f
C29848 a_33188_1636# VGND 0.44029f
C29849 a_32740_1636# VGND 0.44029f
C29850 a_32292_1636# VGND 0.45225f
C29851 a_31708_1592# VGND 0.29459f
C29852 a_31260_1592# VGND 0.2928f
C29853 a_30812_1592# VGND 0.28236f
C29854 a_30364_1592# VGND 0.28236f
C29855 a_29916_1592# VGND 0.28236f
C29856 a_29468_1592# VGND 0.28454f
C29857 a_29020_1592# VGND 0.28651f
C29858 a_28572_1592# VGND 0.28856f
C29859 a_28124_1592# VGND 0.29126f
C29860 a_27676_1592# VGND 0.31964f
C29861 a_27228_1592# VGND 0.29225f
C29862 a_26780_1592# VGND 0.28922f
C29863 a_26332_1592# VGND 0.28922f
C29864 a_25884_1592# VGND 0.28922f
C29865 a_25436_1592# VGND 0.28922f
C29866 a_24988_1592# VGND 0.28922f
C29867 a_24540_1592# VGND 0.29272f
C29868 a_31620_1636# VGND 0.48791f
C29869 a_31172_1636# VGND 0.47466f
C29870 a_30724_1636# VGND 0.44029f
C29871 a_30276_1636# VGND 0.44029f
C29872 a_29828_1636# VGND 0.44029f
C29873 a_29380_1636# VGND 0.44299f
C29874 a_28932_1636# VGND 0.44442f
C29875 a_28484_1636# VGND 0.44656f
C29876 a_28036_1636# VGND 0.45468f
C29877 a_27588_1636# VGND 0.46123f
C29878 a_27140_1636# VGND 0.47363f
C29879 a_26692_1636# VGND 0.474f
C29880 a_26244_1636# VGND 0.474f
C29881 a_25796_1636# VGND 0.474f
C29882 a_25348_1636# VGND 0.474f
C29883 a_24900_1636# VGND 0.474f
C29884 a_24452_1636# VGND 0.48596f
C29885 a_23868_1592# VGND 0.28772f
C29886 a_23420_1592# VGND 0.29264f
C29887 a_22972_1592# VGND 0.28922f
C29888 a_22524_1592# VGND 0.28922f
C29889 a_22076_1592# VGND 0.28922f
C29890 a_21628_1592# VGND 0.2921f
C29891 a_21180_1592# VGND 0.29363f
C29892 a_20732_1592# VGND 0.29577f
C29893 a_20284_1592# VGND 0.30012f
C29894 a_19836_1592# VGND 0.31932f
C29895 a_19388_1592# VGND 0.28342f
C29896 a_18940_1592# VGND 0.28236f
C29897 a_18492_1592# VGND 0.28236f
C29898 a_18044_1592# VGND 0.28236f
C29899 a_17596_1592# VGND 0.28236f
C29900 a_17148_1592# VGND 0.28236f
C29901 a_16700_1592# VGND 0.28586f
C29902 a_23780_1636# VGND 0.4542f
C29903 a_23332_1636# VGND 0.47343f
C29904 a_22884_1636# VGND 0.474f
C29905 a_22436_1636# VGND 0.474f
C29906 a_21988_1636# VGND 0.474f
C29907 a_21540_1636# VGND 0.47687f
C29908 a_21092_1636# VGND 0.47841f
C29909 a_20644_1636# VGND 0.48073f
C29910 a_20196_1636# VGND 0.49798f
C29911 a_19748_1636# VGND 0.48872f
C29912 a_19300_1636# VGND 0.44029f
C29913 a_18852_1636# VGND 0.44029f
C29914 a_18404_1636# VGND 0.44029f
C29915 a_17956_1636# VGND 0.44029f
C29916 a_17508_1636# VGND 0.44029f
C29917 a_17060_1636# VGND 0.44029f
C29918 a_16612_1636# VGND 0.45225f
C29919 a_16028_1592# VGND 0.29468f
C29920 a_15580_1592# VGND 0.28584f
C29921 a_15132_1592# VGND 0.28236f
C29922 a_14684_1592# VGND 0.28236f
C29923 a_14236_1592# VGND 0.28236f
C29924 a_13788_1592# VGND 0.28547f
C29925 a_13340_1592# VGND 0.28704f
C29926 a_12892_1592# VGND 0.28925f
C29927 a_12444_1592# VGND 0.30115f
C29928 a_11996_1592# VGND 0.31019f
C29929 a_11548_1592# VGND 0.28926f
C29930 a_11100_1592# VGND 0.28922f
C29931 a_10652_1592# VGND 0.28922f
C29932 a_10204_1592# VGND 0.28922f
C29933 a_9756_1592# VGND 0.28922f
C29934 a_9308_1592# VGND 0.28922f
C29935 a_8860_1592# VGND 0.29272f
C29936 a_15940_1636# VGND 0.48857f
C29937 a_15492_1636# VGND 0.44029f
C29938 a_15044_1636# VGND 0.44029f
C29939 a_14596_1636# VGND 0.44029f
C29940 a_14148_1636# VGND 0.44029f
C29941 a_13700_1636# VGND 0.44334f
C29942 a_13252_1636# VGND 0.44499f
C29943 a_12804_1636# VGND 0.44752f
C29944 a_12356_1636# VGND 0.47129f
C29945 a_11908_1636# VGND 0.48201f
C29946 a_11460_1636# VGND 0.474f
C29947 a_11012_1636# VGND 0.474f
C29948 a_10564_1636# VGND 0.474f
C29949 a_10116_1636# VGND 0.474f
C29950 a_9668_1636# VGND 0.474f
C29951 a_9220_1636# VGND 0.474f
C29952 a_8772_1636# VGND 0.48596f
C29953 a_8188_1592# VGND 0.29452f
C29954 a_7740_1592# VGND 0.2927f
C29955 a_7292_1592# VGND 0.28922f
C29956 a_6844_1592# VGND 0.28922f
C29957 a_6396_1592# VGND 0.28922f
C29958 a_5948_1592# VGND 0.29252f
C29959 a_5500_1592# VGND 0.2942f
C29960 a_5052_1592# VGND 0.29645f
C29961 a_4604_1592# VGND 0.31757f
C29962 a_4156_1592# VGND 0.29327f
C29963 a_3708_1592# VGND 0.28236f
C29964 a_3260_1592# VGND 0.28236f
C29965 a_2812_1592# VGND 0.28236f
C29966 a_2364_1592# VGND 0.28236f
C29967 a_1916_1592# VGND 0.28236f
C29968 a_1468_1592# VGND 0.28236f
C29969 a_1020_1592# VGND 0.29228f
C29970 a_8100_1636# VGND 0.48734f
C29971 a_7652_1636# VGND 0.474f
C29972 a_7204_1636# VGND 0.474f
C29973 a_6756_1636# VGND 0.474f
C29974 a_6308_1636# VGND 0.47451f
C29975 a_5860_1636# VGND 0.47692f
C29976 a_5412_1636# VGND 0.47817f
C29977 a_4964_1636# VGND 0.47846f
C29978 a_4516_1636# VGND 0.51132f
C29979 a_4068_1636# VGND 0.44738f
C29980 a_3620_1636# VGND 0.44029f
C29981 a_3172_1636# VGND 0.44029f
C29982 a_2724_1636# VGND 0.44029f
C29983 a_2276_1636# VGND 0.44029f
C29984 a_1828_1636# VGND 0.44029f
C29985 a_1380_1636# VGND 0.44029f
C29986 a_932_1636# VGND 0.46832f
C29987 a_67908_2824# VGND 0.48748f
C29988 a_67460_2824# VGND 0.4837f
C29989 a_67012_2824# VGND 0.48313f
C29990 a_66564_2824# VGND 0.50992f
C29991 a_66116_2824# VGND 0.4766f
C29992 a_65668_2824# VGND 0.48592f
C29993 a_64996_2824# VGND 0.44211f
C29994 a_64548_2824# VGND 0.43828f
C29995 a_64100_2824# VGND 0.43828f
C29996 a_63652_2824# VGND 0.43828f
C29997 a_63204_2824# VGND 0.46817f
C29998 a_62756_2824# VGND 0.4688f
C29999 a_62308_2824# VGND 0.46875f
C30000 a_61860_2824# VGND 0.48081f
C30001 a_61188_2824# VGND 0.44211f
C30002 a_60740_2824# VGND 0.43862f
C30003 a_60292_2824# VGND 0.44149f
C30004 a_59844_2824# VGND 0.44322f
C30005 a_59396_2824# VGND 0.44589f
C30006 a_58948_2824# VGND 0.47297f
C30007 a_58500_2824# VGND 0.44612f
C30008 a_58052_2824# VGND 0.45034f
C30009 a_57380_2824# VGND 0.47258f
C30010 a_56932_2824# VGND 0.46875f
C30011 a_56484_2824# VGND 0.46875f
C30012 a_56036_2824# VGND 0.46875f
C30013 a_55588_2824# VGND 0.46941f
C30014 a_55140_2824# VGND 0.43828f
C30015 a_54692_2824# VGND 0.43828f
C30016 a_54244_2824# VGND 0.45034f
C30017 a_53572_2824# VGND 0.47258f
C30018 a_53124_2824# VGND 0.46875f
C30019 a_52676_2824# VGND 0.47152f
C30020 a_52228_2824# VGND 0.47299f
C30021 a_51780_2824# VGND 0.47518f
C30022 a_51332_2824# VGND 0.4865f
C30023 a_50884_2824# VGND 0.48692f
C30024 a_50436_2824# VGND 0.48081f
C30025 a_49764_2824# VGND 0.44211f
C30026 a_49316_2824# VGND 0.43828f
C30027 a_48868_2824# VGND 0.43828f
C30028 a_48420_2824# VGND 0.43828f
C30029 a_47972_2824# VGND 0.43828f
C30030 a_47524_2824# VGND 0.46817f
C30031 a_47076_2824# VGND 0.4688f
C30032 a_46628_2824# VGND 0.48081f
C30033 a_45956_2824# VGND 0.44211f
C30034 a_45508_2824# VGND 0.43828f
C30035 a_45060_2824# VGND 0.43984f
C30036 a_44612_2824# VGND 0.44192f
C30037 a_44164_2824# VGND 0.44387f
C30038 a_43716_2824# VGND 0.44685f
C30039 a_43268_2824# VGND 0.47417f
C30040 a_42820_2824# VGND 0.45344f
C30041 a_42148_2824# VGND 0.47258f
C30042 a_41700_2824# VGND 0.46875f
C30043 a_41252_2824# VGND 0.46875f
C30044 a_40804_2824# VGND 0.46875f
C30045 a_40356_2824# VGND 0.46875f
C30046 a_39908_2824# VGND 0.46941f
C30047 a_39460_2824# VGND 0.43828f
C30048 a_39012_2824# VGND 0.45034f
C30049 a_38340_2824# VGND 0.47258f
C30050 a_37892_2824# VGND 0.46875f
C30051 a_37444_2824# VGND 0.46881f
C30052 a_36996_2824# VGND 0.47188f
C30053 a_36548_2824# VGND 0.47357f
C30054 a_36100_2824# VGND 0.47617f
C30055 a_35652_2824# VGND 0.50177f
C30056 a_35204_2824# VGND 0.48908f
C30057 a_34532_2824# VGND 0.44211f
C30058 a_34084_2824# VGND 0.43828f
C30059 a_33636_2824# VGND 0.43828f
C30060 a_33188_2824# VGND 0.43828f
C30061 a_32740_2824# VGND 0.43828f
C30062 a_32292_2824# VGND 0.43828f
C30063 a_31844_2824# VGND 0.46817f
C30064 a_31396_2824# VGND 0.48085f
C30065 a_30724_2824# VGND 0.44211f
C30066 a_30276_2824# VGND 0.43828f
C30067 a_29828_2824# VGND 0.43828f
C30068 a_29380_2824# VGND 0.44098f
C30069 a_28932_2824# VGND 0.44241f
C30070 a_28484_2824# VGND 0.44455f
C30071 a_28036_2824# VGND 0.45229f
C30072 a_27588_2824# VGND 0.47055f
C30073 a_26916_2824# VGND 0.47258f
C30074 a_26468_2824# VGND 0.46875f
C30075 a_26020_2824# VGND 0.46875f
C30076 a_25572_2824# VGND 0.46875f
C30077 a_25124_2824# VGND 0.46875f
C30078 a_24676_2824# VGND 0.46875f
C30079 a_24228_2824# VGND 0.46941f
C30080 a_23780_2824# VGND 0.45034f
C30081 a_23108_2824# VGND 0.47258f
C30082 a_22660_2824# VGND 0.46875f
C30083 a_22212_2824# VGND 0.46875f
C30084 a_21764_2824# VGND 0.47008f
C30085 a_21316_2824# VGND 0.4723f
C30086 a_20868_2824# VGND 0.47421f
C30087 a_20420_2824# VGND 0.47716f
C30088 a_19972_2824# VGND 0.52209f
C30089 a_19300_2824# VGND 0.44218f
C30090 a_18852_2824# VGND 0.43828f
C30091 a_18404_2824# VGND 0.43828f
C30092 a_17956_2824# VGND 0.43828f
C30093 a_17508_2824# VGND 0.43828f
C30094 a_17060_2824# VGND 0.43828f
C30095 a_16612_2824# VGND 0.43828f
C30096 a_16164_2824# VGND 0.48023f
C30097 a_15492_2824# VGND 0.44211f
C30098 a_15044_2824# VGND 0.43828f
C30099 a_14596_2824# VGND 0.43828f
C30100 a_14148_2824# VGND 0.43828f
C30101 a_13700_2824# VGND 0.44133f
C30102 a_13252_2824# VGND 0.44298f
C30103 a_12804_2824# VGND 0.44551f
C30104 a_12356_2824# VGND 0.48022f
C30105 a_11684_2824# VGND 0.47514f
C30106 a_11236_2824# VGND 0.46875f
C30107 a_10788_2824# VGND 0.46875f
C30108 a_10340_2824# VGND 0.46875f
C30109 a_9892_2824# VGND 0.46875f
C30110 a_9444_2824# VGND 0.46875f
C30111 a_8996_2824# VGND 0.46875f
C30112 a_8548_2824# VGND 0.48147f
C30113 a_7876_2824# VGND 0.47263f
C30114 a_7428_2824# VGND 0.46875f
C30115 a_6980_2824# VGND 0.46875f
C30116 a_6532_2824# VGND 0.46875f
C30117 a_6084_2824# VGND 0.47127f
C30118 a_5636_2824# VGND 0.47278f
C30119 a_5188_2824# VGND 0.47489f
C30120 a_4740_2824# VGND 0.49292f
C30121 a_4068_2824# VGND 0.44968f
C30122 a_3620_2824# VGND 0.43828f
C30123 a_3172_2824# VGND 0.43828f
C30124 a_2724_2824# VGND 0.43828f
C30125 a_2276_2824# VGND 0.43828f
C30126 a_1828_2824# VGND 0.43828f
C30127 a_1380_2824# VGND 0.43828f
C30128 a_932_2824# VGND 0.4664f
C30129 a_67996_2727# VGND 0.2898f
C30130 a_67548_2727# VGND 0.2915f
C30131 a_67100_2727# VGND 0.29347f
C30132 a_66652_2727# VGND 0.33039f
C30133 a_66204_2727# VGND 0.29061f
C30134 a_65756_2727# VGND 0.28728f
C30135 a_65084_2727# VGND 0.29253f
C30136 a_64636_2727# VGND 0.28746f
C30137 a_64188_2727# VGND 0.28757f
C30138 a_63740_2727# VGND 0.30341f
C30139 a_63292_2727# VGND 0.30341f
C30140 a_62844_2727# VGND 0.30341f
C30141 a_62396_2727# VGND 0.30341f
C30142 a_61948_2727# VGND 0.30712f
C30143 a_61276_2727# VGND 0.30848f
C30144 a_60828_2727# VGND 0.30341f
C30145 a_60380_2727# VGND 0.30666f
C30146 a_59932_2727# VGND 0.30832f
C30147 a_59484_2727# VGND 0.31056f
C30148 a_59036_2727# VGND 0.32954f
C30149 a_58588_2727# VGND 0.31523f
C30150 a_58140_2727# VGND 0.30712f
C30151 a_57468_2727# VGND 0.30848f
C30152 a_57020_2727# VGND 0.30341f
C30153 a_56572_2727# VGND 0.30341f
C30154 a_56124_2727# VGND 0.30341f
C30155 a_55676_2727# VGND 0.30341f
C30156 a_55228_2727# VGND 0.30341f
C30157 a_54780_2727# VGND 0.30341f
C30158 a_54332_2727# VGND 0.30712f
C30159 a_53660_2727# VGND 0.30848f
C30160 a_53212_2727# VGND 0.30341f
C30161 a_52764_2727# VGND 0.30581f
C30162 a_52316_2727# VGND 0.30765f
C30163 a_51868_2727# VGND 0.30974f
C30164 a_51420_2727# VGND 0.31256f
C30165 a_50972_2727# VGND 0.33819f
C30166 a_50524_2727# VGND 0.30958f
C30167 a_49852_2727# VGND 0.30848f
C30168 a_49404_2727# VGND 0.30341f
C30169 a_48956_2727# VGND 0.30341f
C30170 a_48508_2727# VGND 0.30341f
C30171 a_48060_2727# VGND 0.30341f
C30172 a_47612_2727# VGND 0.30341f
C30173 a_47164_2727# VGND 0.30341f
C30174 a_46716_2727# VGND 0.30712f
C30175 a_46044_2727# VGND 0.30848f
C30176 a_45596_2727# VGND 0.30341f
C30177 a_45148_2727# VGND 0.30419f
C30178 a_44700_2727# VGND 0.30708f
C30179 a_44252_2727# VGND 0.30894f
C30180 a_43804_2727# VGND 0.31126f
C30181 a_43356_2727# VGND 0.34666f
C30182 a_42908_2727# VGND 0.31456f
C30183 a_42236_2727# VGND 0.30848f
C30184 a_41788_2727# VGND 0.30341f
C30185 a_41340_2727# VGND 0.30341f
C30186 a_40892_2727# VGND 0.30341f
C30187 a_40444_2727# VGND 0.30341f
C30188 a_39996_2727# VGND 0.30341f
C30189 a_39548_2727# VGND 0.30341f
C30190 a_39100_2727# VGND 0.30712f
C30191 a_38428_2727# VGND 0.30848f
C30192 a_37980_2727# VGND 0.30341f
C30193 a_37532_2727# VGND 0.30341f
C30194 a_37084_2727# VGND 0.30659f
C30195 a_36636_2727# VGND 0.3082f
C30196 a_36188_2727# VGND 0.31043f
C30197 a_35740_2727# VGND 0.32632f
C30198 a_35292_2727# VGND 0.32264f
C30199 a_34620_2727# VGND 0.30848f
C30200 a_34172_2727# VGND 0.30341f
C30201 a_33724_2727# VGND 0.30341f
C30202 a_33276_2727# VGND 0.30341f
C30203 a_32828_2727# VGND 0.30341f
C30204 a_32380_2727# VGND 0.30341f
C30205 a_31932_2727# VGND 0.30341f
C30206 a_31484_2727# VGND 0.30712f
C30207 a_30812_2727# VGND 0.30848f
C30208 a_30364_2727# VGND 0.30341f
C30209 a_29916_2727# VGND 0.30341f
C30210 a_29468_2727# VGND 0.30558f
C30211 a_29020_2727# VGND 0.30755f
C30212 a_28572_2727# VGND 0.30961f
C30213 a_28124_2727# VGND 0.31231f
C30214 a_27676_2727# VGND 0.34503f
C30215 a_27004_2727# VGND 0.30863f
C30216 a_26556_2727# VGND 0.30341f
C30217 a_26108_2727# VGND 0.30341f
C30218 a_25660_2727# VGND 0.30341f
C30219 a_25212_2727# VGND 0.30341f
C30220 a_24764_2727# VGND 0.30341f
C30221 a_24316_2727# VGND 0.30341f
C30222 a_23868_2727# VGND 0.30712f
C30223 a_23196_2727# VGND 0.30848f
C30224 a_22748_2727# VGND 0.30341f
C30225 a_22300_2727# VGND 0.30341f
C30226 a_21852_2727# VGND 0.30392f
C30227 a_21404_2727# VGND 0.30699f
C30228 a_20956_2727# VGND 0.30881f
C30229 a_20508_2727# VGND 0.31112f
C30230 a_20060_2727# VGND 0.34605f
C30231 a_19388_2727# VGND 0.30977f
C30232 a_18940_2727# VGND 0.30341f
C30233 a_18492_2727# VGND 0.30341f
C30234 a_18044_2727# VGND 0.30341f
C30235 a_17596_2727# VGND 0.30341f
C30236 a_17148_2727# VGND 0.30341f
C30237 a_16700_2727# VGND 0.30341f
C30238 a_16252_2727# VGND 0.30712f
C30239 a_15580_2727# VGND 0.30848f
C30240 a_15132_2727# VGND 0.30341f
C30241 a_14684_2727# VGND 0.30341f
C30242 a_14236_2727# VGND 0.30341f
C30243 a_13788_2727# VGND 0.30652f
C30244 a_13340_2727# VGND 0.30809f
C30245 a_12892_2727# VGND 0.3103f
C30246 a_12444_2727# VGND 0.32694f
C30247 a_11772_2727# VGND 0.3156f
C30248 a_11324_2727# VGND 0.30341f
C30249 a_10876_2727# VGND 0.30341f
C30250 a_10428_2727# VGND 0.30341f
C30251 a_9980_2727# VGND 0.30341f
C30252 a_9532_2727# VGND 0.30341f
C30253 a_9084_2727# VGND 0.30341f
C30254 a_8636_2727# VGND 0.30712f
C30255 a_7964_2727# VGND 0.30848f
C30256 a_7516_2727# VGND 0.30341f
C30257 a_7068_2727# VGND 0.30341f
C30258 a_6620_2727# VGND 0.30341f
C30259 a_6172_2727# VGND 0.30533f
C30260 a_5724_2727# VGND 0.29169f
C30261 a_5276_2727# VGND 0.29209f
C30262 a_4828_2727# VGND 0.29921f
C30263 a_4156_2727# VGND 0.2987f
C30264 a_3708_2727# VGND 0.2812f
C30265 a_3260_2727# VGND 0.2812f
C30266 a_2812_2727# VGND 0.2812f
C30267 a_2364_2727# VGND 0.2812f
C30268 a_1916_2727# VGND 0.2812f
C30269 a_1468_2727# VGND 0.2812f
C30270 a_1020_2727# VGND 0.29134f
C30271 a_67996_3160# VGND 0.29009f
C30272 a_67548_3160# VGND 0.29121f
C30273 a_67100_3160# VGND 0.28927f
C30274 a_66652_3160# VGND 0.3275f
C30275 a_66204_3160# VGND 0.28778f
C30276 a_65756_3160# VGND 0.2812f
C30277 a_65308_3160# VGND 0.28739f
C30278 a_64860_3160# VGND 0.28746f
C30279 a_64412_3160# VGND 0.29654f
C30280 a_67908_3204# VGND 0.4924f
C30281 a_67460_3204# VGND 0.444f
C30282 a_67012_3204# VGND 0.44727f
C30283 a_66564_3204# VGND 0.47245f
C30284 a_66116_3204# VGND 0.44079f
C30285 a_65668_3204# VGND 0.43828f
C30286 a_65220_3204# VGND 0.43828f
C30287 a_64772_3204# VGND 0.43828f
C30288 a_64324_3204# VGND 0.4664f
C30289 a_5052_3160# VGND 0.28763f
C30290 a_4604_3160# VGND 0.31741f
C30291 a_4156_3160# VGND 0.29553f
C30292 a_3708_3160# VGND 0.2812f
C30293 a_3260_3160# VGND 0.2812f
C30294 a_2812_3160# VGND 0.2812f
C30295 a_2364_3160# VGND 0.2812f
C30296 a_1916_3160# VGND 0.2812f
C30297 a_1468_3160# VGND 0.2812f
C30298 a_1020_3160# VGND 0.29134f
C30299 a_4964_3204# VGND 0.47812f
C30300 a_4516_3204# VGND 0.5182f
C30301 a_4068_3204# VGND 0.44538f
C30302 a_3620_3204# VGND 0.43828f
C30303 a_3172_3204# VGND 0.43828f
C30304 a_2724_3204# VGND 0.43828f
C30305 a_2276_3204# VGND 0.43828f
C30306 a_1828_3204# VGND 0.43828f
C30307 a_1380_3204# VGND 0.43828f
C30308 a_932_3204# VGND 0.4664f
C30309 a_67460_4392# VGND 0.45147f
C30310 a_67012_4392# VGND 0.44727f
C30311 a_66564_4392# VGND 0.47245f
C30312 a_66116_4392# VGND 0.44079f
C30313 a_65668_4392# VGND 0.43828f
C30314 a_65220_4392# VGND 0.43828f
C30315 a_64772_4392# VGND 0.43828f
C30316 a_64324_4392# VGND 0.4664f
C30317 a_5300_4392# VGND 0.4913f
C30318 a_4852_4392# VGND 0.48985f
C30319 a_4068_4392# VGND 0.44997f
C30320 a_3620_4392# VGND 0.43828f
C30321 a_3172_4392# VGND 0.43828f
C30322 a_2724_4392# VGND 0.43828f
C30323 a_2276_4392# VGND 0.43828f
C30324 a_1828_4392# VGND 0.43828f
C30325 a_1380_4392# VGND 0.43828f
C30326 a_932_4392# VGND 0.4664f
C30327 a_67548_4295# VGND 0.28805f
C30328 a_67100_4295# VGND 0.28927f
C30329 a_66652_4295# VGND 0.3275f
C30330 a_66204_4295# VGND 0.28778f
C30331 a_65756_4295# VGND 0.2812f
C30332 a_65308_4295# VGND 0.2812f
C30333 a_64860_4295# VGND 0.2812f
C30334 a_64412_4295# VGND 0.29134f
C30335 a_5388_4295# VGND 0.3139f
C30336 a_4940_4295# VGND 0.29949f
C30337 a_4156_4295# VGND 0.28278f
C30338 a_3708_4295# VGND 0.2812f
C30339 a_3260_4295# VGND 0.2812f
C30340 a_2812_4295# VGND 0.2812f
C30341 a_2364_4295# VGND 0.2812f
C30342 a_1916_4295# VGND 0.2812f
C30343 a_1468_4295# VGND 0.2812f
C30344 a_1020_4295# VGND 0.29134f
C30345 a_67996_4728# VGND 0.29348f
C30346 a_67548_4728# VGND 0.29121f
C30347 a_67100_4728# VGND 0.28927f
C30348 a_66652_4728# VGND 0.3275f
C30349 a_66204_4728# VGND 0.28778f
C30350 a_65756_4728# VGND 0.2812f
C30351 a_65308_4728# VGND 0.2812f
C30352 a_64860_4728# VGND 0.2812f
C30353 a_64412_4728# VGND 0.29134f
C30354 a_67908_4772# VGND 0.4924f
C30355 a_67460_4772# VGND 0.444f
C30356 a_67012_4772# VGND 0.44727f
C30357 a_66564_4772# VGND 0.47245f
C30358 a_66116_4772# VGND 0.44079f
C30359 a_65668_4772# VGND 0.43828f
C30360 a_65220_4772# VGND 0.43828f
C30361 a_64772_4772# VGND 0.43828f
C30362 a_64324_4772# VGND 0.4664f
C30363 a_5052_4728# VGND 0.28654f
C30364 a_4604_4728# VGND 0.31699f
C30365 a_4156_4728# VGND 0.29553f
C30366 a_3708_4728# VGND 0.2812f
C30367 a_3260_4728# VGND 0.2812f
C30368 a_2812_4728# VGND 0.2812f
C30369 a_2364_4728# VGND 0.2812f
C30370 a_1916_4728# VGND 0.2812f
C30371 a_1468_4728# VGND 0.2812f
C30372 a_1020_4728# VGND 0.29134f
C30373 a_4964_4772# VGND 0.47812f
C30374 a_4516_4772# VGND 0.5182f
C30375 a_4068_4772# VGND 0.44538f
C30376 a_3620_4772# VGND 0.43828f
C30377 a_3172_4772# VGND 0.43828f
C30378 a_2724_4772# VGND 0.43828f
C30379 a_2276_4772# VGND 0.43828f
C30380 a_1828_4772# VGND 0.43828f
C30381 a_1380_4772# VGND 0.43828f
C30382 a_932_4772# VGND 0.4664f
C30383 a_67460_5960# VGND 0.45147f
C30384 a_67012_5960# VGND 0.44727f
C30385 a_66564_5960# VGND 0.47245f
C30386 a_66116_5960# VGND 0.44079f
C30387 a_65668_5960# VGND 0.43828f
C30388 a_65220_5960# VGND 0.43828f
C30389 a_64772_5960# VGND 0.43828f
C30390 a_64324_5960# VGND 0.4664f
C30391 a_5300_5960# VGND 0.48995f
C30392 a_4852_5960# VGND 0.48956f
C30393 a_4068_5960# VGND 0.44997f
C30394 a_3620_5960# VGND 0.43828f
C30395 a_3172_5960# VGND 0.43828f
C30396 a_2724_5960# VGND 0.43828f
C30397 a_2276_5960# VGND 0.43828f
C30398 a_1828_5960# VGND 0.43828f
C30399 a_1380_5960# VGND 0.43828f
C30400 a_932_5960# VGND 0.4664f
C30401 a_67548_5863# VGND 0.28805f
C30402 a_67100_5863# VGND 0.28927f
C30403 a_66652_5863# VGND 0.3275f
C30404 a_66204_5863# VGND 0.28778f
C30405 a_65756_5863# VGND 0.2812f
C30406 a_65308_5863# VGND 0.2812f
C30407 a_64860_5863# VGND 0.2812f
C30408 a_64412_5863# VGND 0.29134f
C30409 a_5388_5863# VGND 0.3139f
C30410 a_4940_5863# VGND 0.29949f
C30411 a_4156_5863# VGND 0.28278f
C30412 a_3708_5863# VGND 0.2812f
C30413 a_3260_5863# VGND 0.2812f
C30414 a_2812_5863# VGND 0.2812f
C30415 a_2364_5863# VGND 0.2812f
C30416 a_1916_5863# VGND 0.2812f
C30417 a_1468_5863# VGND 0.2812f
C30418 a_1020_5863# VGND 0.29134f
C30419 a_67996_6296# VGND 0.29348f
C30420 a_67548_6296# VGND 0.29121f
C30421 a_67100_6296# VGND 0.28927f
C30422 a_66652_6296# VGND 0.3275f
C30423 a_66204_6296# VGND 0.28778f
C30424 a_65756_6296# VGND 0.2812f
C30425 a_65308_6296# VGND 0.2812f
C30426 a_64860_6296# VGND 0.2812f
C30427 a_64412_6296# VGND 0.29134f
C30428 a_67908_6340# VGND 0.4924f
C30429 a_67460_6340# VGND 0.444f
C30430 a_67012_6340# VGND 0.44727f
C30431 a_66564_6340# VGND 0.47245f
C30432 a_66116_6340# VGND 0.44079f
C30433 a_65668_6340# VGND 0.43828f
C30434 a_65220_6340# VGND 0.43828f
C30435 a_64772_6340# VGND 0.43828f
C30436 a_64324_6340# VGND 0.4664f
C30437 a_5052_6296# VGND 0.28654f
C30438 a_4604_6296# VGND 0.31699f
C30439 a_4156_6296# VGND 0.29553f
C30440 a_3708_6296# VGND 0.2812f
C30441 a_3260_6296# VGND 0.2812f
C30442 a_2812_6296# VGND 0.2812f
C30443 a_2364_6296# VGND 0.2812f
C30444 a_1916_6296# VGND 0.2812f
C30445 a_1468_6296# VGND 0.2812f
C30446 a_1020_6296# VGND 0.29134f
C30447 a_4964_6340# VGND 0.47812f
C30448 a_4516_6340# VGND 0.5182f
C30449 a_4068_6340# VGND 0.44538f
C30450 a_3620_6340# VGND 0.43828f
C30451 a_3172_6340# VGND 0.43828f
C30452 a_2724_6340# VGND 0.43828f
C30453 a_2276_6340# VGND 0.43828f
C30454 a_1828_6340# VGND 0.43828f
C30455 a_1380_6340# VGND 0.43828f
C30456 a_932_6340# VGND 0.4664f
C30457 a_67460_7528# VGND 0.45147f
C30458 a_67012_7528# VGND 0.44727f
C30459 a_66564_7528# VGND 0.47245f
C30460 a_66116_7528# VGND 0.44079f
C30461 a_65668_7528# VGND 0.43828f
C30462 a_65220_7528# VGND 0.43828f
C30463 a_64772_7528# VGND 0.43828f
C30464 a_64324_7528# VGND 0.4664f
C30465 a_5300_7528# VGND 0.48995f
C30466 a_4852_7528# VGND 0.48956f
C30467 a_4068_7528# VGND 0.44997f
C30468 a_3620_7528# VGND 0.43828f
C30469 a_3172_7528# VGND 0.43828f
C30470 a_2724_7528# VGND 0.43828f
C30471 a_2276_7528# VGND 0.43828f
C30472 a_1828_7528# VGND 0.43828f
C30473 a_1380_7528# VGND 0.43828f
C30474 a_932_7528# VGND 0.4664f
C30475 a_67548_7431# VGND 0.28805f
C30476 a_67100_7431# VGND 0.28927f
C30477 a_66652_7431# VGND 0.3275f
C30478 a_66204_7431# VGND 0.28778f
C30479 a_65756_7431# VGND 0.2812f
C30480 a_65308_7431# VGND 0.2812f
C30481 a_64860_7431# VGND 0.2812f
C30482 a_64412_7431# VGND 0.29134f
C30483 a_5388_7431# VGND 0.3139f
C30484 a_4940_7431# VGND 0.29949f
C30485 a_4156_7431# VGND 0.28278f
C30486 a_3708_7431# VGND 0.2812f
C30487 a_3260_7431# VGND 0.2812f
C30488 a_2812_7431# VGND 0.2812f
C30489 a_2364_7431# VGND 0.2812f
C30490 a_1916_7431# VGND 0.2812f
C30491 a_1468_7431# VGND 0.2812f
C30492 a_1020_7431# VGND 0.29134f
C30493 a_67996_7864# VGND 0.29348f
C30494 a_67548_7864# VGND 0.29121f
C30495 a_67100_7864# VGND 0.28927f
C30496 a_66652_7864# VGND 0.3275f
C30497 a_66204_7864# VGND 0.28778f
C30498 a_65756_7864# VGND 0.2812f
C30499 a_65308_7864# VGND 0.2812f
C30500 a_64860_7864# VGND 0.2812f
C30501 a_64412_7864# VGND 0.29134f
C30502 a_67908_7908# VGND 0.49483f
C30503 a_67460_7908# VGND 0.444f
C30504 a_67012_7908# VGND 0.44727f
C30505 a_66564_7908# VGND 0.47245f
C30506 a_66116_7908# VGND 0.44079f
C30507 a_65668_7908# VGND 0.43828f
C30508 a_65220_7908# VGND 0.43828f
C30509 a_64772_7908# VGND 0.43828f
C30510 a_64324_7908# VGND 0.4664f
C30511 a_5052_7864# VGND 0.28654f
C30512 a_4604_7864# VGND 0.31699f
C30513 a_4156_7864# VGND 0.29553f
C30514 a_3708_7864# VGND 0.2812f
C30515 a_3260_7864# VGND 0.2812f
C30516 a_2812_7864# VGND 0.2812f
C30517 a_2364_7864# VGND 0.2812f
C30518 a_1916_7864# VGND 0.2812f
C30519 a_1468_7864# VGND 0.2812f
C30520 a_1020_7864# VGND 0.29134f
C30521 a_4964_7908# VGND 0.47812f
C30522 a_4516_7908# VGND 0.5182f
C30523 a_4068_7908# VGND 0.44538f
C30524 a_3620_7908# VGND 0.43828f
C30525 a_3172_7908# VGND 0.43828f
C30526 a_2724_7908# VGND 0.43828f
C30527 a_2276_7908# VGND 0.43828f
C30528 a_1828_7908# VGND 0.43828f
C30529 a_1380_7908# VGND 0.43828f
C30530 a_932_7908# VGND 0.4664f
C30531 a_67460_9096# VGND 0.45147f
C30532 a_67012_9096# VGND 0.44727f
C30533 a_66564_9096# VGND 0.47245f
C30534 a_66116_9096# VGND 0.44079f
C30535 a_65668_9096# VGND 0.43828f
C30536 a_65220_9096# VGND 0.43828f
C30537 a_64772_9096# VGND 0.43828f
C30538 a_64324_9096# VGND 0.4664f
C30539 a_5300_9096# VGND 0.48995f
C30540 a_4852_9096# VGND 0.48956f
C30541 a_4068_9096# VGND 0.44997f
C30542 a_3620_9096# VGND 0.43828f
C30543 a_3172_9096# VGND 0.43828f
C30544 a_2724_9096# VGND 0.43828f
C30545 a_2276_9096# VGND 0.43828f
C30546 a_1828_9096# VGND 0.43828f
C30547 a_1380_9096# VGND 0.43828f
C30548 a_932_9096# VGND 0.4664f
C30549 a_67548_8999# VGND 0.28805f
C30550 a_67100_8999# VGND 0.28927f
C30551 a_66652_8999# VGND 0.3275f
C30552 a_66204_8999# VGND 0.28778f
C30553 a_65756_8999# VGND 0.2812f
C30554 a_65308_8999# VGND 0.2812f
C30555 a_64860_8999# VGND 0.2812f
C30556 a_64412_8999# VGND 0.29028f
C30557 a_5388_8999# VGND 0.3139f
C30558 a_4940_8999# VGND 0.29949f
C30559 a_4156_8999# VGND 0.28278f
C30560 a_3708_8999# VGND 0.2812f
C30561 a_3260_8999# VGND 0.2812f
C30562 a_2812_8999# VGND 0.2812f
C30563 a_2364_8999# VGND 0.2812f
C30564 a_1916_8999# VGND 0.2812f
C30565 a_1468_8999# VGND 0.2812f
C30566 a_1020_8999# VGND 0.29134f
C30567 a_67548_9432# VGND 0.30676f
C30568 a_67100_9432# VGND 0.28927f
C30569 a_66652_9432# VGND 0.3275f
C30570 a_66204_9432# VGND 0.28778f
C30571 a_65756_9432# VGND 0.2812f
C30572 a_65308_9432# VGND 0.2812f
C30573 a_64860_9432# VGND 0.2812f
C30574 a_64412_9432# VGND 0.28492f
C30575 a_67460_9476# VGND 0.4713f
C30576 a_67012_9476# VGND 0.46622f
C30577 a_66564_9476# VGND 0.49291f
C30578 a_66116_9476# VGND 0.45973f
C30579 a_65668_9476# VGND 0.45723f
C30580 a_65220_9476# VGND 0.45723f
C30581 a_64772_9476# VGND 0.45723f
C30582 a_64324_9476# VGND 0.46809f
C30583 a_63740_9432# VGND 0.30848f
C30584 a_63292_9432# VGND 0.30341f
C30585 a_62844_9432# VGND 0.30341f
C30586 a_62396_9432# VGND 0.30341f
C30587 a_61948_9432# VGND 0.30341f
C30588 a_61500_9432# VGND 0.30341f
C30589 a_61052_9432# VGND 0.30341f
C30590 a_60604_9432# VGND 0.30888f
C30591 a_63652_9476# VGND 0.45972f
C30592 a_63204_9476# VGND 0.45589f
C30593 a_62756_9476# VGND 0.45589f
C30594 a_62308_9476# VGND 0.45589f
C30595 a_61860_9476# VGND 0.45589f
C30596 a_61412_9476# VGND 0.45589f
C30597 a_60964_9476# VGND 0.45589f
C30598 a_60516_9476# VGND 0.47168f
C30599 a_59932_9432# VGND 0.31339f
C30600 a_59484_9432# VGND 0.31056f
C30601 a_59036_9432# VGND 0.32954f
C30602 a_58588_9432# VGND 0.31523f
C30603 a_58140_9432# VGND 0.30341f
C30604 a_57692_9432# VGND 0.30341f
C30605 a_57244_9432# VGND 0.30341f
C30606 a_56796_9432# VGND 0.30712f
C30607 a_59844_9476# VGND 0.46342f
C30608 a_59396_9476# VGND 0.46226f
C30609 a_58948_9476# VGND 0.48975f
C30610 a_58500_9476# VGND 0.46249f
C30611 a_58052_9476# VGND 0.45465f
C30612 a_57604_9476# VGND 0.45465f
C30613 a_57156_9476# VGND 0.45465f
C30614 a_56708_9476# VGND 0.4816f
C30615 a_56124_9432# VGND 0.30848f
C30616 a_55676_9432# VGND 0.30341f
C30617 a_55228_9432# VGND 0.30341f
C30618 a_54780_9432# VGND 0.30341f
C30619 a_54332_9432# VGND 0.30341f
C30620 a_53884_9432# VGND 0.30341f
C30621 a_53436_9432# VGND 0.30341f
C30622 a_52988_9432# VGND 0.30724f
C30623 a_56036_9476# VGND 0.45987f
C30624 a_55588_9476# VGND 0.45604f
C30625 a_55140_9476# VGND 0.45604f
C30626 a_54692_9476# VGND 0.45604f
C30627 a_54244_9476# VGND 0.45604f
C30628 a_53796_9476# VGND 0.45604f
C30629 a_53348_9476# VGND 0.45604f
C30630 a_52900_9476# VGND 0.46909f
C30631 a_52316_9432# VGND 0.31273f
C30632 a_51868_9432# VGND 0.30974f
C30633 a_51420_9432# VGND 0.31256f
C30634 a_50972_9432# VGND 0.33819f
C30635 a_50524_9432# VGND 0.30587f
C30636 a_50076_9432# VGND 0.30341f
C30637 a_49628_9432# VGND 0.30341f
C30638 a_49180_9432# VGND 0.30712f
C30639 a_52228_9476# VGND 0.46531f
C30640 a_51780_9476# VGND 0.46367f
C30641 a_51332_9476# VGND 0.47499f
C30642 a_50884_9476# VGND 0.47478f
C30643 a_50436_9476# VGND 0.45724f
C30644 a_49988_9476# VGND 0.45724f
C30645 a_49540_9476# VGND 0.45724f
C30646 a_49092_9476# VGND 0.4693f
C30647 a_48508_9432# VGND 0.30848f
C30648 a_48060_9432# VGND 0.30341f
C30649 a_47612_9432# VGND 0.30341f
C30650 a_47164_9432# VGND 0.30341f
C30651 a_46716_9432# VGND 0.30341f
C30652 a_46268_9432# VGND 0.30341f
C30653 a_45820_9432# VGND 0.30341f
C30654 a_45372_9432# VGND 0.31355f
C30655 a_48420_9476# VGND 0.44211f
C30656 a_47972_9476# VGND 0.43828f
C30657 a_47524_9476# VGND 0.43828f
C30658 a_47076_9476# VGND 0.43828f
C30659 a_46628_9476# VGND 0.43828f
C30660 a_46180_9476# VGND 0.43828f
C30661 a_45732_9476# VGND 0.43828f
C30662 a_45284_9476# VGND 0.4664f
C30663 a_5052_9432# VGND 0.28654f
C30664 a_4604_9432# VGND 0.31699f
C30665 a_4156_9432# VGND 0.29553f
C30666 a_3708_9432# VGND 0.2812f
C30667 a_3260_9432# VGND 0.2812f
C30668 a_2812_9432# VGND 0.2812f
C30669 a_2364_9432# VGND 0.2812f
C30670 a_1916_9432# VGND 0.2812f
C30671 a_1468_9432# VGND 0.2812f
C30672 a_1020_9432# VGND 0.29134f
C30673 a_4964_9476# VGND 0.47812f
C30674 a_4516_9476# VGND 0.5182f
C30675 a_4068_9476# VGND 0.44538f
C30676 a_3620_9476# VGND 0.43828f
C30677 a_3172_9476# VGND 0.43828f
C30678 a_2724_9476# VGND 0.43828f
C30679 a_2276_9476# VGND 0.43828f
C30680 a_1828_9476# VGND 0.43828f
C30681 a_1380_9476# VGND 0.43828f
C30682 a_932_9476# VGND 0.4664f
C30683 a_68020_10664# VGND 0.48098f
C30684 a_67572_10664# VGND 0.46116f
C30685 a_67124_10664# VGND 0.46394f
C30686 a_66676_10664# VGND 0.49854f
C30687 a_66228_10664# VGND 0.46139f
C30688 a_65780_10664# VGND 0.456f
C30689 a_65332_10664# VGND 0.456f
C30690 a_64884_10664# VGND 0.46806f
C30691 a_64212_10664# VGND 0.47318f
C30692 a_63764_10664# VGND 0.45815f
C30693 a_63316_10664# VGND 0.45848f
C30694 a_62868_10664# VGND 0.45848f
C30695 a_62420_10664# VGND 0.45848f
C30696 a_61972_10664# VGND 0.45848f
C30697 a_61524_10664# VGND 0.45848f
C30698 a_61076_10664# VGND 0.45848f
C30699 a_60628_10664# VGND 0.45986f
C30700 a_60180_10664# VGND 0.47837f
C30701 a_59732_10664# VGND 0.4652f
C30702 a_59284_10664# VGND 0.46815f
C30703 a_58836_10664# VGND 0.50255f
C30704 a_58388_10664# VGND 0.46328f
C30705 a_57940_10664# VGND 0.45971f
C30706 a_57492_10664# VGND 0.45971f
C30707 a_57044_10664# VGND 0.47167f
C30708 a_56372_10664# VGND 0.48871f
C30709 a_55924_10664# VGND 0.45971f
C30710 a_55476_10664# VGND 0.45971f
C30711 a_55028_10664# VGND 0.45971f
C30712 a_54580_10664# VGND 0.45971f
C30713 a_54132_10664# VGND 0.45971f
C30714 a_53684_10664# VGND 0.45971f
C30715 a_53236_10664# VGND 0.45971f
C30716 a_52788_10664# VGND 0.46167f
C30717 a_52340_10664# VGND 0.46228f
C30718 a_51892_10664# VGND 0.4643f
C30719 a_51444_10664# VGND 0.46779f
C30720 a_50996_10664# VGND 0.4917f
C30721 a_50548_10664# VGND 0.46052f
C30722 a_50100_10664# VGND 0.45848f
C30723 a_49652_10664# VGND 0.45848f
C30724 a_49204_10664# VGND 0.47298f
C30725 a_48420_10664# VGND 0.44215f
C30726 a_47972_10664# VGND 0.43828f
C30727 a_47524_10664# VGND 0.43828f
C30728 a_47076_10664# VGND 0.43828f
C30729 a_46628_10664# VGND 0.43828f
C30730 a_46180_10664# VGND 0.43828f
C30731 a_45732_10664# VGND 0.43828f
C30732 a_45284_10664# VGND 0.4664f
C30733 a_5300_10664# VGND 0.48995f
C30734 a_4852_10664# VGND 0.48956f
C30735 a_4068_10664# VGND 0.44997f
C30736 a_3620_10664# VGND 0.43828f
C30737 a_3172_10664# VGND 0.43828f
C30738 a_2724_10664# VGND 0.43828f
C30739 a_2276_10664# VGND 0.43828f
C30740 a_1828_10664# VGND 0.43828f
C30741 a_1380_10664# VGND 0.43828f
C30742 a_932_10664# VGND 0.4664f
C30743 a_68108_10567# VGND 0.31063f
C30744 a_67660_10567# VGND 0.28822f
C30745 a_67212_10567# VGND 0.29048f
C30746 a_66764_10567# VGND 0.31433f
C30747 a_66316_10567# VGND 0.29333f
C30748 a_65868_10567# VGND 0.2831f
C30749 a_65420_10567# VGND 0.2831f
C30750 a_64972_10567# VGND 0.28681f
C30751 a_64300_10567# VGND 0.28946f
C30752 a_63852_10567# VGND 0.28758f
C30753 a_63404_10567# VGND 0.2841f
C30754 a_62956_10567# VGND 0.2841f
C30755 a_62508_10567# VGND 0.2841f
C30756 a_62060_10567# VGND 0.2841f
C30757 a_61612_10567# VGND 0.2841f
C30758 a_61164_10567# VGND 0.2841f
C30759 a_60716_10567# VGND 0.28633f
C30760 a_60268_10567# VGND 0.28787f
C30761 a_59820_10567# VGND 0.28969f
C30762 a_59372_10567# VGND 0.29201f
C30763 a_58924_10567# VGND 0.32367f
C30764 a_58476_10567# VGND 0.29233f
C30765 a_58028_10567# VGND 0.28426f
C30766 a_57580_10567# VGND 0.28426f
C30767 a_57132_10567# VGND 0.28776f
C30768 a_56460_10567# VGND 0.28946f
C30769 a_56012_10567# VGND 0.28758f
C30770 a_55564_10567# VGND 0.2841f
C30771 a_55116_10567# VGND 0.2841f
C30772 a_54668_10567# VGND 0.2841f
C30773 a_54220_10567# VGND 0.2841f
C30774 a_53772_10567# VGND 0.2841f
C30775 a_53324_10567# VGND 0.2841f
C30776 a_52876_10567# VGND 0.28701f
C30777 a_52428_10567# VGND 0.2881f
C30778 a_51980_10567# VGND 0.29002f
C30779 a_51532_10567# VGND 0.2925f
C30780 a_51084_10567# VGND 0.3315f
C30781 a_50636_10567# VGND 0.29011f
C30782 a_50188_10567# VGND 0.28426f
C30783 a_49740_10567# VGND 0.28426f
C30784 a_49292_10567# VGND 0.28799f
C30785 a_48508_10567# VGND 0.26958f
C30786 a_48060_10567# VGND 0.2812f
C30787 a_47612_10567# VGND 0.2812f
C30788 a_47164_10567# VGND 0.2812f
C30789 a_46716_10567# VGND 0.2812f
C30790 a_46268_10567# VGND 0.2812f
C30791 a_45820_10567# VGND 0.2812f
C30792 a_45372_10567# VGND 0.29134f
C30793 a_5388_10567# VGND 0.3139f
C30794 a_4940_10567# VGND 0.29949f
C30795 a_4156_10567# VGND 0.28278f
C30796 a_3708_10567# VGND 0.2812f
C30797 a_3260_10567# VGND 0.2812f
C30798 a_2812_10567# VGND 0.2812f
C30799 a_2364_10567# VGND 0.2812f
C30800 a_1916_10567# VGND 0.2812f
C30801 a_1468_10567# VGND 0.2812f
C30802 a_1020_10567# VGND 0.29134f
C30803 a_67772_11000# VGND 0.28474f
C30804 a_67324_11000# VGND 0.29263f
C30805 a_66876_11000# VGND 0.30298f
C30806 a_66428_11000# VGND 0.30915f
C30807 a_65980_11000# VGND 0.28588f
C30808 a_65532_11000# VGND 0.28581f
C30809 a_65084_11000# VGND 0.28581f
C30810 a_64636_11000# VGND 0.28875f
C30811 a_64188_11000# VGND 0.28594f
C30812 a_63740_11000# VGND 0.28426f
C30813 a_63292_11000# VGND 0.28426f
C30814 a_62844_11000# VGND 0.28426f
C30815 a_62396_11000# VGND 0.28426f
C30816 a_61948_11000# VGND 0.28426f
C30817 a_61500_11000# VGND 0.28426f
C30818 a_61052_11000# VGND 0.28776f
C30819 a_67684_11044# VGND 0.46786f
C30820 a_67236_11044# VGND 0.46378f
C30821 a_66788_11044# VGND 0.48615f
C30822 a_66340_11044# VGND 0.46546f
C30823 a_65892_11044# VGND 0.45666f
C30824 a_65444_11044# VGND 0.45666f
C30825 a_64996_11044# VGND 0.45666f
C30826 a_64548_11044# VGND 0.47155f
C30827 a_64100_11044# VGND 0.45794f
C30828 a_63652_11044# VGND 0.4579f
C30829 a_63204_11044# VGND 0.4579f
C30830 a_62756_11044# VGND 0.4579f
C30831 a_62308_11044# VGND 0.4579f
C30832 a_61860_11044# VGND 0.4579f
C30833 a_61412_11044# VGND 0.4579f
C30834 a_60964_11044# VGND 0.46986f
C30835 a_60380_11000# VGND 0.29443f
C30836 a_59932_11000# VGND 0.29249f
C30837 a_59484_11000# VGND 0.29125f
C30838 a_59036_11000# VGND 0.30936f
C30839 a_58588_11000# VGND 0.29592f
C30840 a_58140_11000# VGND 0.2841f
C30841 a_57692_11000# VGND 0.2841f
C30842 a_57244_11000# VGND 0.2841f
C30843 a_56796_11000# VGND 0.28575f
C30844 a_56348_11000# VGND 0.2859f
C30845 a_55900_11000# VGND 0.28589f
C30846 a_55452_11000# VGND 0.28589f
C30847 a_55004_11000# VGND 0.28589f
C30848 a_54556_11000# VGND 0.28589f
C30849 a_54108_11000# VGND 0.28589f
C30850 a_53660_11000# VGND 0.28589f
C30851 a_53212_11000# VGND 0.28939f
C30852 a_60292_11044# VGND 0.47377f
C30853 a_59844_11044# VGND 0.4616f
C30854 a_59396_11044# VGND 0.46427f
C30855 a_58948_11044# VGND 0.49373f
C30856 a_58500_11044# VGND 0.4645f
C30857 a_58052_11044# VGND 0.45666f
C30858 a_57604_11044# VGND 0.45666f
C30859 a_57156_11044# VGND 0.45666f
C30860 a_56708_11044# VGND 0.47155f
C30861 a_56260_11044# VGND 0.45794f
C30862 a_55812_11044# VGND 0.4579f
C30863 a_55364_11044# VGND 0.4579f
C30864 a_54916_11044# VGND 0.4579f
C30865 a_54468_11044# VGND 0.4579f
C30866 a_54020_11044# VGND 0.4579f
C30867 a_53572_11044# VGND 0.4579f
C30868 a_53124_11044# VGND 0.46986f
C30869 a_52540_11000# VGND 0.2946f
C30870 a_52092_11000# VGND 0.29451f
C30871 a_51644_11000# VGND 0.2933f
C30872 a_51196_11000# VGND 0.32041f
C30873 a_50748_11000# VGND 0.29567f
C30874 a_50300_11000# VGND 0.28581f
C30875 a_49852_11000# VGND 0.28581f
C30876 a_49404_11000# VGND 0.28581f
C30877 a_48956_11000# VGND 0.28879f
C30878 a_48508_11000# VGND 0.28236f
C30879 a_48060_11000# VGND 0.28236f
C30880 a_47612_11000# VGND 0.28236f
C30881 a_47164_11000# VGND 0.28236f
C30882 a_46716_11000# VGND 0.28236f
C30883 a_46268_11000# VGND 0.28236f
C30884 a_45820_11000# VGND 0.28236f
C30885 a_45372_11000# VGND 0.29228f
C30886 a_52452_11044# VGND 0.47398f
C30887 a_52004_11044# VGND 0.46192f
C30888 a_51556_11044# VGND 0.46474f
C30889 a_51108_11044# VGND 0.50076f
C30890 a_50660_11044# VGND 0.46148f
C30891 a_50212_11044# VGND 0.45666f
C30892 a_49764_11044# VGND 0.45666f
C30893 a_49316_11044# VGND 0.45666f
C30894 a_48868_11044# VGND 0.47155f
C30895 a_48420_11044# VGND 0.44029f
C30896 a_47972_11044# VGND 0.44029f
C30897 a_47524_11044# VGND 0.44029f
C30898 a_47076_11044# VGND 0.44029f
C30899 a_46628_11044# VGND 0.44029f
C30900 a_46180_11044# VGND 0.44029f
C30901 a_45732_11044# VGND 0.44029f
C30902 a_45284_11044# VGND 0.46832f
C30903 a_5052_11000# VGND 0.28654f
C30904 a_4604_11000# VGND 0.31699f
C30905 a_4156_11000# VGND 0.29553f
C30906 a_3708_11000# VGND 0.2812f
C30907 a_3260_11000# VGND 0.2812f
C30908 a_2812_11000# VGND 0.2812f
C30909 a_2364_11000# VGND 0.2812f
C30910 a_1916_11000# VGND 0.2812f
C30911 a_1468_11000# VGND 0.2812f
C30912 a_1020_11000# VGND 0.29134f
C30913 a_4964_11044# VGND 0.47812f
C30914 a_4516_11044# VGND 0.5182f
C30915 a_4068_11044# VGND 0.44538f
C30916 a_3620_11044# VGND 0.43828f
C30917 a_3172_11044# VGND 0.43828f
C30918 a_2724_11044# VGND 0.43828f
C30919 a_2276_11044# VGND 0.43828f
C30920 a_1828_11044# VGND 0.43828f
C30921 a_1380_11044# VGND 0.43828f
C30922 a_932_11044# VGND 0.4664f
C30923 a_68020_12232# VGND 0.47855f
C30924 a_67572_12232# VGND 0.46105f
C30925 a_67124_12232# VGND 0.46383f
C30926 a_66676_12232# VGND 0.49822f
C30927 a_66228_12232# VGND 0.46128f
C30928 a_65780_12232# VGND 0.45589f
C30929 a_65332_12232# VGND 0.45589f
C30930 a_64884_12232# VGND 0.46795f
C30931 a_64212_12232# VGND 0.47057f
C30932 a_63764_12232# VGND 0.45666f
C30933 a_63316_12232# VGND 0.45666f
C30934 a_62868_12232# VGND 0.45666f
C30935 a_62420_12232# VGND 0.45666f
C30936 a_61972_12232# VGND 0.45666f
C30937 a_61524_12232# VGND 0.45666f
C30938 a_61076_12232# VGND 0.45666f
C30939 a_60628_12232# VGND 0.47293f
C30940 a_60180_12232# VGND 0.46151f
C30941 a_59732_12232# VGND 0.46339f
C30942 a_59284_12232# VGND 0.46634f
C30943 a_58836_12232# VGND 0.49982f
C30944 a_58388_12232# VGND 0.46146f
C30945 a_57940_12232# VGND 0.4579f
C30946 a_57492_12232# VGND 0.4579f
C30947 a_57044_12232# VGND 0.46986f
C30948 a_56372_12232# VGND 0.47057f
C30949 a_55924_12232# VGND 0.45666f
C30950 a_55476_12232# VGND 0.45666f
C30951 a_55028_12232# VGND 0.45666f
C30952 a_54580_12232# VGND 0.45666f
C30953 a_54132_12232# VGND 0.45666f
C30954 a_53684_12232# VGND 0.45666f
C30955 a_53236_12232# VGND 0.45666f
C30956 a_52788_12232# VGND 0.47351f
C30957 a_52340_12232# VGND 0.46174f
C30958 a_51892_12232# VGND 0.46372f
C30959 a_51444_12232# VGND 0.46721f
C30960 a_50996_12232# VGND 0.49018f
C30961 a_50548_12232# VGND 0.45994f
C30962 a_50100_12232# VGND 0.4579f
C30963 a_49652_12232# VGND 0.4579f
C30964 a_49204_12232# VGND 0.4724f
C30965 a_48420_12232# VGND 0.44215f
C30966 a_47972_12232# VGND 0.43828f
C30967 a_47524_12232# VGND 0.43828f
C30968 a_47076_12232# VGND 0.43828f
C30969 a_46628_12232# VGND 0.43828f
C30970 a_46180_12232# VGND 0.43828f
C30971 a_45732_12232# VGND 0.43828f
C30972 a_45284_12232# VGND 0.4664f
C30973 a_5300_12232# VGND 0.48995f
C30974 a_4852_12232# VGND 0.48956f
C30975 a_4068_12232# VGND 0.44997f
C30976 a_3620_12232# VGND 0.43828f
C30977 a_3172_12232# VGND 0.43828f
C30978 a_2724_12232# VGND 0.43828f
C30979 a_2276_12232# VGND 0.43828f
C30980 a_1828_12232# VGND 0.43828f
C30981 a_1380_12232# VGND 0.43828f
C30982 a_932_12232# VGND 0.4664f
C30983 a_68108_12135# VGND 0.31063f
C30984 a_67660_12135# VGND 0.28822f
C30985 a_67212_12135# VGND 0.29048f
C30986 a_66764_12135# VGND 0.31433f
C30987 a_66316_12135# VGND 0.29333f
C30988 a_65868_12135# VGND 0.2831f
C30989 a_65420_12135# VGND 0.2831f
C30990 a_64972_12135# VGND 0.28681f
C30991 a_64300_12135# VGND 0.28946f
C30992 a_63852_12135# VGND 0.28758f
C30993 a_63404_12135# VGND 0.2841f
C30994 a_62956_12135# VGND 0.2841f
C30995 a_62508_12135# VGND 0.2841f
C30996 a_62060_12135# VGND 0.2841f
C30997 a_61612_12135# VGND 0.2841f
C30998 a_61164_12135# VGND 0.2841f
C30999 a_60716_12135# VGND 0.28633f
C31000 a_60268_12135# VGND 0.28787f
C31001 a_59820_12135# VGND 0.28969f
C31002 a_59372_12135# VGND 0.29201f
C31003 a_58924_12135# VGND 0.32367f
C31004 a_58476_12135# VGND 0.29233f
C31005 a_58028_12135# VGND 0.28426f
C31006 a_57580_12135# VGND 0.28426f
C31007 a_57132_12135# VGND 0.28776f
C31008 a_56460_12135# VGND 0.28946f
C31009 a_56012_12135# VGND 0.28758f
C31010 a_55564_12135# VGND 0.2841f
C31011 a_55116_12135# VGND 0.2841f
C31012 a_54668_12135# VGND 0.2841f
C31013 a_54220_12135# VGND 0.2841f
C31014 a_53772_12135# VGND 0.2841f
C31015 a_53324_12135# VGND 0.2841f
C31016 a_52876_12135# VGND 0.28701f
C31017 a_52428_12135# VGND 0.2881f
C31018 a_51980_12135# VGND 0.29002f
C31019 a_51532_12135# VGND 0.2925f
C31020 a_51084_12135# VGND 0.3315f
C31021 a_50636_12135# VGND 0.29011f
C31022 a_50188_12135# VGND 0.28426f
C31023 a_49740_12135# VGND 0.28426f
C31024 a_49292_12135# VGND 0.28799f
C31025 a_48508_12135# VGND 0.26958f
C31026 a_48060_12135# VGND 0.2812f
C31027 a_47612_12135# VGND 0.2812f
C31028 a_47164_12135# VGND 0.2812f
C31029 a_46716_12135# VGND 0.2812f
C31030 a_46268_12135# VGND 0.2812f
C31031 a_45820_12135# VGND 0.2812f
C31032 a_45372_12135# VGND 0.29134f
C31033 a_5388_12135# VGND 0.3139f
C31034 a_4940_12135# VGND 0.29949f
C31035 a_4156_12135# VGND 0.28278f
C31036 a_3708_12135# VGND 0.2812f
C31037 a_3260_12135# VGND 0.2812f
C31038 a_2812_12135# VGND 0.2812f
C31039 a_2364_12135# VGND 0.2812f
C31040 a_1916_12135# VGND 0.2812f
C31041 a_1468_12135# VGND 0.2812f
C31042 a_1020_12135# VGND 0.29134f
C31043 a_67772_12568# VGND 0.28307f
C31044 a_67324_12568# VGND 0.29092f
C31045 a_66876_12568# VGND 0.30126f
C31046 a_66428_12568# VGND 0.30744f
C31047 a_65980_12568# VGND 0.28416f
C31048 a_65532_12568# VGND 0.2841f
C31049 a_65084_12568# VGND 0.2841f
C31050 a_64636_12568# VGND 0.28575f
C31051 a_64188_12568# VGND 0.28427f
C31052 a_63740_12568# VGND 0.28426f
C31053 a_63292_12568# VGND 0.28426f
C31054 a_62844_12568# VGND 0.28426f
C31055 a_62396_12568# VGND 0.28426f
C31056 a_61948_12568# VGND 0.28426f
C31057 a_61500_12568# VGND 0.28426f
C31058 a_61052_12568# VGND 0.28776f
C31059 a_67684_12612# VGND 0.46786f
C31060 a_67236_12612# VGND 0.46378f
C31061 a_66788_12612# VGND 0.48615f
C31062 a_66340_12612# VGND 0.46546f
C31063 a_65892_12612# VGND 0.45666f
C31064 a_65444_12612# VGND 0.45666f
C31065 a_64996_12612# VGND 0.45666f
C31066 a_64548_12612# VGND 0.47155f
C31067 a_64100_12612# VGND 0.45794f
C31068 a_63652_12612# VGND 0.4579f
C31069 a_63204_12612# VGND 0.4579f
C31070 a_62756_12612# VGND 0.4579f
C31071 a_62308_12612# VGND 0.4579f
C31072 a_61860_12612# VGND 0.4579f
C31073 a_61412_12612# VGND 0.4579f
C31074 a_60964_12612# VGND 0.46986f
C31075 a_60380_12568# VGND 0.29272f
C31076 a_59932_12568# VGND 0.29249f
C31077 a_59484_12568# VGND 0.29125f
C31078 a_59036_12568# VGND 0.30936f
C31079 a_58588_12568# VGND 0.29592f
C31080 a_58140_12568# VGND 0.2841f
C31081 a_57692_12568# VGND 0.2841f
C31082 a_57244_12568# VGND 0.2841f
C31083 a_56796_12568# VGND 0.28575f
C31084 a_56348_12568# VGND 0.28427f
C31085 a_55900_12568# VGND 0.28426f
C31086 a_55452_12568# VGND 0.28426f
C31087 a_55004_12568# VGND 0.28426f
C31088 a_54556_12568# VGND 0.28426f
C31089 a_54108_12568# VGND 0.28426f
C31090 a_53660_12568# VGND 0.28426f
C31091 a_53212_12568# VGND 0.28776f
C31092 a_60292_12612# VGND 0.47512f
C31093 a_59844_12612# VGND 0.46295f
C31094 a_59396_12612# VGND 0.46562f
C31095 a_58948_12612# VGND 0.49531f
C31096 a_58500_12612# VGND 0.46588f
C31097 a_58052_12612# VGND 0.45787f
C31098 a_57604_12612# VGND 0.45666f
C31099 a_57156_12612# VGND 0.45666f
C31100 a_56708_12612# VGND 0.47155f
C31101 a_56260_12612# VGND 0.45794f
C31102 a_55812_12612# VGND 0.4579f
C31103 a_55364_12612# VGND 0.4579f
C31104 a_54916_12612# VGND 0.4579f
C31105 a_54468_12612# VGND 0.4579f
C31106 a_54020_12612# VGND 0.4579f
C31107 a_53572_12612# VGND 0.4579f
C31108 a_53124_12612# VGND 0.46986f
C31109 a_52540_12568# VGND 0.29292f
C31110 a_52092_12568# VGND 0.29279f
C31111 a_51644_12568# VGND 0.29158f
C31112 a_51196_12568# VGND 0.31814f
C31113 a_50748_12568# VGND 0.29396f
C31114 a_50300_12568# VGND 0.2841f
C31115 a_49852_12568# VGND 0.2841f
C31116 a_49404_12568# VGND 0.2841f
C31117 a_48956_12568# VGND 0.28575f
C31118 a_48508_12568# VGND 0.28236f
C31119 a_48060_12568# VGND 0.28236f
C31120 a_47612_12568# VGND 0.28236f
C31121 a_47164_12568# VGND 0.28236f
C31122 a_46716_12568# VGND 0.28236f
C31123 a_46268_12568# VGND 0.28236f
C31124 a_45820_12568# VGND 0.28236f
C31125 a_45372_12568# VGND 0.29228f
C31126 a_52452_12612# VGND 0.47398f
C31127 a_52004_12612# VGND 0.46192f
C31128 a_51556_12612# VGND 0.46474f
C31129 a_51108_12612# VGND 0.50076f
C31130 a_50660_12612# VGND 0.46148f
C31131 a_50212_12612# VGND 0.45666f
C31132 a_49764_12612# VGND 0.45666f
C31133 a_49316_12612# VGND 0.45666f
C31134 a_48868_12612# VGND 0.47155f
C31135 a_48420_12612# VGND 0.44029f
C31136 a_47972_12612# VGND 0.44029f
C31137 a_47524_12612# VGND 0.44029f
C31138 a_47076_12612# VGND 0.44029f
C31139 a_46628_12612# VGND 0.44029f
C31140 a_46180_12612# VGND 0.44029f
C31141 a_45732_12612# VGND 0.44029f
C31142 a_45284_12612# VGND 0.46832f
C31143 a_5052_12568# VGND 0.28654f
C31144 a_4604_12568# VGND 0.31699f
C31145 a_4156_12568# VGND 0.29553f
C31146 a_3708_12568# VGND 0.2812f
C31147 a_3260_12568# VGND 0.2812f
C31148 a_2812_12568# VGND 0.2812f
C31149 a_2364_12568# VGND 0.2812f
C31150 a_1916_12568# VGND 0.2812f
C31151 a_1468_12568# VGND 0.2812f
C31152 a_1020_12568# VGND 0.29134f
C31153 a_4964_12612# VGND 0.47812f
C31154 a_4516_12612# VGND 0.5182f
C31155 a_4068_12612# VGND 0.44538f
C31156 a_3620_12612# VGND 0.43828f
C31157 a_3172_12612# VGND 0.43828f
C31158 a_2724_12612# VGND 0.43828f
C31159 a_2276_12612# VGND 0.43828f
C31160 a_1828_12612# VGND 0.43828f
C31161 a_1380_12612# VGND 0.43828f
C31162 a_932_12612# VGND 0.4664f
C31163 a_68020_13800# VGND 0.47855f
C31164 a_67572_13800# VGND 0.46105f
C31165 a_67124_13800# VGND 0.46383f
C31166 a_66676_13800# VGND 0.49822f
C31167 a_66228_13800# VGND 0.46128f
C31168 a_65780_13800# VGND 0.45589f
C31169 a_65332_13800# VGND 0.45589f
C31170 a_64884_13800# VGND 0.46795f
C31171 a_64212_13800# VGND 0.47057f
C31172 a_63764_13800# VGND 0.45666f
C31173 a_63316_13800# VGND 0.45666f
C31174 a_62868_13800# VGND 0.45666f
C31175 a_62420_13800# VGND 0.45666f
C31176 a_61972_13800# VGND 0.45666f
C31177 a_61524_13800# VGND 0.45666f
C31178 a_61076_13800# VGND 0.45666f
C31179 a_60628_13800# VGND 0.47293f
C31180 a_60180_13800# VGND 0.46151f
C31181 a_59732_13800# VGND 0.46339f
C31182 a_59284_13800# VGND 0.46634f
C31183 a_58836_13800# VGND 0.49982f
C31184 a_58388_13800# VGND 0.46146f
C31185 a_57940_13800# VGND 0.4579f
C31186 a_57492_13800# VGND 0.4579f
C31187 a_57044_13800# VGND 0.46986f
C31188 a_56372_13800# VGND 0.47057f
C31189 a_55924_13800# VGND 0.45666f
C31190 a_55476_13800# VGND 0.45666f
C31191 a_55028_13800# VGND 0.45666f
C31192 a_54580_13800# VGND 0.45666f
C31193 a_54132_13800# VGND 0.45666f
C31194 a_53684_13800# VGND 0.45666f
C31195 a_53236_13800# VGND 0.45666f
C31196 a_52788_13800# VGND 0.47351f
C31197 a_52340_13800# VGND 0.46174f
C31198 a_51892_13800# VGND 0.46372f
C31199 a_51444_13800# VGND 0.46721f
C31200 a_50996_13800# VGND 0.49018f
C31201 a_50548_13800# VGND 0.45994f
C31202 a_50100_13800# VGND 0.4579f
C31203 a_49652_13800# VGND 0.4579f
C31204 a_49204_13800# VGND 0.4724f
C31205 a_48420_13800# VGND 0.44215f
C31206 a_47972_13800# VGND 0.43828f
C31207 a_47524_13800# VGND 0.43828f
C31208 a_47076_13800# VGND 0.43828f
C31209 a_46628_13800# VGND 0.43828f
C31210 a_46180_13800# VGND 0.43828f
C31211 a_45732_13800# VGND 0.43828f
C31212 a_45284_13800# VGND 0.4664f
C31213 a_5300_13800# VGND 0.48995f
C31214 a_4852_13800# VGND 0.48956f
C31215 a_4068_13800# VGND 0.44997f
C31216 a_3620_13800# VGND 0.43828f
C31217 a_3172_13800# VGND 0.43828f
C31218 a_2724_13800# VGND 0.43828f
C31219 a_2276_13800# VGND 0.43828f
C31220 a_1828_13800# VGND 0.43828f
C31221 a_1380_13800# VGND 0.43828f
C31222 a_932_13800# VGND 0.4664f
C31223 a_68108_13703# VGND 0.31354f
C31224 a_67660_13703# VGND 0.28994f
C31225 a_67212_13703# VGND 0.2922f
C31226 a_66764_13703# VGND 0.31659f
C31227 a_66316_13703# VGND 0.29504f
C31228 a_65868_13703# VGND 0.28481f
C31229 a_65420_13703# VGND 0.28481f
C31230 a_64972_13703# VGND 0.28853f
C31231 a_64300_13703# VGND 0.28981f
C31232 a_63852_13703# VGND 0.28793f
C31233 a_63404_13703# VGND 0.28445f
C31234 a_62956_13703# VGND 0.28445f
C31235 a_62508_13703# VGND 0.28445f
C31236 a_62060_13703# VGND 0.28445f
C31237 a_61612_13703# VGND 0.28445f
C31238 a_61164_13703# VGND 0.28445f
C31239 a_60716_13703# VGND 0.28924f
C31240 a_60268_13703# VGND 0.28596f
C31241 a_59820_13703# VGND 0.2878f
C31242 a_59372_13703# VGND 0.29011f
C31243 a_58924_13703# VGND 0.32081f
C31244 a_58476_13703# VGND 0.29043f
C31245 a_58028_13703# VGND 0.28825f
C31246 a_57580_13703# VGND 0.28443f
C31247 a_57132_13703# VGND 0.28949f
C31248 a_56460_13703# VGND 0.29109f
C31249 a_56012_13703# VGND 0.28921f
C31250 a_55564_13703# VGND 0.28573f
C31251 a_55116_13703# VGND 0.28573f
C31252 a_54668_13703# VGND 0.28573f
C31253 a_54220_13703# VGND 0.28573f
C31254 a_53772_13703# VGND 0.28573f
C31255 a_53324_13703# VGND 0.28583f
C31256 a_52876_13703# VGND 0.28873f
C31257 a_52428_13703# VGND 0.28981f
C31258 a_51980_13703# VGND 0.29173f
C31259 a_51532_13703# VGND 0.29421f
C31260 a_51084_13703# VGND 0.33375f
C31261 a_50636_13703# VGND 0.29182f
C31262 a_50188_13703# VGND 0.28597f
C31263 a_49740_13703# VGND 0.28597f
C31264 a_49292_13703# VGND 0.28834f
C31265 a_48508_13703# VGND 0.26958f
C31266 a_48060_13703# VGND 0.2812f
C31267 a_47612_13703# VGND 0.2812f
C31268 a_47164_13703# VGND 0.2812f
C31269 a_46716_13703# VGND 0.2812f
C31270 a_46268_13703# VGND 0.2812f
C31271 a_45820_13703# VGND 0.2812f
C31272 a_45372_13703# VGND 0.29134f
C31273 a_5388_13703# VGND 0.3139f
C31274 a_4940_13703# VGND 0.29949f
C31275 a_4156_13703# VGND 0.28278f
C31276 a_3708_13703# VGND 0.2812f
C31277 a_3260_13703# VGND 0.2812f
C31278 a_2812_13703# VGND 0.2812f
C31279 a_2364_13703# VGND 0.2812f
C31280 a_1916_13703# VGND 0.2812f
C31281 a_1468_13703# VGND 0.2812f
C31282 a_1020_13703# VGND 0.29134f
C31283 a_67772_14136# VGND 0.28307f
C31284 a_67324_14136# VGND 0.29092f
C31285 a_66876_14136# VGND 0.30126f
C31286 a_66428_14136# VGND 0.30744f
C31287 a_65980_14136# VGND 0.28416f
C31288 a_65532_14136# VGND 0.2841f
C31289 a_65084_14136# VGND 0.2841f
C31290 a_64636_14136# VGND 0.28575f
C31291 a_64188_14136# VGND 0.28427f
C31292 a_63740_14136# VGND 0.28426f
C31293 a_63292_14136# VGND 0.28426f
C31294 a_62844_14136# VGND 0.28426f
C31295 a_62396_14136# VGND 0.28426f
C31296 a_61948_14136# VGND 0.28426f
C31297 a_61500_14136# VGND 0.28426f
C31298 a_61052_14136# VGND 0.28799f
C31299 a_67684_14180# VGND 0.45149f
C31300 a_67236_14180# VGND 0.44741f
C31301 a_66788_14180# VGND 0.46978f
C31302 a_66340_14180# VGND 0.44909f
C31303 a_65892_14180# VGND 0.44029f
C31304 a_65444_14180# VGND 0.44029f
C31305 a_64996_14180# VGND 0.44029f
C31306 a_64548_14180# VGND 0.47263f
C31307 a_64100_14180# VGND 0.4732f
C31308 a_63652_14180# VGND 0.4732f
C31309 a_63204_14180# VGND 0.4732f
C31310 a_62756_14180# VGND 0.4732f
C31311 a_62308_14180# VGND 0.4732f
C31312 a_61860_14180# VGND 0.47322f
C31313 a_61412_14180# VGND 0.4721f
C31314 a_60964_14180# VGND 0.48726f
C31315 a_60268_14136# VGND 0.27391f
C31316 a_59820_14136# VGND 0.28953f
C31317 a_59372_14136# VGND 0.29185f
C31318 a_58924_14136# VGND 0.32321f
C31319 a_57692_14136# VGND 0.26067f
C31320 a_57244_14136# VGND 0.28845f
C31321 a_56796_14136# VGND 0.28923f
C31322 a_56348_14136# VGND 0.28659f
C31323 a_55900_14136# VGND 0.2831f
C31324 a_55452_14136# VGND 0.2831f
C31325 a_55004_14136# VGND 0.2831f
C31326 a_54556_14136# VGND 0.2831f
C31327 a_54108_14136# VGND 0.2831f
C31328 a_53660_14136# VGND 0.2831f
C31329 a_53212_14136# VGND 0.28681f
C31330 a_60180_14180# VGND 0.46695f
C31331 a_59732_14180# VGND 0.47743f
C31332 a_59284_14180# VGND 0.47095f
C31333 a_58836_14180# VGND 0.5046f
C31334 a_57604_14180# VGND 0.46418f
C31335 a_57156_14180# VGND 0.47964f
C31336 a_56708_14180# VGND 0.44748f
C31337 a_56260_14180# VGND 0.43828f
C31338 a_55812_14180# VGND 0.43828f
C31339 a_55364_14180# VGND 0.43828f
C31340 a_54916_14180# VGND 0.43828f
C31341 a_54468_14180# VGND 0.43828f
C31342 a_54020_14180# VGND 0.43828f
C31343 a_53572_14180# VGND 0.43828f
C31344 a_53124_14180# VGND 0.48023f
C31345 a_52540_14136# VGND 0.29292f
C31346 a_52092_14136# VGND 0.29279f
C31347 a_51644_14136# VGND 0.29158f
C31348 a_51196_14136# VGND 0.31814f
C31349 a_50748_14136# VGND 0.29396f
C31350 a_50300_14136# VGND 0.2841f
C31351 a_49852_14136# VGND 0.2841f
C31352 a_49404_14136# VGND 0.2841f
C31353 a_48956_14136# VGND 0.28575f
C31354 a_48508_14136# VGND 0.28236f
C31355 a_48060_14136# VGND 0.28236f
C31356 a_47612_14136# VGND 0.28236f
C31357 a_47164_14136# VGND 0.28236f
C31358 a_46716_14136# VGND 0.28236f
C31359 a_46268_14136# VGND 0.28236f
C31360 a_45820_14136# VGND 0.28236f
C31361 a_45372_14136# VGND 0.29228f
C31362 a_52452_14180# VGND 0.45761f
C31363 a_52004_14180# VGND 0.44555f
C31364 a_51556_14180# VGND 0.44837f
C31365 a_51108_14180# VGND 0.48342f
C31366 a_50660_14180# VGND 0.44511f
C31367 a_50212_14180# VGND 0.44029f
C31368 a_49764_14180# VGND 0.44029f
C31369 a_49316_14180# VGND 0.47263f
C31370 a_48868_14180# VGND 0.4732f
C31371 a_48420_14180# VGND 0.4732f
C31372 a_47972_14180# VGND 0.4732f
C31373 a_47524_14180# VGND 0.4732f
C31374 a_47076_14180# VGND 0.4732f
C31375 a_46628_14180# VGND 0.4732f
C31376 a_46180_14180# VGND 0.47322f
C31377 a_45732_14180# VGND 0.47141f
C31378 a_45284_14180# VGND 0.46912f
C31379 a_5052_14136# VGND 0.28654f
C31380 a_4604_14136# VGND 0.31699f
C31381 a_4156_14136# VGND 0.29553f
C31382 a_3708_14136# VGND 0.2812f
C31383 a_3260_14136# VGND 0.2812f
C31384 a_2812_14136# VGND 0.2812f
C31385 a_2364_14136# VGND 0.2812f
C31386 a_1916_14136# VGND 0.2812f
C31387 a_1468_14136# VGND 0.2812f
C31388 a_1020_14136# VGND 0.29134f
C31389 a_4964_14180# VGND 0.47812f
C31390 a_4516_14180# VGND 0.5182f
C31391 a_4068_14180# VGND 0.44538f
C31392 a_3620_14180# VGND 0.43828f
C31393 a_3172_14180# VGND 0.43828f
C31394 a_2724_14180# VGND 0.43828f
C31395 a_2276_14180# VGND 0.43828f
C31396 a_1828_14180# VGND 0.43828f
C31397 a_1380_14180# VGND 0.43828f
C31398 a_932_14180# VGND 0.4664f
C31399 a_67684_15368# VGND 0.46156f
C31400 a_67236_15368# VGND 0.4546f
C31401 a_66788_15368# VGND 0.47695f
C31402 a_66340_15368# VGND 0.45244f
C31403 a_65892_15368# VGND 0.44364f
C31404 a_65444_15368# VGND 0.44364f
C31405 a_64996_15368# VGND 0.45546f
C31406 a_64324_15368# VGND 0.47393f
C31407 a_63876_15368# VGND 0.4701f
C31408 a_63428_15368# VGND 0.4701f
C31409 a_62980_15368# VGND 0.4701f
C31410 a_62532_15368# VGND 0.4701f
C31411 a_62084_15368# VGND 0.4701f
C31412 a_61636_15368# VGND 0.4701f
C31413 a_61188_15368# VGND 0.48746f
C31414 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.I VGND 1.4832f
C31415 a_56708_15368# VGND 0.44276f
C31416 a_56260_15368# VGND 0.43828f
C31417 a_55812_15368# VGND 0.43828f
C31418 a_55364_15368# VGND 0.43828f
C31419 a_54916_15368# VGND 0.43828f
C31420 a_54468_15368# VGND 0.43828f
C31421 a_54020_15368# VGND 0.43828f
C31422 a_53572_15368# VGND 0.45034f
C31423 a_52900_15368# VGND 0.47558f
C31424 a_52452_15368# VGND 0.44169f
C31425 a_52004_15368# VGND 0.44354f
C31426 a_51556_15368# VGND 0.44636f
C31427 a_51108_15368# VGND 0.48142f
C31428 a_50660_15368# VGND 0.4431f
C31429 a_50212_15368# VGND 0.43828f
C31430 a_49764_15368# VGND 0.45034f
C31431 a_49092_15368# VGND 0.47397f
C31432 a_48644_15368# VGND 0.47117f
C31433 a_48196_15368# VGND 0.4712f
C31434 a_47748_15368# VGND 0.4712f
C31435 a_47300_15368# VGND 0.4712f
C31436 a_46852_15368# VGND 0.4712f
C31437 a_46404_15368# VGND 0.4712f
C31438 a_45956_15368# VGND 0.48325f
C31439 a_45284_15368# VGND 0.44211f
C31440 a_44836_15368# VGND 0.474f
C31441 a_44388_15368# VGND 0.47965f
C31442 a_43940_15368# VGND 0.48206f
C31443 a_43492_15368# VGND 0.50285f
C31444 a_43044_15368# VGND 0.48625f
C31445 a_42596_15368# VGND 0.47513f
C31446 a_42148_15368# VGND 0.48718f
C31447 a_41476_15368# VGND 0.47896f
C31448 a_41028_15368# VGND 0.47513f
C31449 a_40580_15368# VGND 0.47513f
C31450 a_40132_15368# VGND 0.47513f
C31451 a_39684_15368# VGND 0.47513f
C31452 a_39236_15368# VGND 0.47513f
C31453 a_38788_15368# VGND 0.47513f
C31454 a_38340_15368# VGND 0.48718f
C31455 a_37668_15368# VGND 0.47896f
C31456 a_37220_15368# VGND 0.47727f
C31457 a_36772_15368# VGND 0.47901f
C31458 a_36324_15368# VGND 0.48106f
C31459 a_35876_15368# VGND 0.48476f
C31460 a_35428_15368# VGND 0.50799f
C31461 a_34980_15368# VGND 0.47673f
C31462 a_34532_15368# VGND 0.48718f
C31463 a_33860_15368# VGND 0.47896f
C31464 a_33412_15368# VGND 0.47513f
C31465 a_32964_15368# VGND 0.47513f
C31466 a_32516_15368# VGND 0.47513f
C31467 a_32068_15368# VGND 0.47513f
C31468 a_31620_15368# VGND 0.47513f
C31469 a_31172_15368# VGND 0.47513f
C31470 a_30724_15368# VGND 0.50325f
C31471 a_5300_15368# VGND 0.48995f
C31472 a_4852_15368# VGND 0.48956f
C31473 a_4068_15368# VGND 0.44997f
C31474 a_3620_15368# VGND 0.43828f
C31475 a_3172_15368# VGND 0.43828f
C31476 a_2724_15368# VGND 0.43828f
C31477 a_2276_15368# VGND 0.43828f
C31478 a_1828_15368# VGND 0.43828f
C31479 a_1380_15368# VGND 0.43828f
C31480 a_932_15368# VGND 0.4664f
C31481 a_67772_15271# VGND 0.28748f
C31482 a_67324_15271# VGND 0.29851f
C31483 a_66876_15271# VGND 0.30871f
C31484 a_66428_15271# VGND 0.31368f
C31485 a_65980_15271# VGND 0.28914f
C31486 a_65532_15271# VGND 0.289f
C31487 a_65084_15271# VGND 0.29217f
C31488 a_64412_15271# VGND 0.28628f
C31489 a_63964_15271# VGND 0.2812f
C31490 a_63516_15271# VGND 0.2812f
C31491 a_63068_15271# VGND 0.2812f
C31492 a_62620_15271# VGND 0.2812f
C31493 a_62172_15271# VGND 0.2812f
C31494 a_61724_15271# VGND 0.28611f
C31495 a_61276_15271# VGND 0.28908f
C31496 vgaringosc.tapped_ring.c13_inv_array\[30\]_pdkinv_notouch_.ZN VGND 1.08658f
C31497 vgaringosc.tapped_ring.c13_inv_array\[31\]_pdkinv_notouch_.ZN VGND 1.02457f
C31498 vgaringosc.tapped_ring.c13_inv_array\[32\]_pdkinv_notouch_.ZN VGND 0.87901f
C31499 a_56796_15271# VGND 0.28764f
C31500 a_56348_15271# VGND 0.28307f
C31501 a_55900_15271# VGND 0.287f
C31502 a_55452_15271# VGND 0.28549f
C31503 a_55004_15271# VGND 0.28611f
C31504 a_54556_15271# VGND 0.2861f
C31505 a_54108_15271# VGND 0.2862f
C31506 a_53660_15271# VGND 0.28492f
C31507 a_52988_15271# VGND 0.29137f
C31508 a_52540_15271# VGND 0.28964f
C31509 a_52092_15271# VGND 0.29139f
C31510 a_51644_15271# VGND 0.29366f
C31511 a_51196_15271# VGND 0.32145f
C31512 a_50748_15271# VGND 0.29606f
C31513 a_50300_15271# VGND 0.28618f
C31514 a_49852_15271# VGND 0.28981f
C31515 a_49180_15271# VGND 0.28628f
C31516 a_48732_15271# VGND 0.2812f
C31517 a_48284_15271# VGND 0.2812f
C31518 a_47836_15271# VGND 0.2812f
C31519 a_47388_15271# VGND 0.2812f
C31520 a_46940_15271# VGND 0.2812f
C31521 a_46492_15271# VGND 0.2812f
C31522 a_46044_15271# VGND 0.28983f
C31523 a_45372_15271# VGND 0.28628f
C31524 a_44924_15271# VGND 0.2842f
C31525 a_44476_15271# VGND 0.28571f
C31526 a_44028_15271# VGND 0.28788f
C31527 a_43580_15271# VGND 0.2953f
C31528 a_43132_15271# VGND 0.30806f
C31529 a_42684_15271# VGND 0.2814f
C31530 a_42236_15271# VGND 0.28492f
C31531 a_41564_15271# VGND 0.29117f
C31532 a_41116_15271# VGND 0.2861f
C31533 a_40668_15271# VGND 0.2861f
C31534 a_40220_15271# VGND 0.2861f
C31535 a_39772_15271# VGND 0.2861f
C31536 a_39324_15271# VGND 0.2861f
C31537 a_38876_15271# VGND 0.2861f
C31538 a_38428_15271# VGND 0.2899f
C31539 a_37756_15271# VGND 0.29127f
C31540 a_37308_15271# VGND 0.28766f
C31541 a_36860_15271# VGND 0.29008f
C31542 a_36412_15271# VGND 0.29204f
C31543 a_35964_15271# VGND 0.2946f
C31544 a_35516_15271# VGND 0.33265f
C31545 a_35068_15271# VGND 0.2914f
C31546 a_34620_15271# VGND 0.28989f
C31547 a_33948_15271# VGND 0.28628f
C31548 a_33500_15271# VGND 0.2812f
C31549 a_33052_15271# VGND 0.2812f
C31550 a_32604_15271# VGND 0.2812f
C31551 a_32156_15271# VGND 0.2812f
C31552 a_31708_15271# VGND 0.2812f
C31553 a_31260_15271# VGND 0.2812f
C31554 a_30812_15271# VGND 0.29134f
C31555 a_5388_15271# VGND 0.3139f
C31556 a_4940_15271# VGND 0.29949f
C31557 a_4156_15271# VGND 0.28278f
C31558 a_3708_15271# VGND 0.2812f
C31559 a_3260_15271# VGND 0.2812f
C31560 a_2812_15271# VGND 0.2812f
C31561 a_2364_15271# VGND 0.2812f
C31562 a_1916_15271# VGND 0.2812f
C31563 a_1468_15271# VGND 0.2812f
C31564 a_1020_15271# VGND 0.29134f
C31565 a_67996_15704# VGND 0.29582f
C31566 a_67548_15704# VGND 0.29777f
C31567 a_67100_15704# VGND 0.29973f
C31568 a_66652_15704# VGND 0.33923f
C31569 a_66204_15704# VGND 0.29688f
C31570 a_65756_15704# VGND 0.29036f
C31571 a_65308_15704# VGND 0.28964f
C31572 a_64860_15704# VGND 0.28756f
C31573 a_64412_15704# VGND 0.2812f
C31574 a_63964_15704# VGND 0.2812f
C31575 a_63516_15704# VGND 0.2812f
C31576 a_63068_15704# VGND 0.2812f
C31577 a_62620_15704# VGND 0.2812f
C31578 a_62172_15704# VGND 0.28515f
C31579 a_67908_15748# VGND 0.47462f
C31580 a_67460_15748# VGND 0.46957f
C31581 a_67012_15748# VGND 0.46899f
C31582 a_66564_15748# VGND 0.49515f
C31583 a_66116_15748# VGND 0.46251f
C31584 a_65668_15748# VGND 0.4749f
C31585 a_65220_15748# VGND 0.45593f
C31586 a_64772_15748# VGND 0.45593f
C31587 a_64324_15748# VGND 0.45588f
C31588 a_63876_15748# VGND 0.45588f
C31589 a_63428_15748# VGND 0.45588f
C31590 a_62980_15748# VGND 0.45588f
C31591 a_62532_15748# VGND 0.45588f
C31592 a_62084_15748# VGND 0.47048f
C31593 a_61388_15704# VGND 0.27283f
C31594 a_60940_15704# VGND 0.29175f
C31595 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.I VGND 0.86769f
C31596 vgaringosc.tapped_ring.c13_inv_array\[29\]_pdkinv_notouch_.I VGND 0.95084f
C31597 a_55228_15704# VGND 0.26731f
C31598 a_54780_15704# VGND 0.29296f
C31599 a_54332_15704# VGND 0.29495f
C31600 a_61300_15748# VGND 0.45134f
C31601 a_60852_15748# VGND 0.47033f
C31602 vgaringosc.tapped_ring.c13_inv_array\[26\]_pdkinv_notouch_.ZN VGND 0.89352f
C31603 vgaringosc.tapped_ring.c13_inv_array\[28\]_pdkinv_notouch_.I VGND 0.94778f
C31604 vgaringosc.tapped_ring.c13_inv_array\[33\]_pdkinv_notouch_.ZN VGND 1.04558f
C31605 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.I VGND 0.85301f
C31606 vgaringosc.tapped_ring.c13_inv_array\[35\]_pdkinv_notouch_.ZN VGND 0.88716f
C31607 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.I VGND 0.88425f
C31608 a_55140_15748# VGND 0.48533f
C31609 a_54692_15748# VGND 0.46513f
C31610 a_54244_15748# VGND 0.47815f
C31611 a_53660_15704# VGND 0.28772f
C31612 a_53212_15704# VGND 0.28904f
C31613 a_52764_15704# VGND 0.29098f
C31614 a_52316_15704# VGND 0.29287f
C31615 a_51868_15704# VGND 0.29495f
C31616 a_51420_15704# VGND 0.29776f
C31617 a_50972_15704# VGND 0.32408f
C31618 a_50524_15704# VGND 0.29107f
C31619 a_50076_15704# VGND 0.28862f
C31620 a_49628_15704# VGND 0.28871f
C31621 a_49180_15704# VGND 0.28236f
C31622 a_48732_15704# VGND 0.28236f
C31623 a_48284_15704# VGND 0.28236f
C31624 a_47836_15704# VGND 0.28236f
C31625 a_47388_15704# VGND 0.28236f
C31626 a_46940_15704# VGND 0.28236f
C31627 a_46492_15704# VGND 0.28586f
C31628 a_53572_15748# VGND 0.47057f
C31629 a_53124_15748# VGND 0.45666f
C31630 a_52676_15748# VGND 0.45942f
C31631 a_52228_15748# VGND 0.4609f
C31632 a_51780_15748# VGND 0.46308f
C31633 a_51332_15748# VGND 0.47509f
C31634 a_50884_15748# VGND 0.47538f
C31635 a_50436_15748# VGND 0.45666f
C31636 a_49988_15748# VGND 0.47155f
C31637 a_49540_15748# VGND 0.45794f
C31638 a_49092_15748# VGND 0.4579f
C31639 a_48644_15748# VGND 0.4579f
C31640 a_48196_15748# VGND 0.4579f
C31641 a_47748_15748# VGND 0.4579f
C31642 a_47300_15748# VGND 0.4579f
C31643 a_46852_15748# VGND 0.4579f
C31644 a_46404_15748# VGND 0.46986f
C31645 a_45820_15704# VGND 0.29108f
C31646 a_45372_15704# VGND 0.28584f
C31647 a_44924_15704# VGND 0.28536f
C31648 a_44476_15704# VGND 0.28687f
C31649 a_44028_15704# VGND 0.28904f
C31650 a_43580_15704# VGND 0.29645f
C31651 a_43132_15704# VGND 0.3092f
C31652 a_42684_15704# VGND 0.28255f
C31653 a_42236_15704# VGND 0.28236f
C31654 a_41788_15704# VGND 0.28916f
C31655 a_41340_15704# VGND 0.28922f
C31656 a_40892_15704# VGND 0.28922f
C31657 a_40444_15704# VGND 0.28922f
C31658 a_39996_15704# VGND 0.28922f
C31659 a_39548_15704# VGND 0.28922f
C31660 a_39100_15704# VGND 0.28922f
C31661 a_38652_15704# VGND 0.29272f
C31662 a_45732_15748# VGND 0.47191f
C31663 a_45284_15748# VGND 0.45801f
C31664 a_44836_15748# VGND 0.46095f
C31665 a_44388_15748# VGND 0.46253f
C31666 a_43940_15748# VGND 0.46496f
C31667 a_43492_15748# VGND 0.48464f
C31668 a_43044_15748# VGND 0.46905f
C31669 a_42596_15748# VGND 0.45668f
C31670 a_42148_15748# VGND 0.4724f
C31671 a_41700_15748# VGND 0.45794f
C31672 a_41252_15748# VGND 0.4579f
C31673 a_40804_15748# VGND 0.45791f
C31674 a_40356_15748# VGND 0.45926f
C31675 a_39908_15748# VGND 0.45844f
C31676 a_39460_15748# VGND 0.45925f
C31677 a_39012_15748# VGND 0.45928f
C31678 a_38564_15748# VGND 0.47087f
C31679 a_37980_15704# VGND 0.29452f
C31680 a_37532_15704# VGND 0.2927f
C31681 a_37084_15704# VGND 0.2924f
C31682 a_36636_15704# VGND 0.29402f
C31683 a_36188_15704# VGND 0.29624f
C31684 a_35740_15704# VGND 0.31295f
C31685 a_35292_15704# VGND 0.30495f
C31686 a_34844_15704# VGND 0.28922f
C31687 a_34396_15704# VGND 0.28932f
C31688 a_33948_15704# VGND 0.28236f
C31689 a_33500_15704# VGND 0.28236f
C31690 a_33052_15704# VGND 0.28236f
C31691 a_32604_15704# VGND 0.28236f
C31692 a_32156_15704# VGND 0.28236f
C31693 a_31708_15704# VGND 0.28236f
C31694 a_31260_15704# VGND 0.28236f
C31695 a_30812_15704# VGND 0.29228f
C31696 a_37892_15748# VGND 0.47057f
C31697 a_37444_15748# VGND 0.45671f
C31698 a_36996_15748# VGND 0.45978f
C31699 a_36548_15748# VGND 0.46148f
C31700 a_36100_15748# VGND 0.46408f
C31701 a_35652_15748# VGND 0.49078f
C31702 a_35204_15748# VGND 0.46493f
C31703 a_34756_15748# VGND 0.45666f
C31704 a_34308_15748# VGND 0.47155f
C31705 a_33860_15748# VGND 0.44029f
C31706 a_33412_15748# VGND 0.44029f
C31707 a_32964_15748# VGND 0.44029f
C31708 a_32516_15748# VGND 0.44029f
C31709 a_32068_15748# VGND 0.44029f
C31710 a_31620_15748# VGND 0.44029f
C31711 a_31172_15748# VGND 0.44029f
C31712 a_30724_15748# VGND 0.46832f
C31713 a_5052_15704# VGND 0.28654f
C31714 a_4604_15704# VGND 0.31699f
C31715 a_4156_15704# VGND 0.29553f
C31716 a_3708_15704# VGND 0.2812f
C31717 a_3260_15704# VGND 0.2812f
C31718 a_2812_15704# VGND 0.2812f
C31719 a_2364_15704# VGND 0.2812f
C31720 a_1916_15704# VGND 0.2812f
C31721 a_1468_15704# VGND 0.2812f
C31722 a_1020_15704# VGND 0.29134f
C31723 a_4964_15748# VGND 0.47812f
C31724 a_4516_15748# VGND 0.5182f
C31725 a_4068_15748# VGND 0.44538f
C31726 a_3620_15748# VGND 0.43828f
C31727 a_3172_15748# VGND 0.43828f
C31728 a_2724_15748# VGND 0.43828f
C31729 a_2276_15748# VGND 0.43828f
C31730 a_1828_15748# VGND 0.43828f
C31731 a_1380_15748# VGND 0.43828f
C31732 a_932_15748# VGND 0.4664f
C31733 a_67796_16936# VGND 0.47918f
C31734 a_67348_16936# VGND 0.46787f
C31735 a_66900_16936# VGND 0.47687f
C31736 a_66452_16936# VGND 0.48229f
C31737 a_66004_16936# VGND 0.47345f
C31738 a_65332_16936# VGND 0.46796f
C31739 a_64884_16936# VGND 0.46413f
C31740 a_64436_16936# VGND 0.456f
C31741 a_63988_16936# VGND 0.456f
C31742 a_63540_16936# VGND 0.456f
C31743 a_63092_16936# VGND 0.456f
C31744 a_62644_16936# VGND 0.456f
C31745 a_62196_16936# VGND 0.456f
C31746 a_61748_16936# VGND 0.47089f
C31747 a_61300_16936# VGND 0.44836f
C31748 vgaringosc.tapped_ring.c13_inv_array\[25\]_pdkinv_notouch_.I VGND 1.20813f
C31749 a_58612_16936# VGND 0.49485f
C31750 a_58164_16936# VGND 0.47447f
C31751 a_57380_16936# VGND 0.48019f
C31752 a_54804_16936# VGND 0.46928f
C31753 a_54356_16936# VGND 0.46413f
C31754 a_53908_16936# VGND 0.48012f
C31755 a_53460_16936# VGND 0.45732f
C31756 a_53012_16936# VGND 0.45618f
C31757 a_52564_16936# VGND 0.45925f
C31758 a_52116_16936# VGND 0.46091f
C31759 a_51668_16936# VGND 0.46345f
C31760 a_51220_16936# VGND 0.48856f
C31761 a_50772_16936# VGND 0.46466f
C31762 a_50324_16936# VGND 0.46824f
C31763 a_49652_16936# VGND 0.47085f
C31764 a_49204_16936# VGND 0.45801f
C31765 a_48756_16936# VGND 0.45801f
C31766 a_48308_16936# VGND 0.45801f
C31767 a_47860_16936# VGND 0.45801f
C31768 a_47412_16936# VGND 0.45801f
C31769 a_46964_16936# VGND 0.45801f
C31770 a_46516_16936# VGND 0.45801f
C31771 a_46068_16936# VGND 0.4729f
C31772 a_45620_16936# VGND 0.45934f
C31773 a_45172_16936# VGND 0.45987f
C31774 a_44724_16936# VGND 0.46255f
C31775 a_44276_16936# VGND 0.46432f
C31776 a_43828_16936# VGND 0.46704f
C31777 a_43380_16936# VGND 0.49786f
C31778 a_42932_16936# VGND 0.46605f
C31779 a_42484_16936# VGND 0.47125f
C31780 a_41812_16936# VGND 0.47196f
C31781 a_41364_16936# VGND 0.45695f
C31782 a_40916_16936# VGND 0.45695f
C31783 a_40468_16936# VGND 0.45695f
C31784 a_40020_16936# VGND 0.45695f
C31785 a_39572_16936# VGND 0.45695f
C31786 a_39124_16936# VGND 0.45695f
C31787 a_38676_16936# VGND 0.45695f
C31788 a_38228_16936# VGND 0.47294f
C31789 a_37780_16936# VGND 0.45823f
C31790 a_37332_16936# VGND 0.45935f
C31791 a_36884_16936# VGND 0.46167f
C31792 a_36436_16936# VGND 0.46355f
C31793 a_35988_16936# VGND 0.46645f
C31794 a_35540_16936# VGND 0.503f
C31795 a_35092_16936# VGND 0.46245f
C31796 a_34644_16936# VGND 0.47269f
C31797 a_33860_16936# VGND 0.44215f
C31798 a_33412_16936# VGND 0.43828f
C31799 a_32964_16936# VGND 0.43828f
C31800 a_32516_16936# VGND 0.43828f
C31801 a_32068_16936# VGND 0.43828f
C31802 a_31620_16936# VGND 0.43828f
C31803 a_31172_16936# VGND 0.43828f
C31804 a_30724_16936# VGND 0.4664f
C31805 a_5300_16936# VGND 0.48995f
C31806 a_4852_16936# VGND 0.48956f
C31807 a_4068_16936# VGND 0.44997f
C31808 a_3620_16936# VGND 0.43828f
C31809 a_3172_16936# VGND 0.43828f
C31810 a_2724_16936# VGND 0.43828f
C31811 a_2276_16936# VGND 0.43828f
C31812 a_1828_16936# VGND 0.43828f
C31813 a_1380_16936# VGND 0.43828f
C31814 a_932_16936# VGND 0.4664f
C31815 a_67884_16839# VGND 0.28654f
C31816 a_67436_16839# VGND 0.29441f
C31817 a_66988_16839# VGND 0.29492f
C31818 a_66540_16839# VGND 0.3229f
C31819 a_66092_16839# VGND 0.29206f
C31820 a_65420_16839# VGND 0.2908f
C31821 a_64972_16839# VGND 0.28921f
C31822 a_64524_16839# VGND 0.28805f
C31823 a_64076_16839# VGND 0.28457f
C31824 a_63628_16839# VGND 0.28457f
C31825 a_63180_16839# VGND 0.28457f
C31826 a_62732_16839# VGND 0.28457f
C31827 a_62284_16839# VGND 0.28457f
C31828 a_61836_16839# VGND 0.28622f
C31829 a_61388_16839# VGND 0.28558f
C31830 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.ZN VGND 0.88209f
C31831 vgaringosc.tapped_ring.c13_inv_array\[24\]_pdkinv_notouch_.I VGND 0.99674f
C31832 a_58700_16839# VGND 0.29661f
C31833 a_58252_16839# VGND 0.293f
C31834 a_57468_16839# VGND 0.27541f
C31835 vgaringosc.tapped_ring.c13_inv_array\[37\]_pdkinv_notouch_.ZN VGND 1.13678f
C31836 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.I VGND 0.88014f
C31837 vgaringosc.tapped_ring.c13_inv_array\[39\]_pdkinv_notouch_.ZN VGND 0.89845f
C31838 a_54892_16839# VGND 0.25893f
C31839 a_54444_16839# VGND 0.28981f
C31840 a_53996_16839# VGND 0.28923f
C31841 a_53548_16839# VGND 0.28659f
C31842 a_53100_16839# VGND 0.2831f
C31843 a_52652_16839# VGND 0.28623f
C31844 a_52204_16839# VGND 0.28781f
C31845 a_51756_16839# VGND 0.29002f
C31846 a_51308_16839# VGND 0.30331f
C31847 a_50860_16839# VGND 0.30292f
C31848 a_50412_16839# VGND 0.28684f
C31849 a_49740_16839# VGND 0.29109f
C31850 a_49292_16839# VGND 0.28793f
C31851 a_48844_16839# VGND 0.28445f
C31852 a_48396_16839# VGND 0.28445f
C31853 a_47948_16839# VGND 0.28445f
C31854 a_47500_16839# VGND 0.28445f
C31855 a_47052_16839# VGND 0.28445f
C31856 a_46604_16839# VGND 0.28445f
C31857 a_46156_16839# VGND 0.28747f
C31858 a_45708_16839# VGND 0.28236f
C31859 a_45260_16839# VGND 0.28236f
C31860 a_44812_16839# VGND 0.28568f
C31861 a_44364_16839# VGND 0.28736f
C31862 a_43916_16839# VGND 0.29106f
C31863 a_43468_16839# VGND 0.3115f
C31864 a_43020_16839# VGND 0.295f
C31865 a_42572_16839# VGND 0.2861f
C31866 a_41900_16839# VGND 0.28773f
C31867 a_41452_16839# VGND 0.28584f
C31868 a_41004_16839# VGND 0.28273f
C31869 a_40556_16839# VGND 0.28405f
C31870 a_40108_16839# VGND 0.28236f
C31871 a_39660_16839# VGND 0.2884f
C31872 a_39212_16839# VGND 0.28475f
C31873 a_38764_16839# VGND 0.28436f
C31874 a_38316_16839# VGND 0.28646f
C31875 a_37868_16839# VGND 0.28456f
C31876 a_37420_16839# VGND 0.28508f
C31877 a_36972_16839# VGND 0.28941f
C31878 a_36524_16839# VGND 0.28957f
C31879 a_36076_16839# VGND 0.29186f
C31880 a_35628_16839# VGND 0.32069f
C31881 a_35180_16839# VGND 0.29346f
C31882 a_34732_16839# VGND 0.28799f
C31883 a_33948_16839# VGND 0.26958f
C31884 a_33500_16839# VGND 0.2812f
C31885 a_33052_16839# VGND 0.2812f
C31886 a_32604_16839# VGND 0.2812f
C31887 a_32156_16839# VGND 0.2812f
C31888 a_31708_16839# VGND 0.2812f
C31889 a_31260_16839# VGND 0.2812f
C31890 a_30812_16839# VGND 0.29134f
C31891 a_5388_16839# VGND 0.3139f
C31892 a_4940_16839# VGND 0.29949f
C31893 a_4156_16839# VGND 0.28278f
C31894 a_3708_16839# VGND 0.2812f
C31895 a_3260_16839# VGND 0.2812f
C31896 a_2812_16839# VGND 0.2812f
C31897 a_2364_16839# VGND 0.2812f
C31898 a_1916_16839# VGND 0.2812f
C31899 a_1468_16839# VGND 0.2812f
C31900 a_1020_16839# VGND 0.29134f
C31901 a_67996_17272# VGND 0.29154f
C31902 a_67548_17272# VGND 0.29324f
C31903 a_67100_17272# VGND 0.29521f
C31904 a_66652_17272# VGND 0.3331f
C31905 a_66204_17272# VGND 0.29235f
C31906 a_65756_17272# VGND 0.28749f
C31907 a_65308_17272# VGND 0.28528f
C31908 a_64860_17272# VGND 0.28311f
C31909 a_64412_17272# VGND 0.2831f
C31910 a_63964_17272# VGND 0.2831f
C31911 a_63516_17272# VGND 0.2831f
C31912 a_63068_17272# VGND 0.2831f
C31913 a_62620_17272# VGND 0.2831f
C31914 a_62172_17272# VGND 0.28681f
C31915 a_43664_17317# VGND 0.01257f
C31916 a_67908_17316# VGND 0.47462f
C31917 a_67460_17316# VGND 0.46957f
C31918 a_67012_17316# VGND 0.46899f
C31919 a_66564_17316# VGND 0.49515f
C31920 a_66116_17316# VGND 0.46251f
C31921 a_65668_17316# VGND 0.4749f
C31922 a_65220_17316# VGND 0.43828f
C31923 a_64772_17316# VGND 0.43828f
C31924 a_64324_17316# VGND 0.43828f
C31925 a_63876_17316# VGND 0.43828f
C31926 a_63428_17316# VGND 0.43828f
C31927 a_62980_17316# VGND 0.43828f
C31928 a_62532_17316# VGND 0.43828f
C31929 a_62084_17316# VGND 0.45034f
C31930 a_61500_17272# VGND 0.29186f
C31931 vgaringosc.tapped_ring.c13_inv_array\[22\]_pdkinv_notouch_.I VGND 0.88355f
C31932 a_58924_17272# VGND 0.30379f
C31933 a_58476_17272# VGND 0.30001f
C31934 a_58028_17272# VGND 0.28919f
C31935 a_57580_17272# VGND 0.28584f
C31936 a_57132_17272# VGND 0.28989f
C31937 a_56684_17272# VGND 0.28798f
C31938 a_61412_17316# VGND 0.49714f
C31939 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.ZN VGND 0.93358f
C31940 vgaringosc.tapped_ring.c13_inv_array\[20\]_pdkinv_notouch_.ZN VGND 0.8732f
C31941 a_58836_17316# VGND 0.52089f
C31942 a_58388_17316# VGND 0.48027f
C31943 a_57940_17316# VGND 0.47481f
C31944 a_57492_17316# VGND 0.44364f
C31945 a_57044_17316# VGND 0.44364f
C31946 a_56596_17316# VGND 0.45371f
C31947 vgaringosc.tapped_ring.c13_inv_array\[41\]_pdkinv_notouch_.ZN VGND 0.85633f
C31948 vgaringosc.tapped_ring.c13_inv_array\[40\]_pdkinv_notouch_.ZN VGND 0.86654f
C31949 vgaringosc.tapped_ring.c13_inv_array\[42\]_pdkinv_notouch_.ZN VGND 1.08112f
C31950 a_53660_17272# VGND 0.29462f
C31951 a_53212_17272# VGND 0.28758f
C31952 a_52764_17272# VGND 0.2865f
C31953 a_52316_17272# VGND 0.28835f
C31954 a_51868_17272# VGND 0.29044f
C31955 a_51420_17272# VGND 0.29324f
C31956 a_50972_17272# VGND 0.31916f
C31957 a_50524_17272# VGND 0.28655f
C31958 a_50076_17272# VGND 0.28575f
C31959 a_49628_17272# VGND 0.28427f
C31960 a_49180_17272# VGND 0.28426f
C31961 a_48732_17272# VGND 0.28426f
C31962 a_48284_17272# VGND 0.28426f
C31963 a_47836_17272# VGND 0.28426f
C31964 a_47388_17272# VGND 0.28426f
C31965 a_46940_17272# VGND 0.28426f
C31966 a_46492_17272# VGND 0.28799f
C31967 a_53572_17316# VGND 0.47417f
C31968 a_53124_17316# VGND 0.45805f
C31969 a_52676_17316# VGND 0.46039f
C31970 a_52228_17316# VGND 0.46188f
C31971 a_51780_17316# VGND 0.46309f
C31972 a_51332_17316# VGND 0.47511f
C31973 a_50884_17316# VGND 0.47682f
C31974 a_50436_17316# VGND 0.45666f
C31975 a_49988_17316# VGND 0.47155f
C31976 a_49540_17316# VGND 0.47091f
C31977 a_49092_17316# VGND 0.47247f
C31978 a_48644_17316# VGND 0.47266f
C31979 a_48196_17316# VGND 0.4721f
C31980 a_47748_17316# VGND 0.4721f
C31981 a_47300_17316# VGND 0.47214f
C31982 a_46852_17316# VGND 0.47204f
C31983 a_46404_17316# VGND 0.48766f
C31984 a_45708_17272# VGND 0.2703f
C31985 a_45260_17272# VGND 0.2841f
C31986 a_44812_17272# VGND 0.28741f
C31987 a_44364_17272# VGND 0.28967f
C31988 a_43932_17800# VGND 0.00263f
C31989 a_41968_17801# VGND 0.00146f
C31990 a_41040_17801# VGND 0.0017f
C31991 a_41432_17801# VGND 0.42088f
C31992 a_41536_17636# VGND 0.29983f
C31993 a_41048_17341# VGND 1.48247f
C31994 a_45620_17316# VGND 0.46649f
C31995 a_45172_17316# VGND 0.4675f
C31996 a_44724_17316# VGND 0.47414f
C31997 a_44276_17316# VGND 0.47312f
C31998 a_40644_17272# VGND 0.4603f
C31999 a_39324_17272# VGND 0.26477f
C32000 a_40040_17675# VGND 1.13857f
C32001 a_39236_17316# VGND 0.48653f
C32002 a_37980_17272# VGND 0.29193f
C32003 a_37532_17272# VGND 0.28758f
C32004 a_37084_17272# VGND 0.28728f
C32005 a_36636_17272# VGND 0.28889f
C32006 a_36188_17272# VGND 0.29112f
C32007 a_35740_17272# VGND 0.30622f
C32008 a_35292_17272# VGND 0.29982f
C32009 a_34844_17272# VGND 0.2841f
C32010 a_34396_17272# VGND 0.28575f
C32011 a_33948_17272# VGND 0.28236f
C32012 a_33500_17272# VGND 0.28236f
C32013 a_33052_17272# VGND 0.28236f
C32014 a_32604_17272# VGND 0.28236f
C32015 a_32156_17272# VGND 0.28236f
C32016 a_31708_17272# VGND 0.28236f
C32017 a_31260_17272# VGND 0.28236f
C32018 a_30812_17272# VGND 0.29228f
C32019 a_37892_17316# VGND 0.48518f
C32020 a_37444_17316# VGND 0.46739f
C32021 a_36996_17316# VGND 0.4672f
C32022 a_36548_17316# VGND 0.46148f
C32023 a_36100_17316# VGND 0.46409f
C32024 a_35652_17316# VGND 0.49086f
C32025 a_35204_17316# VGND 0.46522f
C32026 a_34756_17316# VGND 0.45801f
C32027 a_34308_17316# VGND 0.47155f
C32028 a_33860_17316# VGND 0.44029f
C32029 a_33412_17316# VGND 0.44029f
C32030 a_32964_17316# VGND 0.44029f
C32031 a_32516_17316# VGND 0.44029f
C32032 a_32068_17316# VGND 0.44029f
C32033 a_31620_17316# VGND 0.44029f
C32034 a_31172_17316# VGND 0.44029f
C32035 a_30724_17316# VGND 0.46832f
C32036 a_5052_17272# VGND 0.28654f
C32037 a_4604_17272# VGND 0.31699f
C32038 a_4156_17272# VGND 0.29553f
C32039 a_3708_17272# VGND 0.2812f
C32040 a_3260_17272# VGND 0.2812f
C32041 a_2812_17272# VGND 0.2812f
C32042 a_2364_17272# VGND 0.2812f
C32043 a_1916_17272# VGND 0.2812f
C32044 a_1468_17272# VGND 0.2812f
C32045 a_1020_17272# VGND 0.29134f
C32046 a_4964_17316# VGND 0.47812f
C32047 a_4516_17316# VGND 0.5182f
C32048 a_4068_17316# VGND 0.44538f
C32049 a_3620_17316# VGND 0.43828f
C32050 a_3172_17316# VGND 0.43828f
C32051 a_2724_17316# VGND 0.43828f
C32052 a_2276_17316# VGND 0.43828f
C32053 a_1828_17316# VGND 0.43828f
C32054 a_1380_17316# VGND 0.43828f
C32055 a_932_17316# VGND 0.4664f
C32056 a_67796_18504# VGND 0.47889f
C32057 a_67348_18504# VGND 0.46758f
C32058 a_66900_18504# VGND 0.47658f
C32059 a_66452_18504# VGND 0.48183f
C32060 a_66004_18504# VGND 0.4757f
C32061 a_65220_18504# VGND 0.45423f
C32062 a_64772_18504# VGND 0.43828f
C32063 a_64324_18504# VGND 0.43828f
C32064 a_63876_18504# VGND 0.43828f
C32065 a_63428_18504# VGND 0.43828f
C32066 a_62980_18504# VGND 0.43828f
C32067 a_62532_18504# VGND 0.43828f
C32068 a_62084_18504# VGND 0.43828f
C32069 a_61636_18504# VGND 0.47963f
C32070 vgaringosc.tapped_ring.c13_inv_array\[19\]_pdkinv_notouch_.I VGND 1.08829f
C32071 a_58164_18504# VGND 0.49665f
C32072 a_44704_18191# VGND 0.00184f
C32073 a_43776_18191# VGND 0.0017f
C32074 a_57492_18504# VGND 0.4542f
C32075 a_57044_18504# VGND 0.44748f
C32076 a_56596_18504# VGND 0.45755f
C32077 a_54804_18504# VGND 0.46192f
C32078 a_54356_18504# VGND 0.47671f
C32079 a_53908_18504# VGND 0.47874f
C32080 a_53460_18504# VGND 0.45594f
C32081 a_53012_18504# VGND 0.45589f
C32082 a_52564_18504# VGND 0.45896f
C32083 a_52116_18504# VGND 0.46062f
C32084 a_51668_18504# VGND 0.46316f
C32085 a_51220_18504# VGND 0.48765f
C32086 a_50772_18504# VGND 0.46437f
C32087 a_50324_18504# VGND 0.47364f
C32088 a_49316_18504# VGND 0.4864f
C32089 a_48868_18504# VGND 0.4701f
C32090 a_48420_18504# VGND 0.4701f
C32091 a_47972_18504# VGND 0.4701f
C32092 a_47524_18504# VGND 0.4701f
C32093 a_47076_18504# VGND 0.4701f
C32094 a_46628_18504# VGND 0.4701f
C32095 a_46180_18504# VGND 0.47076f
C32096 a_45732_18504# VGND 0.46316f
C32097 a_43328_18559# VGND 0.00122f
C32098 a_67884_18407# VGND 0.28654f
C32099 a_67436_18407# VGND 0.29441f
C32100 a_66988_18407# VGND 0.29492f
C32101 a_66540_18407# VGND 0.3229f
C32102 a_66092_18407# VGND 0.2923f
C32103 a_65308_18407# VGND 0.27103f
C32104 a_64860_18407# VGND 0.28555f
C32105 a_64412_18407# VGND 0.2812f
C32106 a_63964_18407# VGND 0.2812f
C32107 a_63516_18407# VGND 0.2812f
C32108 a_63068_18407# VGND 0.2812f
C32109 a_62620_18407# VGND 0.2812f
C32110 a_62172_18407# VGND 0.2812f
C32111 a_61724_18407# VGND 0.28537f
C32112 vgaringosc.tapped_ring.c13_inv_array\[16\]_pdkinv_notouch_.ZN VGND 0.93616f
C32113 vgaringosc.tapped_ring.c13_inv_array\[17\]_pdkinv_notouch_.ZN VGND 0.98595f
C32114 a_58252_18407# VGND 0.27337f
C32115 a_57580_18407# VGND 0.28772f
C32116 a_57132_18407# VGND 0.28838f
C32117 a_56684_18407# VGND 0.2903f
C32118 vgaringosc.tapped_ring.c13_inv_array\[44\]_pdkinv_notouch_.ZN VGND 0.83824f
C32119 vgaringosc.tapped_ring.c13_inv_array\[43\]_pdkinv_notouch_.ZN VGND 1.11196f
C32120 a_54892_18407# VGND 0.27935f
C32121 a_54444_18407# VGND 0.28845f
C32122 a_53996_18407# VGND 0.29076f
C32123 a_53548_18407# VGND 0.28705f
C32124 a_53100_18407# VGND 0.28678f
C32125 a_52652_18407# VGND 0.28656f
C32126 a_52204_18407# VGND 0.28817f
C32127 a_51756_18407# VGND 0.29059f
C32128 a_51308_18407# VGND 0.301f
C32129 a_50860_18407# VGND 0.30331f
C32130 a_50412_18407# VGND 0.28549f
C32131 a_49404_18407# VGND 0.26874f
C32132 a_48956_18407# VGND 0.28555f
C32133 a_48508_18407# VGND 0.28722f
C32134 a_48060_18407# VGND 0.28479f
C32135 a_47612_18407# VGND 0.28374f
C32136 a_47164_18407# VGND 0.28329f
C32137 a_46716_18407# VGND 0.28526f
C32138 a_46268_18407# VGND 0.28702f
C32139 a_45820_18407# VGND 0.28149f
C32140 a_44752_18147# VGND 0.83649f
C32141 a_44459_18559# VGND 0.4687f
C32142 a_43452_18191# VGND 0.33052f
C32143 a_43824_18147# VGND 0.42187f
C32144 a_42896_18504# VGND 1.50376f
C32145 a_39216_18191# VGND 0.0017f
C32146 a_38288_18191# VGND 0.00146f
C32147 _452_.D VGND 0.87641f
C32148 _332_.Z VGND 0.51179f
C32149 a_40244_18180# VGND 1.12303f
C32150 a_39264_18147# VGND 0.84338f
C32151 a_38971_18559# VGND 0.46353f
C32152 a_37964_18191# VGND 0.30246f
C32153 a_38336_18147# VGND 0.42485f
C32154 _330_.ZN VGND 0.71283f
C32155 a_37408_18504# VGND 1.4802f
C32156 a_36436_18504# VGND 0.47672f
C32157 a_35988_18504# VGND 0.46951f
C32158 a_35540_18504# VGND 0.50567f
C32159 a_35092_18504# VGND 0.46551f
C32160 a_34644_18504# VGND 0.47561f
C32161 a_33860_18504# VGND 0.44215f
C32162 a_33412_18504# VGND 0.43828f
C32163 a_32964_18504# VGND 0.43828f
C32164 a_32516_18504# VGND 0.43828f
C32165 a_32068_18504# VGND 0.43828f
C32166 a_31620_18504# VGND 0.43828f
C32167 a_31172_18504# VGND 0.43828f
C32168 a_30724_18504# VGND 0.4664f
C32169 a_5300_18504# VGND 0.48995f
C32170 a_4852_18504# VGND 0.48956f
C32171 a_4068_18504# VGND 0.44997f
C32172 a_3620_18504# VGND 0.43828f
C32173 a_3172_18504# VGND 0.43828f
C32174 a_2724_18504# VGND 0.43828f
C32175 a_2276_18504# VGND 0.43828f
C32176 a_1828_18504# VGND 0.43828f
C32177 a_1380_18504# VGND 0.43828f
C32178 a_932_18504# VGND 0.4664f
C32179 a_36524_18407# VGND 0.25368f
C32180 a_36076_18407# VGND 0.29928f
C32181 a_35628_18407# VGND 0.3206f
C32182 a_35180_18407# VGND 0.29584f
C32183 a_34732_18407# VGND 0.29062f
C32184 a_33948_18407# VGND 0.26958f
C32185 a_33500_18407# VGND 0.2812f
C32186 a_33052_18407# VGND 0.2812f
C32187 a_32604_18407# VGND 0.2812f
C32188 a_32156_18407# VGND 0.2812f
C32189 a_31708_18407# VGND 0.2812f
C32190 a_31260_18407# VGND 0.2812f
C32191 a_30812_18407# VGND 0.29134f
C32192 a_5388_18407# VGND 0.3139f
C32193 a_4940_18407# VGND 0.29949f
C32194 a_4156_18407# VGND 0.28278f
C32195 a_3708_18407# VGND 0.2812f
C32196 a_3260_18407# VGND 0.2812f
C32197 a_2812_18407# VGND 0.2812f
C32198 a_2364_18407# VGND 0.2812f
C32199 a_1916_18407# VGND 0.2812f
C32200 a_1468_18407# VGND 0.2812f
C32201 a_1020_18407# VGND 0.29134f
C32202 a_67996_18840# VGND 0.29154f
C32203 a_67548_18840# VGND 0.29324f
C32204 a_67100_18840# VGND 0.29521f
C32205 a_66652_18840# VGND 0.3331f
C32206 a_66204_18840# VGND 0.29235f
C32207 a_65756_18840# VGND 0.28749f
C32208 a_65308_18840# VGND 0.28338f
C32209 a_64860_18840# VGND 0.2812f
C32210 a_64412_18840# VGND 0.2812f
C32211 a_63964_18840# VGND 0.2812f
C32212 a_63516_18840# VGND 0.2812f
C32213 a_63068_18840# VGND 0.2812f
C32214 a_62620_18840# VGND 0.2812f
C32215 a_62172_18840# VGND 0.28558f
C32216 a_51252_19001# VGND 0.00132f
C32217 a_67908_18884# VGND 0.47491f
C32218 a_67460_18884# VGND 0.47092f
C32219 a_67012_18884# VGND 0.46928f
C32220 a_66564_18884# VGND 0.49561f
C32221 a_66116_18884# VGND 0.4628f
C32222 a_65668_18884# VGND 0.4749f
C32223 a_65220_18884# VGND 0.43828f
C32224 a_64772_18884# VGND 0.43828f
C32225 a_64324_18884# VGND 0.43828f
C32226 a_63876_18884# VGND 0.43828f
C32227 a_63428_18884# VGND 0.43828f
C32228 a_62980_18884# VGND 0.43828f
C32229 a_62532_18884# VGND 0.43828f
C32230 a_62084_18884# VGND 0.45681f
C32231 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.I VGND 1.09492f
C32232 vgaringosc.tapped_ring.c13_inv_array\[15\]_pdkinv_notouch_.ZN VGND 0.88868f
C32233 a_58924_18840# VGND 0.30239f
C32234 a_58476_18840# VGND 0.29524f
C32235 a_58028_18840# VGND 0.28747f
C32236 a_57580_18840# VGND 0.28496f
C32237 a_54780_18840# VGND 0.26283f
C32238 a_54332_18840# VGND 0.29264f
C32239 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.ZN VGND 0.9733f
C32240 vgaringosc.tapped_ring.c13_inv_array\[14\]_pdkinv_notouch_.ZN VGND 0.98892f
C32241 a_58836_18884# VGND 0.50621f
C32242 a_58388_18884# VGND 0.47551f
C32243 a_57940_18884# VGND 0.47353f
C32244 a_57492_18884# VGND 0.48387f
C32245 vgaringosc.tapped_ring.c13_inv_array\[46\]_pdkinv_notouch_.ZN VGND 0.86714f
C32246 vgaringosc.tapped_ring.c13_inv_array\[45\]_pdkinv_notouch_.ZN VGND 0.88397f
C32247 a_54692_18884# VGND 0.46858f
C32248 a_54244_18884# VGND 0.48115f
C32249 a_53436_18840# VGND 0.27154f
C32250 a_51308_19369# VGND 0.00143f
C32251 a_50816_19369# VGND 0.00171f
C32252 a_49888_19369# VGND 0.0017f
C32253 a_52228_19368# VGND 0.49585f
C32254 a_50280_19369# VGND 0.42645f
C32255 a_50384_19204# VGND 0.31364f
C32256 a_49896_18909# VGND 1.5176f
C32257 a_53348_18884# VGND 0.48702f
C32258 a_49492_18840# VGND 0.45394f
C32259 a_48172_18840# VGND 0.2626f
C32260 a_47724_18840# VGND 0.28863f
C32261 a_43344_19001# VGND 0.00135f
C32262 a_48888_19243# VGND 1.1175f
C32263 a_48084_18884# VGND 0.46295f
C32264 a_47636_18884# VGND 0.47121f
C32265 a_45820_18840# VGND 0.29271f
C32266 a_40416_18885# VGND 0.00492f
C32267 a_44320_19369# VGND 0.00166f
C32268 a_43392_19369# VGND 0.00269f
C32269 _325_.ZN VGND 0.81221f
C32270 a_43784_19369# VGND 0.42892f
C32271 a_43888_19204# VGND 0.3047f
C32272 a_43400_18909# VGND 1.48952f
C32273 a_45732_18884# VGND 0.49264f
C32274 a_42996_18840# VGND 0.49515f
C32275 a_42392_19243# VGND 1.14191f
C32276 a_41188_18840# VGND 1.14206f
C32277 a_40684_19368# VGND 0.00255f
C32278 _331_.ZN VGND 0.66596f
C32279 a_39648_19435# VGND 0.00376f
C32280 _330_.A2 VGND 0.49418f
C32281 a_38644_19368# VGND 0.7352f
C32282 a_39268_18840# VGND 0.66406f
C32283 a_37312_19369# VGND 0.00174f
C32284 a_36384_19369# VGND 0.00168f
C32285 a_37067_19001# VGND 0.45904f
C32286 a_37360_19325# VGND 0.84311f
C32287 a_36060_19369# VGND 0.30498f
C32288 a_36432_19325# VGND 0.4261f
C32289 a_35504_18955# VGND 1.51647f
C32290 a_34396_18840# VGND 0.2603f
C32291 a_33948_18840# VGND 0.28555f
C32292 a_33500_18840# VGND 0.2812f
C32293 a_33052_18840# VGND 0.2812f
C32294 a_32604_18840# VGND 0.2812f
C32295 a_32156_18840# VGND 0.2812f
C32296 a_31708_18840# VGND 0.2812f
C32297 a_31260_18840# VGND 0.2812f
C32298 a_30812_18840# VGND 0.29134f
C32299 a_34308_18884# VGND 0.48611f
C32300 a_33860_18884# VGND 0.43828f
C32301 a_33412_18884# VGND 0.43828f
C32302 a_32964_18884# VGND 0.43828f
C32303 a_32516_18884# VGND 0.43828f
C32304 a_32068_18884# VGND 0.43828f
C32305 a_31620_18884# VGND 0.43828f
C32306 a_31172_18884# VGND 0.43828f
C32307 a_30724_18884# VGND 0.4664f
C32308 a_5052_18840# VGND 0.28654f
C32309 a_4604_18840# VGND 0.31699f
C32310 a_4156_18840# VGND 0.29553f
C32311 a_3708_18840# VGND 0.2812f
C32312 a_3260_18840# VGND 0.2812f
C32313 a_2812_18840# VGND 0.2812f
C32314 a_2364_18840# VGND 0.2812f
C32315 a_1916_18840# VGND 0.2812f
C32316 a_1468_18840# VGND 0.2812f
C32317 a_1020_18840# VGND 0.29134f
C32318 a_4964_18884# VGND 0.47812f
C32319 a_4516_18884# VGND 0.5182f
C32320 a_4068_18884# VGND 0.44538f
C32321 a_3620_18884# VGND 0.43828f
C32322 a_3172_18884# VGND 0.43828f
C32323 a_2724_18884# VGND 0.43828f
C32324 a_2276_18884# VGND 0.43828f
C32325 a_1828_18884# VGND 0.43828f
C32326 a_1380_18884# VGND 0.43828f
C32327 a_932_18884# VGND 0.4664f
C32328 a_67796_20072# VGND 0.47889f
C32329 a_67348_20072# VGND 0.46758f
C32330 a_66900_20072# VGND 0.47658f
C32331 a_66452_20072# VGND 0.48183f
C32332 a_66004_20072# VGND 0.4757f
C32333 a_65220_20072# VGND 0.45134f
C32334 a_64772_20072# VGND 0.44748f
C32335 a_64324_20072# VGND 0.43828f
C32336 a_63876_20072# VGND 0.43828f
C32337 a_63428_20072# VGND 0.43828f
C32338 a_62980_20072# VGND 0.43828f
C32339 a_62532_20072# VGND 0.43828f
C32340 a_62084_20072# VGND 0.43828f
C32341 a_61636_20072# VGND 0.46817f
C32342 a_61188_20072# VGND 0.47758f
C32343 vgaringosc.tapped_ring.c13_inv_array\[12\]_pdkinv_notouch_.I VGND 1.07584f
C32344 a_52944_19759# VGND 0.00155f
C32345 a_52016_19759# VGND 0.0019f
C32346 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.I VGND 1.14585f
C32347 a_55252_20072# VGND 0.48077f
C32348 a_54804_20072# VGND 0.46384f
C32349 a_49672_19668# VGND 0.00568f
C32350 a_54356_20072# VGND 0.47231f
C32351 _424_.ZN VGND 0.49757f
C32352 a_67884_19975# VGND 0.28963f
C32353 a_67436_19975# VGND 0.29732f
C32354 a_66988_19975# VGND 0.29907f
C32355 a_66540_19975# VGND 0.32562f
C32356 a_66092_19975# VGND 0.29658f
C32357 a_65308_19975# VGND 0.27429f
C32358 a_64860_19975# VGND 0.28981f
C32359 a_64412_19975# VGND 0.28468f
C32360 a_63964_19975# VGND 0.28501f
C32361 a_63516_19975# VGND 0.28409f
C32362 a_63068_19975# VGND 0.28478f
C32363 a_62620_19975# VGND 0.28537f
C32364 a_62172_19975# VGND 0.28294f
C32365 a_61724_19975# VGND 0.28457f
C32366 a_61276_19975# VGND 0.28394f
C32367 vgaringosc.tapped_ring.c13_inv_array\[9\]_pdkinv_notouch_.ZN VGND 0.95191f
C32368 vgaringosc.tapped_ring.c13_inv_array\[10\]_pdkinv_notouch_.ZN VGND 0.89256f
C32369 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.ZN VGND 0.99614f
C32370 vgaringosc.tapped_ring.c13_inv_array\[50\]_pdkinv_notouch_.ZN VGND 0.85502f
C32371 vgaringosc.tapped_ring.c13_inv_array\[49\]_pdkinv_notouch_.ZN VGND 1.09467f
C32372 vgaringosc.tapped_ring.c13_inv_array\[47\]_pdkinv_notouch_.ZN VGND 0.97475f
C32373 a_55340_19975# VGND 0.26366f
C32374 a_54892_19975# VGND 0.2888f
C32375 a_54444_19975# VGND 0.28793f
C32376 a_52408_19759# VGND 0.4232f
C32377 a_52512_19715# VGND 0.29662f
C32378 a_52024_20083# VGND 1.4662f
C32379 a_51620_19911# VGND 0.47412f
C32380 a_49448_20072# VGND 0.00372f
C32381 a_47504_19759# VGND 0.0017f
C32382 a_46576_19759# VGND 0.00146f
C32383 a_44484_19668# VGND 0.0027f
C32384 a_43668_19668# VGND 0.65423f
C32385 a_43444_19668# VGND 0.00938f
C32386 a_42811_19668# VGND 0.0026f
C32387 a_51240_19624# VGND 0.88493f
C32388 a_48776_20204# VGND 0.7323f
C32389 a_47552_19715# VGND 0.83088f
C32390 a_47259_20127# VGND 0.44797f
C32391 a_46252_19759# VGND 0.29712f
C32392 a_46624_19715# VGND 0.42459f
C32393 _416_.ZN VGND 0.82765f
C32394 a_45696_20072# VGND 1.47341f
C32395 a_44276_20072# VGND 0.00867f
C32396 a_43892_20072# VGND 0.00105f
C32397 _325_.B VGND 1.06394f
C32398 a_37772_19759# VGND 0.00145f
C32399 _450_.D VGND 0.84441f
C32400 a_40580_20072# VGND 0.46444f
C32401 a_40132_20072# VGND 0.45712f
C32402 a_39684_20072# VGND 0.4673f
C32403 a_39236_20072# VGND 0.46618f
C32404 a_38788_20072# VGND 0.48095f
C32405 _328_.A2 VGND 0.79345f
C32406 _327_.Z VGND 1.95488f
C32407 a_40668_19975# VGND 0.26046f
C32408 a_40220_19975# VGND 0.28627f
C32409 a_39772_19975# VGND 0.2841f
C32410 a_39324_19975# VGND 0.28573f
C32411 a_38876_19975# VGND 0.28829f
C32412 a_37384_19624# VGND 0.57687f
C32413 a_36612_20072# VGND 0.00121f
C32414 _448_.D VGND 0.86547f
C32415 a_35716_20072# VGND 0.00406f
C32416 a_35492_20072# VGND 0.00318f
C32417 a_34644_20072# VGND 0.49698f
C32418 a_33860_20072# VGND 0.44215f
C32419 a_33412_20072# VGND 0.43828f
C32420 a_32964_20072# VGND 0.43828f
C32421 a_32516_20072# VGND 0.43828f
C32422 a_32068_20072# VGND 0.43828f
C32423 a_31620_20072# VGND 0.43828f
C32424 a_31172_20072# VGND 0.43828f
C32425 a_30724_20072# VGND 0.4664f
C32426 a_5300_20072# VGND 0.48995f
C32427 a_4852_20072# VGND 0.48956f
C32428 a_4068_20072# VGND 0.44997f
C32429 a_3620_20072# VGND 0.43828f
C32430 a_3172_20072# VGND 0.43828f
C32431 a_2724_20072# VGND 0.43828f
C32432 a_2276_20072# VGND 0.43828f
C32433 a_1828_20072# VGND 0.43828f
C32434 a_1380_20072# VGND 0.43828f
C32435 a_932_20072# VGND 0.4664f
C32436 _323_.A3 VGND 0.53506f
C32437 _325_.A2 VGND 3.20604f
C32438 a_34732_19975# VGND 0.25558f
C32439 a_33948_19975# VGND 0.27294f
C32440 a_33500_19975# VGND 0.28759f
C32441 a_33052_19975# VGND 0.28473f
C32442 a_32604_19975# VGND 0.28473f
C32443 a_32156_19975# VGND 0.28473f
C32444 a_31708_19975# VGND 0.28473f
C32445 a_31260_19975# VGND 0.28473f
C32446 a_30812_19975# VGND 0.29381f
C32447 a_5388_19975# VGND 0.3139f
C32448 a_4940_19975# VGND 0.29949f
C32449 a_4156_19975# VGND 0.28278f
C32450 a_3708_19975# VGND 0.2812f
C32451 a_3260_19975# VGND 0.2812f
C32452 a_2812_19975# VGND 0.2812f
C32453 a_2364_19975# VGND 0.2812f
C32454 a_1916_19975# VGND 0.2812f
C32455 a_1468_19975# VGND 0.2812f
C32456 a_1020_19975# VGND 0.29134f
C32457 a_68108_20408# VGND 0.31676f
C32458 a_68020_20452# VGND 0.50792f
C32459 a_67212_20408# VGND 0.27978f
C32460 a_66764_20408# VGND 0.32383f
C32461 a_66316_20408# VGND 0.30149f
C32462 a_67124_20452# VGND 0.47821f
C32463 a_66676_20452# VGND 0.51878f
C32464 a_66228_20452# VGND 0.47438f
C32465 a_63404_20408# VGND 0.27244f
C32466 a_62060_20408# VGND 0.26337f
C32467 a_61612_20408# VGND 0.29023f
C32468 a_61164_20408# VGND 0.28857f
C32469 vgaringosc.tapped_ring.c13_inv_array\[8\]_pdkinv_notouch_.I VGND 1.27131f
C32470 a_63316_20452# VGND 0.47433f
C32471 a_61972_20452# VGND 0.46921f
C32472 a_61524_20452# VGND 0.46634f
C32473 a_61076_20452# VGND 0.4881f
C32474 vgaringosc.tapped_ring.c13_inv_array\[6\]_pdkinv_notouch_.ZN VGND 0.93677f
C32475 a_58476_20408# VGND 0.27325f
C32476 a_58028_20408# VGND 0.28984f
C32477 a_51912_20452# VGND 0.00646f
C32478 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.ZN VGND 0.91099f
C32479 a_58388_20452# VGND 0.47158f
C32480 a_57940_20452# VGND 0.47344f
C32481 vgaringosc.tapped_ring.c13_inv_array\[52\]_pdkinv_notouch_.ZN VGND 0.9007f
C32482 vgaringosc.tapped_ring.c13_inv_array\[51\]_pdkinv_notouch_.ZN VGND 0.85545f
C32483 a_55228_20408# VGND 0.26175f
C32484 a_54780_20408# VGND 0.28601f
C32485 a_54332_20408# VGND 0.28601f
C32486 a_53884_20408# VGND 0.28806f
C32487 a_52997_20936# VGND 0.00252f
C32488 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.I VGND 0.97971f
C32489 a_55140_20452# VGND 0.47641f
C32490 a_54692_20452# VGND 0.47426f
C32491 a_54244_20452# VGND 0.47519f
C32492 a_53796_20452# VGND 0.48052f
C32493 a_52136_20936# VGND 0.00597f
C32494 _424_.B2 VGND 0.73837f
C32495 a_51240_20452# VGND 0.74114f
C32496 a_50748_20408# VGND 0.2649f
C32497 a_50300_20408# VGND 0.2901f
C32498 a_50660_20452# VGND 0.46604f
C32499 a_50212_20452# VGND 0.47186f
C32500 a_49068_20408# VGND 1.41754f
C32501 a_47728_20937# VGND 0.0017f
C32502 a_46800_20937# VGND 0.00146f
C32503 a_47483_20569# VGND 0.45794f
C32504 a_47776_20893# VGND 0.83625f
C32505 a_46476_20937# VGND 0.2957f
C32506 a_46848_20893# VGND 0.42219f
C32507 a_45920_20523# VGND 1.47354f
C32508 a_43380_20452# VGND 0.00659f
C32509 a_43156_20452# VGND 0.00117f
C32510 a_44491_20936# VGND 0.0027f
C32511 a_42252_20936# VGND 2.09847f
C32512 a_40668_20408# VGND 0.27481f
C32513 a_40220_20408# VGND 0.28671f
C32514 a_39772_20408# VGND 0.28568f
C32515 a_39333_20936# VGND 0.00278f
C32516 a_38764_20408# VGND 0.26583f
C32517 a_38316_20408# VGND 0.2902f
C32518 _319_.A2 VGND 0.64421f
C32519 a_40580_20452# VGND 0.47514f
C32520 a_40132_20452# VGND 0.46637f
C32521 a_39684_20452# VGND 0.45823f
C32522 a_38676_20452# VGND 0.46558f
C32523 a_38228_20452# VGND 0.48555f
C32524 a_35968_20937# VGND 0.00176f
C32525 a_35040_20937# VGND 0.00146f
C32526 a_35723_20569# VGND 0.48478f
C32527 a_36016_20893# VGND 0.83925f
C32528 a_34716_20937# VGND 0.30122f
C32529 a_35088_20893# VGND 0.43539f
C32530 _319_.ZN VGND 0.77228f
C32531 a_34160_20523# VGND 1.50217f
C32532 a_33164_20408# VGND 0.29052f
C32533 a_32716_20408# VGND 0.28457f
C32534 a_32268_20408# VGND 0.28457f
C32535 a_31820_20408# VGND 0.28457f
C32536 a_31372_20408# VGND 0.28457f
C32537 a_30924_20408# VGND 0.28457f
C32538 a_30476_20408# VGND 0.28765f
C32539 a_30028_20408# VGND 0.30712f
C32540 a_33076_20452# VGND 0.46169f
C32541 a_32628_20452# VGND 0.45724f
C32542 a_32180_20452# VGND 0.45589f
C32543 a_31732_20452# VGND 0.45589f
C32544 a_31284_20452# VGND 0.45589f
C32545 a_30836_20452# VGND 0.45589f
C32546 a_30388_20452# VGND 0.45589f
C32547 a_29940_20452# VGND 0.4693f
C32548 a_29356_20408# VGND 0.31154f
C32549 a_28908_20408# VGND 0.308f
C32550 a_28460_20408# VGND 0.31019f
C32551 a_28012_20408# VGND 0.32062f
C32552 a_27564_20408# VGND 0.32724f
C32553 a_27116_20408# VGND 0.30349f
C32554 a_26668_20408# VGND 0.30341f
C32555 a_26220_20408# VGND 0.30712f
C32556 a_29268_20452# VGND 0.46147f
C32557 a_28820_20452# VGND 0.45926f
C32558 a_28372_20452# VGND 0.46173f
C32559 a_27924_20452# VGND 0.48201f
C32560 a_27476_20452# VGND 0.46383f
C32561 a_27028_20452# VGND 0.45465f
C32562 a_26580_20452# VGND 0.45465f
C32563 a_26132_20452# VGND 0.4816f
C32564 a_25548_20408# VGND 0.30848f
C32565 a_25100_20408# VGND 0.30341f
C32566 a_24652_20408# VGND 0.30341f
C32567 a_24204_20408# VGND 0.30341f
C32568 a_23756_20408# VGND 0.30341f
C32569 a_23308_20408# VGND 0.30341f
C32570 a_22860_20408# VGND 0.30341f
C32571 a_22412_20408# VGND 0.30712f
C32572 a_25460_20452# VGND 0.45987f
C32573 a_25012_20452# VGND 0.45604f
C32574 a_24564_20452# VGND 0.45604f
C32575 a_24116_20452# VGND 0.45604f
C32576 a_23668_20452# VGND 0.45604f
C32577 a_23220_20452# VGND 0.45604f
C32578 a_22772_20452# VGND 0.45604f
C32579 a_22324_20452# VGND 0.46809f
C32580 a_21740_20408# VGND 0.31018f
C32581 a_21292_20408# VGND 0.30738f
C32582 a_20844_20408# VGND 0.30937f
C32583 a_20396_20408# VGND 0.312f
C32584 a_19948_20408# VGND 0.34662f
C32585 a_19500_20408# VGND 0.30798f
C32586 a_19052_20408# VGND 0.30341f
C32587 a_18604_20408# VGND 0.30712f
C32588 a_21652_20452# VGND 0.4634f
C32589 a_21204_20452# VGND 0.46119f
C32590 a_20756_20452# VGND 0.46327f
C32591 a_20308_20452# VGND 0.46718f
C32592 a_19860_20452# VGND 0.4832f
C32593 a_19412_20452# VGND 0.4584f
C32594 a_18964_20452# VGND 0.45724f
C32595 a_18516_20452# VGND 0.4693f
C32596 a_17932_20408# VGND 0.30848f
C32597 a_17484_20408# VGND 0.30341f
C32598 a_17036_20408# VGND 0.30341f
C32599 a_16588_20408# VGND 0.30341f
C32600 a_16140_20408# VGND 0.30341f
C32601 a_15692_20408# VGND 0.30341f
C32602 a_15244_20408# VGND 0.30341f
C32603 a_14796_20408# VGND 0.31355f
C32604 a_17844_20452# VGND 0.44211f
C32605 a_17396_20452# VGND 0.43828f
C32606 a_16948_20452# VGND 0.43828f
C32607 a_16500_20452# VGND 0.43828f
C32608 a_16052_20452# VGND 0.43828f
C32609 a_15604_20452# VGND 0.43828f
C32610 a_15156_20452# VGND 0.43828f
C32611 a_14708_20452# VGND 0.4664f
C32612 a_5052_20408# VGND 0.28654f
C32613 a_4604_20408# VGND 0.31699f
C32614 a_4156_20408# VGND 0.29553f
C32615 a_3708_20408# VGND 0.2812f
C32616 a_3260_20408# VGND 0.2812f
C32617 a_2812_20408# VGND 0.2812f
C32618 a_2364_20408# VGND 0.2812f
C32619 a_1916_20408# VGND 0.2812f
C32620 a_1468_20408# VGND 0.2812f
C32621 a_1020_20408# VGND 0.29134f
C32622 a_4964_20452# VGND 0.47812f
C32623 a_4516_20452# VGND 0.5182f
C32624 a_4068_20452# VGND 0.44538f
C32625 a_3620_20452# VGND 0.43828f
C32626 a_3172_20452# VGND 0.43828f
C32627 a_2724_20452# VGND 0.43828f
C32628 a_2276_20452# VGND 0.43828f
C32629 a_1828_20452# VGND 0.43828f
C32630 a_1380_20452# VGND 0.43828f
C32631 a_932_20452# VGND 0.4664f
C32632 a_67684_21640# VGND 0.49795f
C32633 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.I VGND 1.12659f
C32634 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.I VGND 1.13992f
C32635 a_52452_21236# VGND 0.50551f
C32636 a_52081_21236# VGND 0.00652f
C32637 a_51877_21236# VGND 0.00767f
C32638 a_49988_21236# VGND 0.5346f
C32639 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.I VGND 1.17247f
C32640 vgaringosc.tapped_ring.c13_inv_array\[5\]_pdkinv_notouch_.I VGND 1.26345f
C32641 a_58500_21640# VGND 0.48617f
C32642 a_55364_21640# VGND 0.4832f
C32643 a_54916_21640# VGND 0.47548f
C32644 a_54468_21640# VGND 0.47548f
C32645 a_54020_21640# VGND 0.47549f
C32646 a_53572_21640# VGND 0.48516f
C32647 a_67772_21543# VGND 0.28755f
C32648 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.ZN VGND 0.95238f
C32649 vgaringosc.tapped_ring.c12_inv_array\[25\]_pdkinv_notouch_.ZN VGND 1.02218f
C32650 vgaringosc.tapped_ring.c12_inv_array\[27\]_pdkinv_notouch_.I VGND 0.95534f
C32651 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.I VGND 0.89687f
C32652 vgaringosc.tapped_ring.c12_inv_array\[28\]_pdkinv_notouch_.ZN VGND 0.87987f
C32653 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.ZN VGND 1.0452f
C32654 vgaringosc.tapped_ring.c13_inv_array\[4\]_pdkinv_notouch_.I VGND 0.90323f
C32655 a_58588_21543# VGND 0.27526f
C32656 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.ZN VGND 1.11806f
C32657 vgaringosc.tapped_ring.c13_inv_array\[54\]_pdkinv_notouch_.ZN VGND 1.21811f
C32658 vgaringosc.tapped_ring.c13_inv_array\[56\]_pdkinv_notouch_.I VGND 0.93533f
C32659 a_55452_21543# VGND 0.25893f
C32660 a_55004_21543# VGND 0.28627f
C32661 a_54556_21543# VGND 0.2864f
C32662 a_54108_21543# VGND 0.2867f
C32663 a_53660_21543# VGND 0.28873f
C32664 _422_.ZN VGND 0.55278f
C32665 a_51108_21640# VGND 0.51531f
C32666 _474_.D VGND 0.86616f
C32667 a_48068_21236# VGND 0.00256f
C32668 a_47531_21258# VGND 0.00124f
C32669 a_46389_21236# VGND 0.00247f
C32670 a_45564_21236# VGND 0.00385f
C32671 a_45156_21236# VGND 0.00687f
C32672 a_44290_21236# VGND 0.00238f
C32673 _416_.A2 VGND 0.8949f
C32674 a_47860_21640# VGND 0.00492f
C32675 _475_.D VGND 1.12982f
C32676 a_47271_21640# VGND 0.04512f
C32677 a_43646_21236# VGND 0.0032f
C32678 a_43254_21236# VGND 0.00332f
C32679 a_51196_21543# VGND 0.27145f
C32680 _417_.Z VGND 0.72165f
C32681 _419_.Z VGND 1.96385f
C32682 a_42630_21236# VGND 0.00307f
C32683 a_44038_21236# VGND 0.66009f
C32684 a_43814_21236# VGND 0.75652f
C32685 a_39873_21236# VGND 0.00661f
C32686 a_39669_21236# VGND 0.00757f
C32687 a_39475_21236# VGND 0.00803f
C32688 a_38548_21327# VGND 0.00145f
C32689 a_36204_21327# VGND 0.00168f
C32690 a_40692_21640# VGND 0.46931f
C32691 a_40244_21640# VGND 0.46714f
C32692 a_42982_21730# VGND 0.97446f
C32693 a_42778_21812# VGND 0.75823f
C32694 a_42154_21236# VGND 0.77348f
C32695 a_40780_21543# VGND 0.26715f
C32696 a_40332_21543# VGND 0.28694f
C32697 a_38340_21327# VGND 0.5518f
C32698 a_37444_21640# VGND 0.47684f
C32699 a_36996_21640# VGND 0.48227f
C32700 a_36548_21640# VGND 0.47493f
C32701 _319_.A3 VGND 1.45823f
C32702 a_37532_21543# VGND 0.28866f
C32703 a_37084_21543# VGND 0.29339f
C32704 a_36636_21543# VGND 0.29309f
C32705 a_35816_21192# VGND 0.59927f
C32706 a_34308_21640# VGND 0.4867f
C32707 a_33636_21640# VGND 0.47955f
C32708 a_33188_21640# VGND 0.45805f
C32709 a_32740_21640# VGND 0.45805f
C32710 a_32292_21640# VGND 0.45805f
C32711 a_31844_21640# VGND 0.45805f
C32712 a_31396_21640# VGND 0.45805f
C32713 a_30948_21640# VGND 0.45805f
C32714 a_30500_21640# VGND 0.45805f
C32715 a_30052_21640# VGND 0.45848f
C32716 a_29604_21640# VGND 0.47558f
C32717 a_29156_21640# VGND 0.46304f
C32718 a_28708_21640# VGND 0.46484f
C32719 a_28260_21640# VGND 0.46761f
C32720 a_27812_21640# VGND 0.50235f
C32721 a_27364_21640# VGND 0.4654f
C32722 a_26916_21640# VGND 0.45971f
C32723 a_26468_21640# VGND 0.47167f
C32724 a_25796_21640# VGND 0.48871f
C32725 a_25348_21640# VGND 0.45971f
C32726 a_24900_21640# VGND 0.45971f
C32727 a_24452_21640# VGND 0.45971f
C32728 a_24004_21640# VGND 0.45971f
C32729 a_23556_21640# VGND 0.45971f
C32730 a_23108_21640# VGND 0.45971f
C32731 a_22660_21640# VGND 0.45971f
C32732 a_22212_21640# VGND 0.45971f
C32733 a_21764_21640# VGND 0.45981f
C32734 a_21316_21640# VGND 0.46203f
C32735 a_20868_21640# VGND 0.46394f
C32736 a_20420_21640# VGND 0.46688f
C32737 a_19972_21640# VGND 0.50223f
C32738 a_19524_21640# VGND 0.46219f
C32739 a_19076_21640# VGND 0.45848f
C32740 a_18628_21640# VGND 0.47298f
C32741 a_17844_21640# VGND 0.44215f
C32742 a_17396_21640# VGND 0.43828f
C32743 a_16948_21640# VGND 0.43828f
C32744 a_16500_21640# VGND 0.43828f
C32745 a_16052_21640# VGND 0.43828f
C32746 a_15604_21640# VGND 0.43828f
C32747 a_15156_21640# VGND 0.43828f
C32748 a_14708_21640# VGND 0.4664f
C32749 a_5300_21640# VGND 0.48995f
C32750 a_4852_21640# VGND 0.48956f
C32751 a_4068_21640# VGND 0.44997f
C32752 a_3620_21640# VGND 0.43828f
C32753 a_3172_21640# VGND 0.43828f
C32754 a_2724_21640# VGND 0.43828f
C32755 a_2276_21640# VGND 0.43828f
C32756 a_1828_21640# VGND 0.43828f
C32757 a_1380_21640# VGND 0.43828f
C32758 a_932_21640# VGND 0.4664f
C32759 a_34396_21543# VGND 0.24383f
C32760 a_33724_21543# VGND 0.29068f
C32761 a_33276_21543# VGND 0.28608f
C32762 a_32828_21543# VGND 0.28389f
C32763 a_32380_21543# VGND 0.2841f
C32764 a_31932_21543# VGND 0.2841f
C32765 a_31484_21543# VGND 0.2841f
C32766 a_31036_21543# VGND 0.2841f
C32767 a_30588_21543# VGND 0.2841f
C32768 a_30140_21543# VGND 0.28575f
C32769 a_29692_21543# VGND 0.28427f
C32770 a_29244_21543# VGND 0.28763f
C32771 a_28796_21543# VGND 0.28935f
C32772 a_28348_21543# VGND 0.29161f
C32773 a_27900_21543# VGND 0.31464f
C32774 a_27452_21543# VGND 0.29456f
C32775 a_27004_21543# VGND 0.28426f
C32776 a_26556_21543# VGND 0.28776f
C32777 a_25884_21543# VGND 0.28946f
C32778 a_25436_21543# VGND 0.28758f
C32779 a_24988_21543# VGND 0.2841f
C32780 a_24540_21543# VGND 0.2841f
C32781 a_24092_21543# VGND 0.2841f
C32782 a_23644_21543# VGND 0.2841f
C32783 a_23196_21543# VGND 0.2841f
C32784 a_22748_21543# VGND 0.2841f
C32785 a_22300_21543# VGND 0.28575f
C32786 a_21852_21543# VGND 0.28478f
C32787 a_21404_21543# VGND 0.28784f
C32788 a_20956_21543# VGND 0.28967f
C32789 a_20508_21543# VGND 0.29198f
C32790 a_20060_21543# VGND 0.32287f
C32791 a_19612_21543# VGND 0.29254f
C32792 a_19164_21543# VGND 0.28426f
C32793 a_18716_21543# VGND 0.28799f
C32794 a_17932_21543# VGND 0.26958f
C32795 a_17484_21543# VGND 0.2812f
C32796 a_17036_21543# VGND 0.2812f
C32797 a_16588_21543# VGND 0.2812f
C32798 a_16140_21543# VGND 0.2812f
C32799 a_15692_21543# VGND 0.2812f
C32800 a_15244_21543# VGND 0.2812f
C32801 a_14796_21543# VGND 0.29134f
C32802 a_5388_21543# VGND 0.3139f
C32803 a_4940_21543# VGND 0.29949f
C32804 a_4156_21543# VGND 0.28278f
C32805 a_3708_21543# VGND 0.2812f
C32806 a_3260_21543# VGND 0.2812f
C32807 a_2812_21543# VGND 0.2812f
C32808 a_2364_21543# VGND 0.2812f
C32809 a_1916_21543# VGND 0.2812f
C32810 a_1468_21543# VGND 0.2812f
C32811 a_1020_21543# VGND 0.29134f
C32812 a_67996_21976# VGND 0.29567f
C32813 vgaringosc.tapped_ring.c12_inv_array\[14\]_pdkinv_notouch_.I VGND 0.88994f
C32814 vgaringosc.tapped_ring.c12_inv_array\[17\]_pdkinv_notouch_.I VGND 0.85158f
C32815 vgaringosc.tapped_ring.c12_inv_array\[20\]_pdkinv_notouch_.I VGND 0.97878f
C32816 vgaringosc.tapped_ring.c12_inv_array\[24\]_pdkinv_notouch_.I VGND 0.93482f
C32817 a_62508_21976# VGND 0.26625f
C32818 a_67908_22020# VGND 0.50285f
C32819 vgaringosc.tapped_ring.c12_inv_array\[12\]_pdkinv_notouch_.I VGND 0.96349f
C32820 vgaringosc.tapped_ring.c12_inv_array\[13\]_pdkinv_notouch_.I VGND 0.93183f
C32821 vgaringosc.tapped_ring.c12_inv_array\[15\]_pdkinv_notouch_.ZN VGND 1.04068f
C32822 vgaringosc.tapped_ring.c12_inv_array\[18\]_pdkinv_notouch_.ZN VGND 0.96039f
C32823 vgaringosc.tapped_ring.c12_inv_array\[21\]_pdkinv_notouch_.ZN VGND 0.96074f
C32824 vgaringosc.tapped_ring.c12_inv_array\[23\]_pdkinv_notouch_.I VGND 0.89415f
C32825 a_62420_22020# VGND 0.4634f
C32826 vgaringosc.tapped_ring.c12_inv_array\[29\]_pdkinv_notouch_.ZN VGND 0.91261f
C32827 vgaringosc.tapped_ring.c13_inv_array\[2\]_pdkinv_notouch_.I VGND 0.99619f
C32828 a_59260_21976# VGND 0.26842f
C32829 a_55744_22505# VGND 0.00146f
C32830 a_54816_22505# VGND 0.0017f
C32831 _427_.ZN VGND 0.70054f
C32832 a_55208_22505# VGND 0.42486f
C32833 a_55312_22340# VGND 0.30199f
C32834 a_54824_22045# VGND 1.47217f
C32835 vgaringosc.tapped_ring.c13_inv_array\[1\]_pdkinv_notouch_.I VGND 0.97283f
C32836 a_59172_22020# VGND 0.47414f
C32837 vgaringosc.tapped_ring.c13_inv_array\[59\]_pdkinv_notouch_.ZN VGND 0.87792f
C32838 vgaringosc.tapped_ring.c13_inv_array\[58\]_pdkinv_notouch_.ZN VGND 0.86882f
C32839 vgaringosc.tapped_ring.c13_inv_array\[57\]_pdkinv_notouch_.ZN VGND 0.93562f
C32840 a_54420_21976# VGND 0.46279f
C32841 a_54040_22366# VGND 0.84312f
C32842 a_53003_22504# VGND 0.0028f
C32843 a_52434_22504# VGND 0.00734f
C32844 a_52240_22504# VGND 0.00554f
C32845 a_52036_22504# VGND 0.00613f
C32846 a_51618_22504# VGND 0.00209f
C32847 a_51414_22504# VGND 0.00242f
C32848 a_51220_22504# VGND 0.00439f
C32849 a_47524_22021# VGND 0.00492f
C32850 a_46352_22021# VGND 0.00492f
C32851 _424_.A1 VGND 1.71851f
C32852 _427_.B2 VGND 0.92392f
C32853 _281_.A1 VGND 1.62275f
C32854 _476_.Q VGND 2.19926f
C32855 _473_.Q VGND 2.10235f
C32856 _421_.B VGND 0.72669f
C32857 a_47732_22504# VGND 0.00255f
C32858 a_46620_22504# VGND 0.00256f
C32859 a_48529_22460# VGND 0.54966f
C32860 _475_.Q VGND 2.36141f
C32861 _416_.A3 VGND 1.01764f
C32862 a_43600_22504# VGND 0.00489f
C32863 a_43192_22504# VGND 0.00271f
C32864 a_42784_22504# VGND 0.00242f
C32865 a_42376_22504# VGND 0.00515f
C32866 a_37296_22020# VGND 0.00128f
C32867 a_42168_22504# VGND 3.73582f
C32868 _304_.ZN VGND 1.50698f
C32869 _327_.A2 VGND 2.50488f
C32870 a_40452_22504# VGND 0.00487f
C32871 a_39796_22504# VGND 0.6031f
C32872 _302_.Z VGND 1.25712f
C32873 _301_.Z VGND 0.407f
C32874 _300_.A2 VGND 0.96689f
C32875 _316_.A3 VGND 0.71745f
C32876 a_38576_22504# VGND 1.39362f
C32877 _317_.A2 VGND 1.41365f
C32878 a_36148_21976# VGND 1.16365f
C32879 a_34960_22505# VGND 0.0017f
C32880 a_34032_22505# VGND 0.00146f
C32881 a_34715_22137# VGND 0.46515f
C32882 a_35008_22461# VGND 0.89022f
C32883 a_33708_22505# VGND 0.30081f
C32884 a_34080_22461# VGND 0.42549f
C32885 _316_.ZN VGND 0.76316f
C32886 a_33152_22091# VGND 1.47856f
C32887 a_32268_21976# VGND 0.25116f
C32888 a_31820_21976# VGND 0.28817f
C32889 a_31372_21976# VGND 0.286f
C32890 a_30924_21976# VGND 0.286f
C32891 a_30476_21976# VGND 0.28918f
C32892 a_32180_22020# VGND 0.47136f
C32893 a_31732_22020# VGND 0.46125f
C32894 a_31284_22020# VGND 0.46125f
C32895 a_30836_22020# VGND 0.46125f
C32896 a_30388_22020# VGND 0.47307f
C32897 a_29804_21976# VGND 0.29118f
C32898 a_29356_21976# VGND 0.29063f
C32899 a_28908_21976# VGND 0.2887f
C32900 a_28460_21976# VGND 0.29089f
C32901 a_28012_21976# VGND 0.30056f
C32902 a_27564_21976# VGND 0.30832f
C32903 a_27116_21976# VGND 0.28418f
C32904 a_26668_21976# VGND 0.2841f
C32905 a_26220_21976# VGND 0.28575f
C32906 a_25772_21976# VGND 0.2859f
C32907 a_25324_21976# VGND 0.28589f
C32908 a_24876_21976# VGND 0.28589f
C32909 a_24428_21976# VGND 0.28589f
C32910 a_23980_21976# VGND 0.28589f
C32911 a_23532_21976# VGND 0.28589f
C32912 a_23084_21976# VGND 0.28589f
C32913 a_22636_21976# VGND 0.28939f
C32914 a_29716_22020# VGND 0.47057f
C32915 a_29268_22020# VGND 0.46057f
C32916 a_28820_22020# VGND 0.46206f
C32917 a_28372_22020# VGND 0.46374f
C32918 a_27924_22020# VGND 0.48549f
C32919 a_27476_22020# VGND 0.46584f
C32920 a_27028_22020# VGND 0.45666f
C32921 a_26580_22020# VGND 0.45666f
C32922 a_26132_22020# VGND 0.47155f
C32923 a_25684_22020# VGND 0.45794f
C32924 a_25236_22020# VGND 0.4579f
C32925 a_24788_22020# VGND 0.4579f
C32926 a_24340_22020# VGND 0.4579f
C32927 a_23892_22020# VGND 0.4579f
C32928 a_23444_22020# VGND 0.4579f
C32929 a_22996_22020# VGND 0.4579f
C32930 a_22548_22020# VGND 0.46986f
C32931 a_21964_21976# VGND 0.29114f
C32932 a_21516_21976# VGND 0.29253f
C32933 a_21068_21976# VGND 0.2907f
C32934 a_20620_21976# VGND 0.29294f
C32935 a_20172_21976# VGND 0.3107f
C32936 a_19724_21976# VGND 0.2982f
C32937 a_19276_21976# VGND 0.28581f
C32938 a_18828_21976# VGND 0.28581f
C32939 a_18380_21976# VGND 0.28879f
C32940 a_17932_21976# VGND 0.28236f
C32941 a_17484_21976# VGND 0.28236f
C32942 a_17036_21976# VGND 0.28236f
C32943 a_16588_21976# VGND 0.28236f
C32944 a_16140_21976# VGND 0.28236f
C32945 a_15692_21976# VGND 0.28236f
C32946 a_15244_21976# VGND 0.28236f
C32947 a_14796_21976# VGND 0.29228f
C32948 a_21876_22020# VGND 0.47083f
C32949 a_21428_22020# VGND 0.45984f
C32950 a_20980_22020# VGND 0.46157f
C32951 a_20532_22020# VGND 0.46423f
C32952 a_20084_22020# VGND 0.49306f
C32953 a_19636_22020# VGND 0.46467f
C32954 a_19188_22020# VGND 0.45666f
C32955 a_18740_22020# VGND 0.45666f
C32956 a_18292_22020# VGND 0.47155f
C32957 a_17844_22020# VGND 0.44029f
C32958 a_17396_22020# VGND 0.44029f
C32959 a_16948_22020# VGND 0.44029f
C32960 a_16500_22020# VGND 0.44029f
C32961 a_16052_22020# VGND 0.44029f
C32962 a_15604_22020# VGND 0.44029f
C32963 a_15156_22020# VGND 0.44029f
C32964 a_14708_22020# VGND 0.46832f
C32965 a_5052_21976# VGND 0.28654f
C32966 a_4604_21976# VGND 0.31699f
C32967 a_4156_21976# VGND 0.29553f
C32968 a_3708_21976# VGND 0.2812f
C32969 a_3260_21976# VGND 0.2812f
C32970 a_2812_21976# VGND 0.2812f
C32971 a_2364_21976# VGND 0.2812f
C32972 a_1916_21976# VGND 0.2812f
C32973 a_1468_21976# VGND 0.2812f
C32974 a_1020_21976# VGND 0.29134f
C32975 a_4964_22020# VGND 0.47812f
C32976 a_4516_22020# VGND 0.5182f
C32977 a_4068_22020# VGND 0.44538f
C32978 a_3620_22020# VGND 0.43828f
C32979 a_3172_22020# VGND 0.43828f
C32980 a_2724_22020# VGND 0.43828f
C32981 a_2276_22020# VGND 0.43828f
C32982 a_1828_22020# VGND 0.43828f
C32983 a_1380_22020# VGND 0.43828f
C32984 a_932_22020# VGND 0.4664f
C32985 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.I VGND 1.13598f
C32986 vgaringosc.tapped_ring.c12_inv_array\[10\]_pdkinv_notouch_.ZN VGND 1.00004f
C32987 a_65668_23208# VGND 0.49805f
C32988 a_64660_23208# VGND 0.46613f
C32989 a_64212_23208# VGND 0.47091f
C32990 a_63764_23208# VGND 0.45197f
C32991 a_63316_23208# VGND 0.44984f
C32992 a_62868_23208# VGND 0.46889f
C32993 a_62420_23208# VGND 0.43828f
C32994 a_61972_23208# VGND 0.45106f
C32995 a_61524_23208# VGND 0.47067f
C32996 a_61076_23208# VGND 0.47352f
C32997 a_59620_23208# VGND 0.48715f
C32998 a_59172_23208# VGND 0.46829f
C32999 a_54624_22895# VGND 0.00146f
C33000 a_53696_22895# VGND 0.0017f
C33001 a_56932_23208# VGND 0.48621f
C33002 a_56484_23208# VGND 0.46903f
C33003 a_56036_23208# VGND 0.47681f
C33004 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.ZN VGND 1.19776f
C33005 vgaringosc.tapped_ring.c12_inv_array\[9\]_pdkinv_notouch_.ZN VGND 1.23447f
C33006 a_65756_23111# VGND 0.26693f
C33007 a_64748_23111# VGND 0.26669f
C33008 a_64300_23111# VGND 0.28555f
C33009 a_63852_23111# VGND 0.2812f
C33010 a_63404_23111# VGND 0.2812f
C33011 a_62956_23111# VGND 0.2812f
C33012 a_62508_23111# VGND 0.28601f
C33013 a_62060_23111# VGND 0.28505f
C33014 a_61612_23111# VGND 0.28735f
C33015 a_61164_23111# VGND 0.28645f
C33016 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.I VGND 1.13968f
C33017 a_59708_23111# VGND 0.27278f
C33018 a_59260_23111# VGND 0.2957f
C33019 vgaringosc.tapped_ring.c13_inv_array\[61\]_pdkinv_notouch_.ZN VGND 0.88188f
C33020 vgaringosc.tapped_ring.c13_inv_array\[60\]_pdkinv_notouch_.ZN VGND 1.22044f
C33021 a_57020_23111# VGND 0.27015f
C33022 a_56572_23111# VGND 0.29023f
C33023 a_56124_23111# VGND 0.28945f
C33024 a_54088_22895# VGND 0.42145f
C33025 a_54192_22851# VGND 0.30301f
C33026 a_53704_23219# VGND 1.47612f
C33027 a_53300_23047# VGND 0.46685f
C33028 a_50196_22805# VGND 0.71236f
C33029 a_49405_22805# VGND 0.00499f
C33030 a_49013_22805# VGND 0.0022f
C33031 a_50732_23233# VGND 0.00111f
C33032 a_48321_23208# VGND 0.0582f
C33033 a_52920_22760# VGND 0.83616f
C33034 a_51240_23340# VGND 0.87835f
C33035 _395_.A3 VGND 0.65673f
C33036 _218_.ZN VGND 1.03755f
C33037 _399_.A1 VGND 0.85643f
C33038 _324_.B VGND 3.50172f
C33039 a_47860_23208# VGND 0.4894f
C33040 a_39780_22805# VGND 0.71078f
C33041 a_38529_22804# VGND 0.00648f
C33042 a_38325_22804# VGND 0.0075f
C33043 a_38131_22804# VGND 0.00823f
C33044 a_35188_22895# VGND 0.00167f
C33045 a_47948_23111# VGND 0.26368f
C33046 _438_.ZN VGND 0.83852f
C33047 _303_.ZN VGND 1.18524f
C33048 _301_.A1 VGND 2.61142f
C33049 a_36772_23208# VGND 0.48989f
C33050 a_36288_23208# VGND 0.00106f
C33051 a_36860_23111# VGND 0.28177f
C33052 _311_.Z VGND 1.2243f
C33053 a_34980_22895# VGND 0.60742f
C33054 _312_.ZN VGND 0.60096f
C33055 a_33636_23208# VGND 0.48488f
C33056 a_33188_23208# VGND 0.46734f
C33057 a_32740_23208# VGND 0.46406f
C33058 a_32292_23208# VGND 0.45666f
C33059 a_31844_23208# VGND 0.45666f
C33060 a_31396_23208# VGND 0.45666f
C33061 a_30948_23208# VGND 0.45666f
C33062 a_30500_23208# VGND 0.45666f
C33063 a_30052_23208# VGND 0.47155f
C33064 a_29604_23208# VGND 0.45872f
C33065 a_29156_23208# VGND 0.46123f
C33066 a_28708_23208# VGND 0.46303f
C33067 a_28260_23208# VGND 0.46579f
C33068 a_27812_23208# VGND 0.49961f
C33069 a_27364_23208# VGND 0.46359f
C33070 a_26916_23208# VGND 0.4579f
C33071 a_26468_23208# VGND 0.46986f
C33072 a_25796_23208# VGND 0.47057f
C33073 a_25348_23208# VGND 0.45666f
C33074 a_24900_23208# VGND 0.45666f
C33075 a_24452_23208# VGND 0.45666f
C33076 a_24004_23208# VGND 0.45666f
C33077 a_23556_23208# VGND 0.45666f
C33078 a_23108_23208# VGND 0.45666f
C33079 a_22660_23208# VGND 0.45666f
C33080 a_22212_23208# VGND 0.47155f
C33081 a_21764_23208# VGND 0.45927f
C33082 a_21316_23208# VGND 0.46144f
C33083 a_20868_23208# VGND 0.46336f
C33084 a_20420_23208# VGND 0.4663f
C33085 a_19972_23208# VGND 0.50071f
C33086 a_19524_23208# VGND 0.46161f
C33087 a_19076_23208# VGND 0.4579f
C33088 a_18628_23208# VGND 0.4724f
C33089 a_17844_23208# VGND 0.44215f
C33090 a_17396_23208# VGND 0.43828f
C33091 a_16948_23208# VGND 0.43828f
C33092 a_16500_23208# VGND 0.43828f
C33093 a_16052_23208# VGND 0.43828f
C33094 a_15604_23208# VGND 0.43828f
C33095 a_15156_23208# VGND 0.43828f
C33096 a_14708_23208# VGND 0.4664f
C33097 a_5300_23208# VGND 0.48995f
C33098 a_4852_23208# VGND 0.48956f
C33099 a_4068_23208# VGND 0.44997f
C33100 a_3620_23208# VGND 0.43828f
C33101 a_3172_23208# VGND 0.43828f
C33102 a_2724_23208# VGND 0.43828f
C33103 a_2276_23208# VGND 0.43828f
C33104 a_1828_23208# VGND 0.43828f
C33105 a_1380_23208# VGND 0.43828f
C33106 a_932_23208# VGND 0.4664f
C33107 a_33724_23111# VGND 0.29035f
C33108 a_33276_23111# VGND 0.28597f
C33109 a_32828_23111# VGND 0.28774f
C33110 a_32380_23111# VGND 0.28542f
C33111 a_31932_23111# VGND 0.28458f
C33112 a_31484_23111# VGND 0.28462f
C33113 a_31036_23111# VGND 0.28449f
C33114 a_30588_23111# VGND 0.28435f
C33115 a_30140_23111# VGND 0.28639f
C33116 a_29692_23111# VGND 0.2859f
C33117 a_29244_23111# VGND 0.28811f
C33118 a_28796_23111# VGND 0.28934f
C33119 a_28348_23111# VGND 0.29325f
C33120 a_27900_23111# VGND 0.3168f
C33121 a_27452_23111# VGND 0.29483f
C33122 a_27004_23111# VGND 0.28496f
C33123 a_26556_23111# VGND 0.28893f
C33124 a_25884_23111# VGND 0.28946f
C33125 a_25436_23111# VGND 0.28758f
C33126 a_24988_23111# VGND 0.2841f
C33127 a_24540_23111# VGND 0.2841f
C33128 a_24092_23111# VGND 0.2841f
C33129 a_23644_23111# VGND 0.2841f
C33130 a_23196_23111# VGND 0.2841f
C33131 a_22748_23111# VGND 0.2841f
C33132 a_22300_23111# VGND 0.28575f
C33133 a_21852_23111# VGND 0.28478f
C33134 a_21404_23111# VGND 0.28784f
C33135 a_20956_23111# VGND 0.28967f
C33136 a_20508_23111# VGND 0.29198f
C33137 a_20060_23111# VGND 0.32287f
C33138 a_19612_23111# VGND 0.29254f
C33139 a_19164_23111# VGND 0.28426f
C33140 a_18716_23111# VGND 0.28799f
C33141 a_17932_23111# VGND 0.26958f
C33142 a_17484_23111# VGND 0.2812f
C33143 a_17036_23111# VGND 0.2812f
C33144 a_16588_23111# VGND 0.2812f
C33145 a_16140_23111# VGND 0.2812f
C33146 a_15692_23111# VGND 0.2812f
C33147 a_15244_23111# VGND 0.2812f
C33148 a_14796_23111# VGND 0.29134f
C33149 a_5388_23111# VGND 0.3139f
C33150 a_4940_23111# VGND 0.29949f
C33151 a_4156_23111# VGND 0.28278f
C33152 a_3708_23111# VGND 0.2812f
C33153 a_3260_23111# VGND 0.2812f
C33154 a_2812_23111# VGND 0.2812f
C33155 a_2364_23111# VGND 0.2812f
C33156 a_1916_23111# VGND 0.2812f
C33157 a_1468_23111# VGND 0.2812f
C33158 a_1020_23111# VGND 0.29134f
C33159 vgaringosc.tapped_ring.c12_inv_array\[7\]_pdkinv_notouch_.I VGND 1.05877f
C33160 a_65644_23544# VGND 0.28093f
C33161 a_65196_23544# VGND 0.29012f
C33162 a_64748_23544# VGND 0.2854f
C33163 a_64300_23544# VGND 0.2841f
C33164 a_63852_23544# VGND 0.2841f
C33165 a_63404_23544# VGND 0.28476f
C33166 a_62284_23544# VGND 0.26755f
C33167 a_61836_23544# VGND 0.29278f
C33168 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.ZN VGND 0.94357f
C33169 a_65556_23588# VGND 0.46631f
C33170 a_65108_23588# VGND 0.46496f
C33171 a_64660_23588# VGND 0.47418f
C33172 a_64212_23588# VGND 0.47194f
C33173 a_63764_23588# VGND 0.46142f
C33174 a_63316_23588# VGND 0.46326f
C33175 a_62196_23588# VGND 0.47753f
C33176 a_61748_23588# VGND 0.48058f
C33177 a_59260_23544# VGND 0.27023f
C33178 _231_.I VGND 0.67462f
C33179 a_57580_23544# VGND 0.26258f
C33180 a_57132_23544# VGND 0.28444f
C33181 a_56684_23544# VGND 0.28459f
C33182 a_56236_23544# VGND 0.2833f
C33183 a_55788_23544# VGND 0.28422f
C33184 a_55340_23544# VGND 0.28146f
C33185 a_54892_23544# VGND 0.28259f
C33186 a_54444_23544# VGND 0.28408f
C33187 a_48308_23588# VGND 0.05674f
C33188 a_59172_23588# VGND 0.48434f
C33189 vgaringosc.tapped_ring.c13_inv_array\[62\]_pdkinv_notouch_.ZN VGND 0.95362f
C33190 a_57492_23588# VGND 0.47318f
C33191 a_57044_23588# VGND 0.46869f
C33192 a_56596_23588# VGND 0.45577f
C33193 a_56148_23588# VGND 0.43828f
C33194 a_55700_23588# VGND 0.43828f
C33195 a_55252_23588# VGND 0.43828f
C33196 a_54804_23588# VGND 0.43828f
C33197 a_54356_23588# VGND 0.44258f
C33198 _384_.A1 VGND 1.67413f
C33199 a_52660_24072# VGND 0.00157f
C33200 a_52452_24072# VGND 0.5596f
C33201 a_51988_24072# VGND 0.00566f
C33202 _427_.A2 VGND 0.9738f
C33203 a_51332_24072# VGND 0.62349f
C33204 a_50940_24072# VGND 0.00419f
C33205 a_50532_24072# VGND 0.00683f
C33206 a_48908_24080# VGND 0.00222f
C33207 _399_.A2 VGND 1.32558f
C33208 a_48516_24080# VGND 0.00488f
C33209 _417_.A2 VGND 2.57744f
C33210 _397_.Z VGND 0.74737f
C33211 a_46984_23588# VGND 0.86668f
C33212 _402_.B VGND 0.69021f
C33213 a_46356_24072# VGND 0.17297f
C33214 _399_.ZN VGND 2.20817f
C33215 a_44906_24164# VGND 0.00317f
C33216 a_44282_24164# VGND 0.00308f
C33217 a_43890_24164# VGND 0.00319f
C33218 a_43246_24163# VGND 0.00259f
C33219 _305_.A2 VGND 1.47121f
C33220 _226_.ZN VGND 0.83086f
C33221 a_44786_24120# VGND 0.75554f
C33222 a_44162_24120# VGND 0.75608f
C33223 a_43750_23544# VGND 0.94537f
C33224 a_43126_24119# VGND 0.76512f
C33225 a_42796_23981# VGND 0.67817f
C33226 a_41488_24072# VGND 1.37375f
C33227 _325_.A1 VGND 4.92053f
C33228 _300_.ZN VGND 0.75315f
C33229 _434_.ZN VGND 0.74008f
C33230 _441_.B VGND 0.47672f
C33231 a_38759_24072# VGND 0.00759f
C33232 a_38575_24072# VGND 0.00667f
C33233 _437_.ZN VGND 0.49264f
C33234 _439_.ZN VGND 0.99004f
C33235 a_37644_23544# VGND 0.29588f
C33236 a_37196_23544# VGND 0.2886f
C33237 a_36748_23544# VGND 0.29114f
C33238 a_36300_23544# VGND 0.29385f
C33239 _304_.A1 VGND 4.50507f
C33240 a_35184_24073# VGND 0.0019f
C33241 a_34256_24073# VGND 0.00146f
C33242 a_37556_23588# VGND 0.46398f
C33243 a_37108_23588# VGND 0.47036f
C33244 a_36660_23588# VGND 0.47261f
C33245 a_36212_23588# VGND 0.48002f
C33246 a_34939_23705# VGND 0.48247f
C33247 a_35232_24029# VGND 0.88347f
C33248 a_33932_24073# VGND 0.30188f
C33249 a_34304_24029# VGND 0.42246f
C33250 _313_.ZN VGND 0.84695f
C33251 a_33376_23659# VGND 1.47109f
C33252 a_32268_23544# VGND 0.25877f
C33253 a_31820_23544# VGND 0.28817f
C33254 a_31372_23544# VGND 0.286f
C33255 a_30924_23544# VGND 0.286f
C33256 a_30476_23544# VGND 0.28918f
C33257 a_32180_23588# VGND 0.4701f
C33258 a_31732_23588# VGND 0.46759f
C33259 a_31284_23588# VGND 0.46839f
C33260 a_30836_23588# VGND 0.46736f
C33261 a_30388_23588# VGND 0.47826f
C33262 a_29804_23544# VGND 0.28994f
C33263 a_29028_24072# VGND 0.00147f
C33264 a_29716_23588# VGND 0.48572f
C33265 a_28820_24072# VGND 0.56622f
C33266 a_28460_23544# VGND 0.24963f
C33267 a_28012_23544# VGND 0.304f
C33268 a_27564_23544# VGND 0.31133f
C33269 a_27116_23544# VGND 0.28591f
C33270 a_26668_23544# VGND 0.28584f
C33271 a_26220_23544# VGND 0.28749f
C33272 a_25772_23544# VGND 0.28528f
C33273 a_25324_23544# VGND 0.2831f
C33274 a_24876_23544# VGND 0.2831f
C33275 a_24428_23544# VGND 0.2831f
C33276 a_23980_23544# VGND 0.2831f
C33277 a_23532_23544# VGND 0.2831f
C33278 a_23084_23544# VGND 0.2831f
C33279 a_22636_23544# VGND 0.28681f
C33280 a_28372_23588# VGND 0.47249f
C33281 a_27924_23588# VGND 0.47629f
C33282 a_27476_23588# VGND 0.46907f
C33283 a_27028_23588# VGND 0.45593f
C33284 a_26580_23588# VGND 0.46161f
C33285 a_26132_23588# VGND 0.47597f
C33286 a_25684_23588# VGND 0.45595f
C33287 a_25236_23588# VGND 0.45589f
C33288 a_24788_23588# VGND 0.45589f
C33289 a_24340_23588# VGND 0.45595f
C33290 a_23892_23588# VGND 0.4559f
C33291 a_23444_23588# VGND 0.45724f
C33292 a_22996_23588# VGND 0.45589f
C33293 a_22548_23588# VGND 0.46795f
C33294 a_21964_23544# VGND 0.28946f
C33295 a_21516_23544# VGND 0.29082f
C33296 a_21068_23544# VGND 0.28898f
C33297 a_20620_23544# VGND 0.29122f
C33298 a_20172_23544# VGND 0.30865f
C33299 a_19724_23544# VGND 0.29648f
C33300 a_19276_23544# VGND 0.2841f
C33301 a_18828_23544# VGND 0.2841f
C33302 a_18380_23544# VGND 0.28575f
C33303 a_17932_23544# VGND 0.28236f
C33304 a_17484_23544# VGND 0.28236f
C33305 a_17036_23544# VGND 0.28236f
C33306 a_16588_23544# VGND 0.28236f
C33307 a_16140_23544# VGND 0.28236f
C33308 a_15692_23544# VGND 0.28236f
C33309 a_15244_23544# VGND 0.28236f
C33310 a_14796_23544# VGND 0.29228f
C33311 a_21876_23588# VGND 0.47083f
C33312 a_21428_23588# VGND 0.45984f
C33313 a_20980_23588# VGND 0.46157f
C33314 a_20532_23588# VGND 0.46423f
C33315 a_20084_23588# VGND 0.49306f
C33316 a_19636_23588# VGND 0.46467f
C33317 a_19188_23588# VGND 0.45666f
C33318 a_18740_23588# VGND 0.45666f
C33319 a_18292_23588# VGND 0.47155f
C33320 a_17844_23588# VGND 0.44029f
C33321 a_17396_23588# VGND 0.44029f
C33322 a_16948_23588# VGND 0.44029f
C33323 a_16500_23588# VGND 0.44029f
C33324 a_16052_23588# VGND 0.44029f
C33325 a_15604_23588# VGND 0.44029f
C33326 a_15156_23588# VGND 0.44029f
C33327 a_14708_23588# VGND 0.46832f
C33328 a_5052_23544# VGND 0.28654f
C33329 a_4604_23544# VGND 0.31699f
C33330 a_4156_23544# VGND 0.29553f
C33331 a_3708_23544# VGND 0.2812f
C33332 a_3260_23544# VGND 0.2812f
C33333 a_2812_23544# VGND 0.2812f
C33334 a_2364_23544# VGND 0.2812f
C33335 a_1916_23544# VGND 0.2812f
C33336 a_1468_23544# VGND 0.2812f
C33337 a_1020_23544# VGND 0.29134f
C33338 a_4964_23588# VGND 0.47812f
C33339 a_4516_23588# VGND 0.5182f
C33340 a_4068_23588# VGND 0.44538f
C33341 a_3620_23588# VGND 0.43828f
C33342 a_3172_23588# VGND 0.43828f
C33343 a_2724_23588# VGND 0.43828f
C33344 a_2276_23588# VGND 0.43828f
C33345 a_1828_23588# VGND 0.43828f
C33346 a_1380_23588# VGND 0.43828f
C33347 a_932_23588# VGND 0.4664f
C33348 a_67684_24776# VGND 0.4787f
C33349 vgaringosc.tapped_ring.c12_inv_array\[5\]_pdkinv_notouch_.I VGND 1.29411f
C33350 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.I VGND 1.01635f
C33351 a_52852_24372# VGND 0.1953f
C33352 a_51332_24372# VGND 0.49726f
C33353 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.I VGND 0.95366f
C33354 a_56148_24776# VGND 0.45197f
C33355 a_55700_24776# VGND 0.44748f
C33356 a_55252_24776# VGND 0.44748f
C33357 a_54804_24776# VGND 0.44364f
C33358 a_54356_24776# VGND 0.44364f
C33359 a_53908_24776# VGND 0.45533f
C33360 a_53460_24776# VGND 0.47535f
C33361 _478_.D VGND 0.60583f
C33362 a_51988_24776# VGND 0.00101f
C33363 a_43819_24372# VGND 0.00269f
C33364 a_43245_24373# VGND 0.00497f
C33365 a_42853_24373# VGND 0.00204f
C33366 _441_.A2 VGND 0.83649f
C33367 a_67772_24679# VGND 0.28259f
C33368 vgaringosc.tapped_ring.c12_inv_array\[3\]_pdkinv_notouch_.ZN VGND 1.05121f
C33369 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.ZN VGND 0.89169f
C33370 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.ZN VGND 1.19353f
C33371 vgaringosc.tapped_ring.c06_inv_array\[2\]_pdkinv_notouch_.ZN VGND 0.85514f
C33372 vgaringosc.tapped_ring.c06_inv_array\[1\]_pdkinv_notouch_.ZN VGND 0.88444f
C33373 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.ZN VGND 1.11889f
C33374 vgaringosc.tapped_ring.c05_inv_array\[2\]_pdkinv_notouch_.ZN VGND 1.07484f
C33375 vgaringosc.tapped_ring.c05_inv_array\[1\]_pdkinv_notouch_.I VGND 0.83916f
C33376 vgaringosc.tapped_ring.c04_inv_array\[2\]_pdkinv_notouch_.ZN VGND 0.9532f
C33377 vgaringosc.tapped_ring.c04_inv_array\[1\]_pdkinv_notouch_.ZN VGND 0.9062f
C33378 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.ZN VGND 1.03192f
C33379 a_56236_24679# VGND 0.26633f
C33380 a_55788_24679# VGND 0.28671f
C33381 a_55340_24679# VGND 0.28584f
C33382 a_54892_24679# VGND 0.2854f
C33383 a_54444_24679# VGND 0.2841f
C33384 a_53996_24679# VGND 0.2841f
C33385 a_53548_24679# VGND 0.28876f
C33386 _427_.B1 VGND 0.9291f
C33387 _428_.Z VGND 0.73227f
C33388 a_50084_24328# VGND 0.96521f
C33389 _448_.Q VGND 4.88055f
C33390 _447_.Q VGND 5.25209f
C33391 a_42161_24776# VGND 0.07065f
C33392 a_40565_24394# VGND 0.00124f
C33393 a_39985_24372# VGND 0.00661f
C33394 a_39781_24372# VGND 0.00757f
C33395 a_39587_24372# VGND 0.00803f
C33396 a_39004_24463# VGND 0.00145f
C33397 a_37424_24463# VGND 0.00176f
C33398 a_36496_24463# VGND 0.00166f
C33399 hold1.Z VGND 1.09934f
C33400 _260_.ZN VGND 1.22618f
C33401 a_41476_24776# VGND 0.49235f
C33402 a_40357_24776# VGND 0.04787f
C33403 _441_.A3 VGND 1.0857f
C33404 a_41564_24679# VGND 0.29288f
C33405 _432_.ZN VGND 0.98721f
C33406 _433_.ZN VGND 0.83136f
C33407 _435_.ZN VGND 0.91783f
C33408 _452_.Q VGND 5.73425f
C33409 _430_.ZN VGND 0.93541f
C33410 a_38616_24328# VGND 0.56353f
C33411 a_32048_24463# VGND 0.0017f
C33412 a_31120_24463# VGND 0.00146f
C33413 a_37472_24419# VGND 0.84732f
C33414 a_37179_24831# VGND 0.45207f
C33415 a_36172_24463# VGND 0.30204f
C33416 a_36544_24419# VGND 0.43007f
C33417 a_35616_24776# VGND 1.51537f
C33418 a_34756_24776# VGND 0.47264f
C33419 a_34308_24776# VGND 0.49024f
C33420 a_33524_24776# VGND 0.47414f
C33421 a_33076_24776# VGND 0.48128f
C33422 a_29163_24394# VGND 0.00126f
C33423 a_27552_24397# VGND 0.00424f
C33424 a_34844_24679# VGND 0.24844f
C33425 a_34396_24679# VGND 0.28927f
C33426 a_33612_24679# VGND 0.27074f
C33427 a_33164_24679# VGND 0.29036f
C33428 a_32096_24419# VGND 0.8482f
C33429 a_31803_24831# VGND 0.44973f
C33430 a_30796_24463# VGND 0.29387f
C33431 a_31168_24419# VGND 0.42413f
C33432 a_30240_24776# VGND 1.46951f
C33433 a_28903_24776# VGND 0.0596f
C33434 a_28679_24776# VGND 0.00109f
C33435 a_26548_24372# VGND 0.7352f
C33436 a_27924_24776# VGND 0.48208f
C33437 a_25796_24776# VGND 0.47128f
C33438 a_25348_24776# VGND 0.45666f
C33439 a_24900_24776# VGND 0.45666f
C33440 a_24452_24776# VGND 0.45666f
C33441 a_24004_24776# VGND 0.45666f
C33442 a_23556_24776# VGND 0.45666f
C33443 a_23108_24776# VGND 0.45666f
C33444 a_22660_24776# VGND 0.45666f
C33445 a_22212_24776# VGND 0.47155f
C33446 a_21764_24776# VGND 0.45927f
C33447 a_21316_24776# VGND 0.46144f
C33448 a_20868_24776# VGND 0.46336f
C33449 a_20420_24776# VGND 0.4663f
C33450 a_19972_24776# VGND 0.50071f
C33451 a_19524_24776# VGND 0.46161f
C33452 a_19076_24776# VGND 0.4579f
C33453 a_18628_24776# VGND 0.4724f
C33454 a_17844_24776# VGND 0.44215f
C33455 a_17396_24776# VGND 0.43828f
C33456 a_16948_24776# VGND 0.43828f
C33457 a_16500_24776# VGND 0.43828f
C33458 a_16052_24776# VGND 0.43828f
C33459 a_15604_24776# VGND 0.43828f
C33460 a_15156_24776# VGND 0.43828f
C33461 a_14708_24776# VGND 0.4664f
C33462 a_5300_24776# VGND 0.48995f
C33463 a_4852_24776# VGND 0.48956f
C33464 a_4068_24776# VGND 0.44997f
C33465 a_3620_24776# VGND 0.43828f
C33466 a_3172_24776# VGND 0.43828f
C33467 a_2724_24776# VGND 0.43828f
C33468 a_2276_24776# VGND 0.43828f
C33469 a_1828_24776# VGND 0.43828f
C33470 a_1380_24776# VGND 0.43828f
C33471 a_932_24776# VGND 0.4664f
C33472 a_28012_24679# VGND 0.26144f
C33473 a_27172_24328# VGND 0.69622f
C33474 a_25884_24679# VGND 0.28953f
C33475 a_25436_24679# VGND 0.28584f
C33476 a_24988_24679# VGND 0.28236f
C33477 a_24540_24679# VGND 0.28458f
C33478 a_24092_24679# VGND 0.28262f
C33479 a_23644_24679# VGND 0.28581f
C33480 a_23196_24679# VGND 0.28582f
C33481 a_22748_24679# VGND 0.28575f
C33482 a_22300_24679# VGND 0.28652f
C33483 a_21852_24679# VGND 0.28537f
C33484 a_21404_24679# VGND 0.28816f
C33485 a_20956_24679# VGND 0.28996f
C33486 a_20508_24679# VGND 0.29249f
C33487 a_20060_24679# VGND 0.32519f
C33488 a_19612_24679# VGND 0.29254f
C33489 a_19164_24679# VGND 0.28426f
C33490 a_18716_24679# VGND 0.28799f
C33491 a_17932_24679# VGND 0.26958f
C33492 a_17484_24679# VGND 0.2812f
C33493 a_17036_24679# VGND 0.2812f
C33494 a_16588_24679# VGND 0.2812f
C33495 a_16140_24679# VGND 0.2812f
C33496 a_15692_24679# VGND 0.2812f
C33497 a_15244_24679# VGND 0.2812f
C33498 a_14796_24679# VGND 0.29134f
C33499 a_5388_24679# VGND 0.3139f
C33500 a_4940_24679# VGND 0.29949f
C33501 a_4156_24679# VGND 0.28278f
C33502 a_3708_24679# VGND 0.2812f
C33503 a_3260_24679# VGND 0.2812f
C33504 a_2812_24679# VGND 0.2812f
C33505 a_2364_24679# VGND 0.2812f
C33506 a_1916_24679# VGND 0.2812f
C33507 a_1468_24679# VGND 0.2812f
C33508 a_1020_24679# VGND 0.29134f
C33509 a_59226_25156# VGND 0.00252f
C33510 vgaringosc.tapped_ring.c12_inv_array\[1\]_pdkinv_notouch_.I VGND 0.89534f
C33511 a_62796_25640# VGND 0.00951f
C33512 a_62404_25640# VGND 0.00198f
C33513 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.ZN VGND 0.98635f
C33514 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.I VGND 1.04602f
C33515 vgaringosc.tapped_ring.c11_inv_array\[14\]_pdkinv_notouch_.ZN VGND 0.90895f
C33516 vgaringosc.tapped_ring.c07_inv_array\[1\]_pdkinv_notouch_.ZN VGND 0.87216f
C33517 vgaringosc.tapped_ring.c07_inv_array\[0\]_pdkinv_notouch_.I VGND 1.51596f
C33518 a_62560_25112# VGND 0.45621f
C33519 a_61836_25515# VGND 1.03321f
C33520 a_60524_25640# VGND 0.00205f
C33521 a_60084_25640# VGND 0.01024f
C33522 a_60212_25156# VGND 1.0362f
C33523 vgaringosc.tapped_ring.c06_inv_array\[0\]_pdkinv_notouch_.I VGND 1.28909f
C33524 a_59652_25640# VGND 0.46338f
C33525 vgaringosc.tapped_ring.c04_inv_array\[3\]_pdkinv_notouch_.ZN VGND 1.37942f
C33526 vgaringosc.tapped_ring.c12_inv_array\[31\]_pdkinv_notouch_.ZN VGND 1.58651f
C33527 a_58364_25112# VGND 0.2742f
C33528 a_57916_25112# VGND 0.28647f
C33529 a_55788_25112# VGND 0.26105f
C33530 a_55340_25112# VGND 0.28627f
C33531 a_54892_25112# VGND 0.2841f
C33532 a_54444_25112# VGND 0.2841f
C33533 a_53996_25112# VGND 0.28756f
C33534 a_44028_25156# VGND 0.00127f
C33535 clkbuf_1_0__f_clk.I VGND 8.93737f
C33536 a_58276_25156# VGND 0.48636f
C33537 a_57828_25156# VGND 0.46277f
C33538 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.ZN VGND 0.86744f
C33539 a_55700_25156# VGND 0.4851f
C33540 a_55252_25156# VGND 0.45642f
C33541 a_54804_25156# VGND 0.46001f
C33542 a_54356_25156# VGND 0.46764f
C33543 a_53908_25156# VGND 0.48967f
C33544 _474_.Q VGND 4.45669f
C33545 _279_.Z VGND 1.46768f
C33546 a_47297_25596# VGND 0.54363f
C33547 _281_.ZN VGND 2.03127f
C33548 a_46156_25112# VGND 0.2727f
C33549 a_46068_25156# VGND 0.4918f
C33550 a_40468_25157# VGND 0.00492f
C33551 a_43600_25640# VGND 0.00514f
C33552 a_43192_25640# VGND 0.00295f
C33553 a_42784_25640# VGND 0.00242f
C33554 a_42376_25640# VGND 0.00534f
C33555 _260_.A2 VGND 1.30615f
C33556 hold2.I VGND 2.71832f
C33557 _264_.B VGND 1.01527f
C33558 a_40676_25640# VGND 0.00256f
C33559 _444_.D VGND 1.05961f
C33560 _260_.A1 VGND 2.55262f
C33561 _261_.ZN VGND 0.63421f
C33562 _441_.ZN VGND 0.5778f
C33563 _436_.ZN VGND 1.04772f
C33564 _311_.A2 VGND 2.88804f
C33565 a_37532_25112# VGND 0.27527f
C33566 a_37084_25112# VGND 0.28907f
C33567 a_36636_25112# VGND 0.28832f
C33568 a_36188_25112# VGND 0.29471f
C33569 a_35740_25112# VGND 0.30771f
C33570 a_34400_25641# VGND 0.0017f
C33571 a_33472_25641# VGND 0.00146f
C33572 a_37444_25156# VGND 0.45603f
C33573 a_36996_25156# VGND 0.44657f
C33574 a_36548_25156# VGND 0.44815f
C33575 a_36100_25156# VGND 0.45026f
C33576 a_35652_25156# VGND 0.48459f
C33577 a_34155_25273# VGND 0.4677f
C33578 a_34448_25597# VGND 1.11865f
C33579 a_33148_25641# VGND 0.30019f
C33580 a_33520_25597# VGND 0.4167f
C33581 a_32592_25227# VGND 1.47833f
C33582 a_31820_25112# VGND 0.24504f
C33583 _459_.D VGND 0.6646f
C33584 a_31732_25156# VGND 0.47942f
C33585 a_30476_25112# VGND 0.24405f
C33586 a_30388_25156# VGND 0.49531f
C33587 a_29136_25641# VGND 0.00185f
C33588 a_28208_25641# VGND 0.00172f
C33589 a_28891_25273# VGND 0.45876f
C33590 a_29184_25597# VGND 0.83805f
C33591 a_27884_25641# VGND 0.32298f
C33592 a_28256_25597# VGND 0.42956f
C33593 _355_.ZN VGND 1.39551f
C33594 a_27328_25227# VGND 1.49879f
C33595 a_25888_25641# VGND 0.0017f
C33596 a_24960_25641# VGND 0.00146f
C33597 a_25643_25273# VGND 0.4662f
C33598 a_25936_25597# VGND 0.8387f
C33599 a_24636_25641# VGND 0.29991f
C33600 a_25008_25597# VGND 0.42419f
C33601 a_24080_25227# VGND 1.47742f
C33602 a_23084_25112# VGND 0.25499f
C33603 a_22636_25112# VGND 0.29059f
C33604 a_22996_25156# VGND 0.47473f
C33605 a_22548_25156# VGND 0.47421f
C33606 a_21964_25112# VGND 0.28946f
C33607 a_21516_25112# VGND 0.29082f
C33608 a_21068_25112# VGND 0.28898f
C33609 a_20620_25112# VGND 0.29122f
C33610 a_20172_25112# VGND 0.30865f
C33611 a_19724_25112# VGND 0.29648f
C33612 a_19276_25112# VGND 0.2841f
C33613 a_18828_25112# VGND 0.2841f
C33614 a_18380_25112# VGND 0.28575f
C33615 a_17932_25112# VGND 0.28236f
C33616 a_17484_25112# VGND 0.28236f
C33617 a_17036_25112# VGND 0.28236f
C33618 a_16588_25112# VGND 0.28236f
C33619 a_16140_25112# VGND 0.28236f
C33620 a_15692_25112# VGND 0.28236f
C33621 a_15244_25112# VGND 0.28236f
C33622 a_14796_25112# VGND 0.29228f
C33623 a_21876_25156# VGND 0.47732f
C33624 a_21428_25156# VGND 0.47309f
C33625 a_20980_25156# VGND 0.47611f
C33626 a_20532_25156# VGND 0.47491f
C33627 a_20084_25156# VGND 0.50137f
C33628 a_19636_25156# VGND 0.46606f
C33629 a_19188_25156# VGND 0.45666f
C33630 a_18740_25156# VGND 0.45666f
C33631 a_18292_25156# VGND 0.47156f
C33632 a_17844_25156# VGND 0.44029f
C33633 a_17396_25156# VGND 0.44029f
C33634 a_16948_25156# VGND 0.44029f
C33635 a_16500_25156# VGND 0.44029f
C33636 a_16052_25156# VGND 0.44029f
C33637 a_15604_25156# VGND 0.44029f
C33638 a_15156_25156# VGND 0.44029f
C33639 a_14708_25156# VGND 0.46832f
C33640 a_5052_25112# VGND 0.28654f
C33641 a_4604_25112# VGND 0.31699f
C33642 a_4156_25112# VGND 0.29553f
C33643 a_3708_25112# VGND 0.2812f
C33644 a_3260_25112# VGND 0.2812f
C33645 a_2812_25112# VGND 0.2812f
C33646 a_2364_25112# VGND 0.2812f
C33647 a_1916_25112# VGND 0.2812f
C33648 a_1468_25112# VGND 0.2812f
C33649 a_1020_25112# VGND 0.29134f
C33650 a_4964_25156# VGND 0.47812f
C33651 a_4516_25156# VGND 0.5182f
C33652 a_4068_25156# VGND 0.44538f
C33653 a_3620_25156# VGND 0.43828f
C33654 a_3172_25156# VGND 0.43828f
C33655 a_2724_25156# VGND 0.43828f
C33656 a_2276_25156# VGND 0.43828f
C33657 a_1828_25156# VGND 0.43828f
C33658 a_1380_25156# VGND 0.43828f
C33659 a_932_25156# VGND 0.4664f
C33660 vgaringosc.tapped_ring.c11_inv_array\[10\]_pdkinv_notouch_.I VGND 1.00566f
C33661 vgaringosc.tapped_ring.c11_inv_array\[13\]_pdkinv_notouch_.I VGND 1.25491f
C33662 a_65668_26344# VGND 0.48254f
C33663 a_59605_25962# VGND 0.00133f
C33664 a_56828_25940# VGND 0.00198f
C33665 a_56388_25940# VGND 0.00951f
C33666 a_64772_26344# VGND 0.49462f
C33667 _245_.I1 VGND 1.43053f
C33668 a_62308_26344# VGND 0.46264f
C33669 a_61860_26344# VGND 0.45838f
C33670 a_61412_26344# VGND 0.47582f
C33671 a_60964_26344# VGND 0.46236f
C33672 a_60516_26344# VGND 0.47761f
C33673 a_59397_26344# VGND 0.05f
C33674 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.ZN VGND 0.99608f
C33675 vgaringosc.tapped_ring.c11_inv_array\[11\]_pdkinv_notouch_.ZN VGND 1.30397f
C33676 a_65756_26247# VGND 0.26433f
C33677 a_64860_26247# VGND 0.27132f
C33678 vgaringosc.tapped_ring.c08_inv_array\[1\]_pdkinv_notouch_.ZN VGND 0.82627f
C33679 vgaringosc.tapped_ring.c08_inv_array\[0\]_pdkinv_notouch_.ZN VGND 0.90729f
C33680 vgaringosc.tapped_ring.c07_inv_array\[2\]_pdkinv_notouch_.ZN VGND 0.99056f
C33681 a_62396_26247# VGND 0.26331f
C33682 a_61948_26247# VGND 0.28801f
C33683 a_61500_26247# VGND 0.28749f
C33684 a_61052_26247# VGND 0.28721f
C33685 a_60604_26247# VGND 0.28979f
C33686 _251_.ZN VGND 0.68763f
C33687 _231_.ZN VGND 0.94998f
C33688 a_58948_26344# VGND 0.50521f
C33689 a_58500_26344# VGND 0.49462f
C33690 a_53280_26031# VGND 0.00146f
C33691 a_52352_26031# VGND 0.00186f
C33692 a_51016_25940# VGND 0.00558f
C33693 a_54692_26344# VGND 0.4801f
C33694 _412_.ZN VGND 0.61728f
C33695 a_59036_26247# VGND 0.29921f
C33696 a_58588_26247# VGND 0.30308f
C33697 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.ZN VGND 0.9754f
C33698 a_56516_26344# VGND 1.03014f
C33699 vgaringosc.tapped_ring.c04_inv_array\[0\]_pdkinv_notouch_.I VGND 1.29111f
C33700 a_55956_25940# VGND 0.46778f
C33701 vgaringosc.tapped_ring.c03_inv_array\[0\]_pdkinv_notouch_.I VGND 1.62404f
C33702 a_54780_26247# VGND 0.26126f
C33703 a_52744_26031# VGND 0.42052f
C33704 a_52848_25987# VGND 0.29992f
C33705 a_52360_26355# VGND 1.47831f
C33706 a_51956_26183# VGND 0.4648f
C33707 _412_.B2 VGND 0.87047f
C33708 a_50792_26344# VGND 0.01028f
C33709 a_47636_25940# VGND 2.08997f
C33710 a_47291_25940# VGND 0.00253f
C33711 a_45664_26031# VGND 0.00146f
C33712 a_44736_26031# VGND 0.00173f
C33713 _284_.B VGND 1.62769f
C33714 a_43253_25940# VGND 0.00299f
C33715 a_42587_25940# VGND 0.00251f
C33716 _402_.ZN VGND 0.87462f
C33717 a_51576_25896# VGND 0.84528f
C33718 a_50120_26476# VGND 0.73977f
C33719 _381_.A2 VGND 1.81582f
C33720 _282_.ZN VGND 0.77192f
C33721 _421_.A1 VGND 1.60754f
C33722 a_45128_26031# VGND 0.41758f
C33723 a_45232_25987# VGND 0.29654f
C33724 a_44744_26355# VGND 1.47494f
C33725 a_44340_26183# VGND 0.45756f
C33726 _435_.A3 VGND 1.36424f
C33727 a_34516_25940# VGND 0.00262f
C33728 a_33188_25940# VGND 0.15067f
C33729 a_43736_25896# VGND 1.1145f
C33730 _451_.Q VGND 4.07074f
C33731 hold2.Z VGND 0.65666f
C33732 a_41476_26344# VGND 0.47312f
C33733 a_41028_26344# VGND 0.47704f
C33734 a_40580_26344# VGND 0.45426f
C33735 a_40132_26344# VGND 0.46667f
C33736 a_39684_26344# VGND 0.46454f
C33737 a_39236_26344# VGND 0.48683f
C33738 _431_.A3 VGND 0.97569f
C33739 a_37892_26344# VGND 0.48694f
C33740 a_37444_26344# VGND 0.44753f
C33741 a_36996_26344# VGND 0.4506f
C33742 a_36548_26344# VGND 0.44845f
C33743 a_36100_26344# VGND 0.45106f
C33744 a_35652_26344# VGND 0.4763f
C33745 a_35204_26344# VGND 0.47026f
C33746 a_34308_26344# VGND 0.00492f
C33747 a_41564_26247# VGND 0.29371f
C33748 a_41116_26247# VGND 0.28593f
C33749 a_40668_26247# VGND 0.2854f
C33750 a_40220_26247# VGND 0.28669f
C33751 a_39772_26247# VGND 0.28425f
C33752 a_39324_26247# VGND 0.28887f
C33753 _438_.A2 VGND 1.85892f
C33754 a_37980_26247# VGND 0.26457f
C33755 a_37532_26247# VGND 0.28671f
C33756 a_37084_26247# VGND 0.28902f
C33757 a_36636_26247# VGND 0.2902f
C33758 a_36188_26247# VGND 0.29112f
C33759 a_35740_26247# VGND 0.30757f
C33760 a_35292_26247# VGND 0.29679f
C33761 _460_.D VGND 0.47832f
C33762 a_32292_26344# VGND 0.4752f
C33763 a_31844_26344# VGND 0.47084f
C33764 a_30036_25940# VGND 0.00255f
C33765 a_29348_25940# VGND 0.00366f
C33766 a_29164_25940# VGND 0.00353f
C33767 a_28756_25940# VGND 0.00638f
C33768 a_28552_25940# VGND 0.00899f
C33769 _358_.A2 VGND 0.79953f
C33770 a_29828_26344# VGND 0.00492f
C33771 _359_.ZN VGND 0.90351f
C33772 _360_.ZN VGND 0.47061f
C33773 a_32380_26247# VGND 0.28741f
C33774 a_31932_26247# VGND 0.28941f
C33775 a_30724_26020# VGND 1.12817f
C33776 a_27588_26344# VGND 0.49242f
C33777 a_27140_26344# VGND 0.47448f
C33778 _457_.D VGND 0.68772f
C33779 a_22304_26031# VGND 0.0017f
C33780 a_21376_26031# VGND 0.00161f
C33781 a_24228_26344# VGND 0.47743f
C33782 a_23780_26344# VGND 0.47408f
C33783 a_23332_26344# VGND 0.48632f
C33784 a_27676_26247# VGND 0.29894f
C33785 a_27228_26247# VGND 0.28787f
C33786 _352_.ZN VGND 0.46061f
C33787 a_24316_26247# VGND 0.25545f
C33788 a_23868_26247# VGND 0.289f
C33789 a_23420_26247# VGND 0.28834f
C33790 a_22352_25987# VGND 0.84262f
C33791 a_22059_26399# VGND 0.45111f
C33792 a_21052_26031# VGND 0.3071f
C33793 a_21424_25987# VGND 0.4253f
C33794 a_20496_26344# VGND 1.48198f
C33795 a_19524_26344# VGND 0.47598f
C33796 a_19076_26344# VGND 0.46508f
C33797 a_18628_26344# VGND 0.47931f
C33798 a_17844_26344# VGND 0.44215f
C33799 a_17396_26344# VGND 0.43828f
C33800 a_16948_26344# VGND 0.43828f
C33801 a_16500_26344# VGND 0.43828f
C33802 a_16052_26344# VGND 0.43828f
C33803 a_15604_26344# VGND 0.43828f
C33804 a_15156_26344# VGND 0.43828f
C33805 a_14708_26344# VGND 0.4664f
C33806 a_5300_26344# VGND 0.48995f
C33807 a_4852_26344# VGND 0.48956f
C33808 a_4068_26344# VGND 0.44997f
C33809 a_3620_26344# VGND 0.43828f
C33810 a_3172_26344# VGND 0.43828f
C33811 a_2724_26344# VGND 0.43828f
C33812 a_2276_26344# VGND 0.43828f
C33813 a_1828_26344# VGND 0.43828f
C33814 a_1380_26344# VGND 0.43828f
C33815 a_932_26344# VGND 0.4664f
C33816 a_19612_26247# VGND 0.26455f
C33817 a_19164_26247# VGND 0.28671f
C33818 a_18716_26247# VGND 0.29263f
C33819 a_17932_26247# VGND 0.26996f
C33820 a_17484_26247# VGND 0.2812f
C33821 a_17036_26247# VGND 0.28121f
C33822 a_16588_26247# VGND 0.28136f
C33823 a_16140_26247# VGND 0.28133f
C33824 a_15692_26247# VGND 0.28431f
C33825 a_15244_26247# VGND 0.2812f
C33826 a_14796_26247# VGND 0.29134f
C33827 a_5388_26247# VGND 0.3139f
C33828 a_4940_26247# VGND 0.29949f
C33829 a_4156_26247# VGND 0.28278f
C33830 a_3708_26247# VGND 0.2812f
C33831 a_3260_26247# VGND 0.2812f
C33832 a_2812_26247# VGND 0.2812f
C33833 a_2364_26247# VGND 0.2812f
C33834 a_1916_26247# VGND 0.2812f
C33835 a_1468_26247# VGND 0.2812f
C33836 a_1020_26247# VGND 0.29134f
C33837 vgaringosc.tapped_ring.c11_inv_array\[8\]_pdkinv_notouch_.I VGND 0.9931f
C33838 a_64972_26680# VGND 0.26485f
C33839 a_63180_26680# VGND 0.26435f
C33840 a_62732_26680# VGND 0.2879f
C33841 a_62284_26680# VGND 0.28601f
C33842 a_61836_26680# VGND 0.28974f
C33843 a_51968_26724# VGND 0.00181f
C33844 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.ZN VGND 1.18388f
C33845 vgaringosc.tapped_ring.c11_inv_array\[6\]_pdkinv_notouch_.ZN VGND 0.97149f
C33846 a_64884_26724# VGND 0.47885f
C33847 vgaringosc.tapped_ring.c08_inv_array\[3\]_pdkinv_notouch_.ZN VGND 0.85963f
C33848 vgaringosc.tapped_ring.c08_inv_array\[2\]_pdkinv_notouch_.ZN VGND 0.83876f
C33849 a_63092_26724# VGND 0.47498f
C33850 a_62644_26724# VGND 0.4619f
C33851 a_62196_26724# VGND 0.46251f
C33852 a_61748_26724# VGND 0.48014f
C33853 a_60828_26680# VGND 0.27099f
C33854 a_59620_27208# VGND 0.48742f
C33855 a_59260_26680# VGND 0.24959f
C33856 a_58140_26680# VGND 0.25414f
C33857 a_57276_27208# VGND 0.00198f
C33858 a_56836_27208# VGND 0.00951f
C33859 a_55340_26680# VGND 0.26213f
C33860 a_54892_26680# VGND 0.28584f
C33861 a_54444_26680# VGND 0.28591f
C33862 a_53996_26680# VGND 0.28809f
C33863 a_60740_26724# VGND 0.49657f
C33864 _244_.Z VGND 0.7065f
C33865 _245_.Z VGND 0.73249f
C33866 a_59172_26724# VGND 0.47213f
C33867 a_58052_26724# VGND 0.47296f
C33868 a_56964_26724# VGND 1.04816f
C33869 vgaringosc.tapped_ring.c02_inv_array\[0\]_pdkinv_notouch_.I VGND 1.27285f
C33870 a_56404_27208# VGND 0.45784f
C33871 a_55252_26724# VGND 0.46253f
C33872 a_54804_26724# VGND 0.46253f
C33873 a_54356_26724# VGND 0.45954f
C33874 a_53908_26724# VGND 0.49271f
C33875 a_52988_26680# VGND 0.26731f
C33876 a_51436_27208# VGND 0.00146f
C33877 _398_.C VGND 3.14011f
C33878 _384_.A3 VGND 3.65821f
C33879 a_52900_26724# VGND 0.49305f
C33880 _284_.A2 VGND 2.12477f
C33881 a_51048_26680# VGND 0.60576f
C33882 _395_.A2 VGND 1.30596f
C33883 clkload0.Z VGND 0.3795f
C33884 a_48384_26724# VGND 1.44512f
C33885 a_43440_26841# VGND 0.00127f
C33886 a_49764_26724# VGND 0.96524f
C33887 _419_.A4 VGND 1.50434f
C33888 _412_.A1 VGND 1.45794f
C33889 a_47173_27208# VGND 0.00266f
C33890 _424_.A2 VGND 3.91571f
C33891 a_46198_27060# VGND 0.73309f
C33892 a_44816_27209# VGND 0.00176f
C33893 a_43888_27209# VGND 0.00158f
C33894 a_43396_27209# VGND 0.00107f
C33895 a_44571_26841# VGND 0.45813f
C33896 a_44864_27165# VGND 0.83966f
C33897 a_43564_27209# VGND 0.31287f
C33898 a_43936_27165# VGND 0.42606f
C33899 a_43008_26795# VGND 1.5142f
C33900 a_41344_27209# VGND 0.0017f
C33901 a_40416_27209# VGND 0.00146f
C33902 a_41099_26841# VGND 0.46302f
C33903 a_41392_27165# VGND 0.85219f
C33904 a_40092_27209# VGND 0.29442f
C33905 a_40464_27165# VGND 0.42356f
C33906 _442_.ZN VGND 0.76832f
C33907 a_39536_26795# VGND 1.47437f
C33908 a_37532_26680# VGND 0.2721f
C33909 a_37084_26680# VGND 0.28687f
C33910 a_36636_26680# VGND 0.28821f
C33911 a_36188_26680# VGND 0.29066f
C33912 a_32628_26725# VGND 0.00492f
C33913 a_35756_27216# VGND 0.00176f
C33914 a_37444_26724# VGND 0.48026f
C33915 a_36996_26724# VGND 0.47371f
C33916 a_36548_26724# VGND 0.47142f
C33917 a_36100_26724# VGND 0.48926f
C33918 a_35140_26680# VGND 1.19604f
C33919 a_34532_27208# VGND 0.00861f
C33920 a_34348_27208# VGND 0.00586f
C33921 a_33940_27208# VGND 0.00324f
C33922 a_33764_27208# VGND 0.00344f
C33923 a_32836_27208# VGND 0.00258f
C33924 a_28596_26725# VGND 0.00792f
C33925 _358_.A3 VGND 2.47381f
C33926 a_31484_26680# VGND 0.26348f
C33927 a_31031_27208# VGND 0.00761f
C33928 a_30847_27208# VGND 0.00657f
C33929 a_31396_26724# VGND 0.48362f
C33930 _336_.Z VGND 1.70639f
C33931 _355_.B VGND 0.67633f
C33932 a_28804_27208# VGND 0.00271f
C33933 a_28124_26680# VGND 0.26619f
C33934 a_27676_26680# VGND 0.32172f
C33935 a_27228_26680# VGND 0.28753f
C33936 a_26112_27209# VGND 0.0017f
C33937 a_25184_27209# VGND 0.00146f
C33938 _336_.A1 VGND 1.73966f
C33939 _336_.A2 VGND 3.25378f
C33940 a_28036_26724# VGND 0.48447f
C33941 a_27588_26724# VGND 0.48931f
C33942 a_27140_26724# VGND 0.48406f
C33943 a_25867_26841# VGND 0.46827f
C33944 a_26160_27165# VGND 0.84765f
C33945 a_24860_27209# VGND 0.29963f
C33946 a_25232_27165# VGND 0.41967f
C33947 _351_.ZN VGND 0.67668f
C33948 a_24304_26795# VGND 1.47881f
C33949 a_21600_26725# VGND 0.00624f
C33950 a_21868_27208# VGND 0.00259f
C33951 _455_.D VGND 0.73383f
C33952 a_20844_26680# VGND 0.25945f
C33953 a_20396_26680# VGND 0.2954f
C33954 a_19948_26680# VGND 0.33481f
C33955 a_18048_27209# VGND 0.00146f
C33956 a_17120_27209# VGND 0.00146f
C33957 a_16796_27209# VGND 0.29374f
C33958 a_17168_27165# VGND 0.41897f
C33959 a_16240_26795# VGND 1.47004f
C33960 a_20756_26724# VGND 0.47129f
C33961 a_20308_26724# VGND 0.45646f
C33962 a_19860_26724# VGND 0.48275f
C33963 a_18096_27165# VGND 1.69111f
C33964 a_17803_26841# VGND 0.67416f
C33965 a_15244_26680# VGND 0.25309f
C33966 a_14796_26680# VGND 0.29512f
C33967 a_15156_26724# VGND 0.45148f
C33968 a_14708_26724# VGND 0.47523f
C33969 a_5052_26680# VGND 0.28654f
C33970 a_4604_26680# VGND 0.31699f
C33971 a_4156_26680# VGND 0.29553f
C33972 a_3708_26680# VGND 0.2812f
C33973 a_3260_26680# VGND 0.2812f
C33974 a_2812_26680# VGND 0.2812f
C33975 a_2364_26680# VGND 0.2812f
C33976 a_1916_26680# VGND 0.2812f
C33977 a_1468_26680# VGND 0.2812f
C33978 a_1020_26680# VGND 0.29134f
C33979 a_4964_26724# VGND 0.47812f
C33980 a_4516_26724# VGND 0.5182f
C33981 a_4068_26724# VGND 0.44538f
C33982 a_3620_26724# VGND 0.43828f
C33983 a_3172_26724# VGND 0.43828f
C33984 a_2724_26724# VGND 0.43828f
C33985 a_2276_26724# VGND 0.43828f
C33986 a_1828_26724# VGND 0.43828f
C33987 a_1380_26724# VGND 0.43828f
C33988 a_932_26724# VGND 0.4664f
C33989 vgaringosc.tapped_ring.c11_inv_array\[5\]_pdkinv_notouch_.I VGND 1.18005f
C33990 a_65668_27912# VGND 0.4818f
C33991 a_59380_27508# VGND 0.00278f
C33992 a_58020_27508# VGND 0.51709f
C33993 a_51883_27508# VGND 0.00261f
C33994 a_51317_27508# VGND 0.00359f
C33995 a_50068_27508# VGND 0.52017f
C33996 a_64100_27912# VGND 0.47455f
C33997 a_62756_27912# VGND 0.4697f
C33998 a_62308_27912# VGND 0.46384f
C33999 a_61860_27912# VGND 0.46384f
C34000 a_61412_27912# VGND 0.4749f
C34001 a_60964_27912# VGND 0.47287f
C34002 a_60516_27912# VGND 0.47608f
C34003 a_60068_27912# VGND 0.46867f
C34004 a_59172_27912# VGND 0.01245f
C34005 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.ZN VGND 0.97214f
C34006 a_65756_27815# VGND 0.26179f
C34007 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.I VGND 1.10948f
C34008 a_64188_27815# VGND 0.26036f
C34009 vgaringosc.tapped_ring.c08_inv_array\[4\]_pdkinv_notouch_.ZN VGND 1.0444f
C34010 a_62844_27815# VGND 0.2626f
C34011 a_62396_27815# VGND 0.28909f
C34012 a_61948_27815# VGND 0.29011f
C34013 a_61500_27815# VGND 0.29175f
C34014 a_61052_27815# VGND 0.28747f
C34015 a_60604_27815# VGND 0.28852f
C34016 a_60156_27815# VGND 0.29069f
C34017 _247_.B VGND 0.57374f
C34018 _243_.ZN VGND 0.70309f
C34019 a_49172_27508# VGND 0.0035f
C34020 a_48988_27508# VGND 0.00329f
C34021 a_48580_27508# VGND 0.00589f
C34022 a_48376_27508# VGND 0.00863f
C34023 a_57156_27912# VGND 0.46633f
C34024 vgaringosc.tapped_ring.c01_inv_array\[1\]_pdkinv_notouch_.I VGND 1.0807f
C34025 a_56036_27912# VGND 0.46971f
C34026 a_55588_27912# VGND 0.47699f
C34027 a_55140_27912# VGND 0.4699f
C34028 a_53572_27912# VGND 0.47621f
C34029 a_53124_27912# VGND 0.47287f
C34030 a_52676_27912# VGND 0.47757f
C34031 a_52228_27912# VGND 0.47835f
C34032 _243_.B2 VGND 0.59195f
C34033 _242_.Z VGND 0.64079f
C34034 _241_.Z VGND 0.66737f
C34035 a_57244_27815# VGND 0.2936f
C34036 a_56124_27815# VGND 0.26154f
C34037 a_55676_27815# VGND 0.28671f
C34038 a_55228_27815# VGND 0.28645f
C34039 a_53660_27815# VGND 0.26885f
C34040 a_53212_27815# VGND 0.28824f
C34041 a_52764_27815# VGND 0.28704f
C34042 a_52316_27815# VGND 0.2925f
C34043 _407_.ZN VGND 0.46747f
C34044 a_46171_27508# VGND 0.00262f
C34045 a_45577_27509# VGND 0.00383f
C34046 a_45169_27509# VGND 0.006f
C34047 a_38768_27599# VGND 0.0017f
C34048 a_37840_27599# VGND 0.00146f
C34049 _411_.A2 VGND 2.85669f
C34050 _408_.ZN VGND 0.56597f
C34051 _424_.B1 VGND 4.21237f
C34052 _397_.A4 VGND 1.67303f
C34053 _470_.D VGND 0.57436f
C34054 a_44961_27912# VGND 0.02773f
C34055 _400_.ZN VGND 0.73817f
C34056 _403_.ZN VGND 0.5591f
C34057 _330_.A1 VGND 6.80689f
C34058 a_44388_27912# VGND 0.4751f
C34059 a_43940_27912# VGND 0.48295f
C34060 a_43492_27912# VGND 0.49991f
C34061 a_43044_27912# VGND 0.48115f
C34062 a_42596_27912# VGND 0.46839f
C34063 a_42148_27912# VGND 0.4928f
C34064 a_41140_27912# VGND 0.47266f
C34065 a_40692_27912# VGND 0.47976f
C34066 a_39796_27912# VGND 0.48078f
C34067 a_35660_27508# VGND 0.74537f
C34068 a_35216_27533# VGND 0.00403f
C34069 a_44476_27815# VGND 0.25626f
C34070 a_44028_27815# VGND 0.29545f
C34071 a_43580_27815# VGND 0.29772f
C34072 a_43132_27815# VGND 0.3114f
C34073 a_42684_27815# VGND 0.28429f
C34074 a_42236_27815# VGND 0.28784f
C34075 a_41228_27815# VGND 0.26863f
C34076 a_40780_27815# VGND 0.28981f
C34077 _436_.B VGND 1.15607f
C34078 a_39884_27815# VGND 0.28717f
C34079 a_38816_27555# VGND 0.83943f
C34080 a_38523_27967# VGND 0.46542f
C34081 a_37516_27599# VGND 0.30314f
C34082 a_37888_27555# VGND 0.42459f
C34083 _443_.D VGND 0.66509f
C34084 a_36960_27912# VGND 1.4786f
C34085 _452_.CLK VGND 11.49706f
C34086 a_35874_27937# VGND 0.00103f
C34087 a_30912_27508# VGND 0.00458f
C34088 a_30520_27508# VGND 0.00233f
C34089 a_30128_27508# VGND 0.00412f
C34090 a_29736_27508# VGND 0.00476f
C34091 a_25108_27508# VGND 0.00255f
C34092 a_23872_27599# VGND 0.0017f
C34093 a_22944_27599# VGND 0.00146f
C34094 a_28112_27912# VGND 0.00226f
C34095 a_27908_27912# VGND 0.00388f
C34096 a_26916_27912# VGND 0.48502f
C34097 a_26468_27912# VGND 0.48974f
C34098 a_25796_27912# VGND 0.48771f
C34099 _351_.A2 VGND 0.76867f
C34100 a_24900_27912# VGND 0.00492f
C34101 a_35008_27533# VGND 0.71606f
C34102 _371_.A3 VGND 1.36226f
C34103 a_27004_27815# VGND 0.26213f
C34104 a_26556_27815# VGND 0.29118f
C34105 a_25884_27815# VGND 0.28843f
C34106 a_21044_27508# VGND 0.15997f
C34107 a_23920_27555# VGND 0.83534f
C34108 a_23627_27967# VGND 0.45901f
C34109 a_22620_27599# VGND 0.30016f
C34110 a_22992_27555# VGND 0.42064f
C34111 _454_.D VGND 0.78295f
C34112 a_22064_27912# VGND 1.48321f
C34113 _346_.ZN VGND 0.59085f
C34114 a_20308_27912# VGND 0.46155f
C34115 a_19860_27912# VGND 0.47345f
C34116 a_19412_27912# VGND 0.4663f
C34117 a_17844_27912# VGND 0.46496f
C34118 a_17396_27912# VGND 0.46114f
C34119 a_16948_27912# VGND 0.45916f
C34120 a_16500_27912# VGND 0.45916f
C34121 a_16052_27912# VGND 0.45983f
C34122 a_15604_27912# VGND 0.46751f
C34123 a_15156_27912# VGND 0.43828f
C34124 a_14708_27912# VGND 0.4664f
C34125 a_5300_27912# VGND 0.48995f
C34126 a_4852_27912# VGND 0.48956f
C34127 a_4068_27912# VGND 0.44997f
C34128 a_3620_27912# VGND 0.43828f
C34129 a_3172_27912# VGND 0.43828f
C34130 a_2724_27912# VGND 0.43828f
C34131 a_2276_27912# VGND 0.43828f
C34132 a_1828_27912# VGND 0.43828f
C34133 a_1380_27912# VGND 0.43828f
C34134 a_932_27912# VGND 0.4664f
C34135 a_20396_27815# VGND 0.26881f
C34136 a_19948_27815# VGND 0.33371f
C34137 a_19500_27815# VGND 0.29395f
C34138 a_17932_27815# VGND 0.27564f
C34139 a_17484_27815# VGND 0.28146f
C34140 a_17036_27815# VGND 0.28473f
C34141 a_16588_27815# VGND 0.2812f
C34142 a_16140_27815# VGND 0.2812f
C34143 a_15692_27815# VGND 0.2812f
C34144 a_15244_27815# VGND 0.2812f
C34145 a_14796_27815# VGND 0.29134f
C34146 a_5388_27815# VGND 0.31553f
C34147 a_4940_27815# VGND 0.29984f
C34148 a_4156_27815# VGND 0.28278f
C34149 a_3708_27815# VGND 0.2812f
C34150 a_3260_27815# VGND 0.2812f
C34151 a_2812_27815# VGND 0.2812f
C34152 a_2364_27815# VGND 0.2812f
C34153 a_1916_27815# VGND 0.2812f
C34154 a_1468_27815# VGND 0.2812f
C34155 a_1020_27815# VGND 0.29134f
C34156 a_63105_28293# VGND 0.0268f
C34157 a_62503_28293# VGND 0.04574f
C34158 vgaringosc.tapped_ring.c11_inv_array\[3\]_pdkinv_notouch_.I VGND 0.88733f
C34159 a_63721_28776# VGND 0.00383f
C34160 a_63313_28776# VGND 0.0059f
C34161 a_62763_28776# VGND 0.00124f
C34162 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.ZN VGND 0.88988f
C34163 vgaringosc.tapped_ring.c09_inv_array\[7\]_pdkinv_notouch_.I VGND 0.87738f
C34164 vgaringosc.tapped_ring.c08_inv_array\[6\]_pdkinv_notouch_.ZN VGND 0.87968f
C34165 vgaringosc.tapped_ring.c08_inv_array\[5\]_pdkinv_notouch_.ZN VGND 0.86376f
C34166 vgaringosc.tapped_ring.c11_inv_array\[15\]_pdkinv_notouch_.ZN VGND 1.9009f
C34167 _250_.A2 VGND 0.4018f
C34168 a_60940_28248# VGND 0.27292f
C34169 a_60492_28248# VGND 0.29181f
C34170 a_60059_28776# VGND 0.00263f
C34171 _243_.A1 VGND 0.64771f
C34172 _252_.B VGND 1.24808f
C34173 _241_.I0 VGND 1.31797f
C34174 a_56124_28248# VGND 0.26105f
C34175 a_55676_28248# VGND 0.28671f
C34176 a_55228_28248# VGND 0.28645f
C34177 a_60852_28292# VGND 0.46949f
C34178 a_60404_28292# VGND 0.46764f
C34179 vgaringosc.tapped_ring.c00_inv_array\[1\]_pdkinv_notouch_.I VGND 0.95235f
C34180 a_56036_28292# VGND 0.46763f
C34181 a_55588_28292# VGND 0.45991f
C34182 a_55140_28292# VGND 0.48364f
C34183 a_52891_28776# VGND 0.00252f
C34184 a_51084_28248# VGND 0.30967f
C34185 _407_.A1 VGND 1.16758f
C34186 a_50197_28776# VGND 0.00278f
C34187 a_49637_28776# VGND 0.00266f
C34188 vgaringosc.ro_inv1.inv_array_notouch_\[1\].ZN VGND 0.60245f
C34189 vgaringosc.ro_inv1.inv_array_notouch_\[2\].ZN VGND 0.52594f
C34190 a_50996_28292# VGND 0.50915f
C34191 _404_.A1 VGND 1.12506f
C34192 _395_.A1 VGND 1.99867f
C34193 _381_.Z VGND 1.03582f
C34194 _470_.Q VGND 2.03528f
C34195 _393_.A3 VGND 0.56767f
C34196 _389_.ZN VGND 0.8636f
C34197 a_45484_28248# VGND 0.29263f
C34198 a_45036_28248# VGND 0.29022f
C34199 a_39256_28292# VGND 0.00372f
C34200 a_43248_28777# VGND 0.00182f
C34201 a_42320_28777# VGND 0.00146f
C34202 a_45396_28292# VGND 0.48356f
C34203 a_44948_28292# VGND 0.48464f
C34204 a_43003_28409# VGND 0.48558f
C34205 a_43296_28733# VGND 0.87924f
C34206 a_41996_28777# VGND 0.30315f
C34207 a_42368_28733# VGND 0.42039f
C34208 _265_.ZN VGND 0.67697f
C34209 a_41440_28363# VGND 1.47984f
C34210 a_39480_28776# VGND 0.00526f
C34211 _234_.ZN VGND 0.53783f
C34212 a_40038_28720# VGND 0.98626f
C34213 a_38584_28292# VGND 0.7353f
C34214 _437_.A1 VGND 3.88324f
C34215 a_37324_28776# VGND 0.00172f
C34216 a_36828_28776# VGND 0.00158f
C34217 a_36420_28776# VGND 0.00157f
C34218 a_29575_28293# VGND 0.04718f
C34219 a_35914_28776# VGND 0.00212f
C34220 a_35710_28776# VGND 0.00534f
C34221 a_35516_28776# VGND 0.00436f
C34222 a_35108_28776# VGND 0.0041f
C34223 a_34700_28776# VGND 0.0041f
C34224 a_34292_28776# VGND 0.00504f
C34225 a_34084_28776# VGND 3.23779f
C34226 a_33720_28776# VGND 0.00503f
C34227 a_33312_28776# VGND 0.00242f
C34228 a_32904_28776# VGND 0.00242f
C34229 a_32476_28776# VGND 0.00413f
C34230 _223_.ZN VGND 1.20015f
C34231 _335_.ZN VGND 1.53319f
C34232 _371_.A1 VGND 3.26813f
C34233 a_30388_28776# VGND 3.71637f
C34234 a_29835_28776# VGND 0.00127f
C34235 _337_.ZN VGND 1.80745f
C34236 _369_.ZN VGND 0.51193f
C34237 _352_.A2 VGND 5.21113f
C34238 a_28364_28776# VGND 0.00143f
C34239 a_27868_28776# VGND 0.00358f
C34240 a_27460_28776# VGND 0.00142f
C34241 _371_.A2 VGND 1.75112f
C34242 a_26954_28776# VGND 0.00175f
C34243 a_26750_28776# VGND 0.00226f
C34244 a_26556_28776# VGND 0.00308f
C34245 a_26148_28776# VGND 0.0041f
C34246 a_25740_28776# VGND 0.0041f
C34247 a_25332_28776# VGND 0.00496f
C34248 a_25124_28776# VGND 3.23429f
C34249 a_24780_28776# VGND 0.00145f
C34250 _346_.A2 VGND 1.89295f
C34251 _345_.A2 VGND 0.54154f
C34252 _337_.A3 VGND 4.10117f
C34253 _455_.Q VGND 3.31557f
C34254 a_24392_28248# VGND 0.55798f
C34255 _454_.Q VGND 2.11148f
C34256 a_23084_28248# VGND 0.26367f
C34257 a_22636_28248# VGND 0.29465f
C34258 a_22996_28292# VGND 0.45104f
C34259 a_22548_28292# VGND 0.46485f
C34260 a_21628_28248# VGND 0.27314f
C34261 a_19280_28777# VGND 0.00146f
C34262 a_18352_28777# VGND 0.00146f
C34263 a_18028_28777# VGND 0.29666f
C34264 a_18400_28733# VGND 0.4187f
C34265 _378_.ZN VGND 0.51499f
C34266 a_17472_28363# VGND 1.4791f
C34267 a_21540_28292# VGND 0.47962f
C34268 a_19328_28733# VGND 1.74552f
C34269 a_19035_28409# VGND 0.68258f
C34270 a_16588_28248# VGND 0.24926f
C34271 a_16140_28248# VGND 0.28627f
C34272 a_15692_28248# VGND 0.2841f
C34273 a_15244_28248# VGND 0.2841f
C34274 a_14796_28248# VGND 0.2937f
C34275 a_16500_28292# VGND 0.47278f
C34276 a_16052_28292# VGND 0.46157f
C34277 a_15604_28292# VGND 0.46136f
C34278 a_15156_28292# VGND 0.46136f
C34279 a_14708_28292# VGND 0.49005f
C34280 a_5052_28248# VGND 0.28654f
C34281 a_4604_28248# VGND 0.31699f
C34282 a_4156_28248# VGND 0.29553f
C34283 a_3708_28248# VGND 0.2812f
C34284 a_3260_28248# VGND 0.2812f
C34285 a_2812_28248# VGND 0.2812f
C34286 a_2364_28248# VGND 0.2812f
C34287 a_1916_28248# VGND 0.2812f
C34288 a_1468_28248# VGND 0.2812f
C34289 a_1020_28248# VGND 0.29134f
C34290 a_4964_28292# VGND 0.49253f
C34291 a_4516_28292# VGND 0.51849f
C34292 a_4068_28292# VGND 0.44538f
C34293 a_3620_28292# VGND 0.43828f
C34294 a_3172_28292# VGND 0.43828f
C34295 a_2724_28292# VGND 0.43828f
C34296 a_2276_28292# VGND 0.43828f
C34297 a_1828_28292# VGND 0.43828f
C34298 a_1380_28292# VGND 0.43828f
C34299 a_932_28292# VGND 0.4664f
C34300 a_64220_29098# VGND 0.00231f
C34301 vgaringosc.tapped_ring.c11_inv_array\[1\]_pdkinv_notouch_.I VGND 1.07742f
C34302 vgaringosc.tapped_ring.c09_inv_array\[6\]_pdkinv_notouch_.I VGND 1.03841f
C34303 a_63524_29098# VGND 0.00477f
C34304 a_62944_29101# VGND 0.0039f
C34305 _250_.B VGND 0.94252f
C34306 a_63952_29480# VGND 0.02887f
C34307 a_61940_29076# VGND 0.7352f
C34308 a_59572_29076# VGND 0.5977f
C34309 a_59348_29076# VGND 0.00566f
C34310 a_58709_29076# VGND 0.00271f
C34311 a_63336_29480# VGND 0.01496f
C34312 _248_.B1 VGND 1.70073f
C34313 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.ZN VGND 0.88641f
C34314 _250_.C VGND 0.44298f
C34315 a_62564_29032# VGND 0.67975f
C34316 _238_.I VGND 1.00345f
C34317 _250_.ZN VGND 1.26007f
C34318 _252_.ZN VGND 1.39439f
C34319 a_60276_29032# VGND 0.97247f
C34320 _247_.ZN VGND 0.74485f
C34321 _238_.ZN VGND 0.49233f
C34322 _257_.B VGND 0.45732f
C34323 a_52756_29076# VGND 0.4195f
C34324 vgaringosc.tapped_ring.c00_inv_array\[0\]_pdkinv_notouch_.I VGND 1.06881f
C34325 a_56484_29480# VGND 0.49357f
C34326 vgaringosc.ro_inv4.inv_array_notouch_\[1\].I VGND 1.79341f
C34327 a_48859_29076# VGND 0.00247f
C34328 a_53616_29480# VGND 0.00124f
C34329 a_52068_29480# VGND 0.00168f
C34330 a_51050_29480# VGND 0.00467f
C34331 a_47733_29098# VGND 0.00124f
C34332 a_46837_29076# VGND 0.00249f
C34333 a_45040_29167# VGND 0.00181f
C34334 a_44112_29167# VGND 0.00169f
C34335 a_49652_29480# VGND 0.47996f
C34336 _392_.A2 VGND 0.66279f
C34337 _258_.ZN VGND 0.81348f
C34338 a_56572_29383# VGND 0.26328f
C34339 vgaringosc.ro_inv4.inv_array_notouch_\[3\].ZN VGND 1.67133f
C34340 _267_.ZN VGND 0.62892f
C34341 a_49740_29383# VGND 0.27577f
C34342 _402_.A1 VGND 5.35194f
C34343 _390_.ZN VGND 1.0264f
C34344 _393_.A1 VGND 1.24968f
C34345 a_47525_29480# VGND 0.05673f
C34346 _386_.A4 VGND 0.96788f
C34347 _383_.ZN VGND 0.94084f
C34348 _384_.ZN VGND 1.56947f
C34349 _386_.ZN VGND 0.98087f
C34350 _397_.A1 VGND 4.24926f
C34351 _383_.A2 VGND 0.87417f
C34352 a_45088_29123# VGND 0.84082f
C34353 a_44795_29535# VGND 0.46755f
C34354 a_43788_29167# VGND 0.3075f
C34355 a_44160_29123# VGND 0.42963f
C34356 _480_.Q VGND 0.69239f
C34357 a_43232_29480# VGND 1.51658f
C34358 a_37536_29167# VGND 0.0017f
C34359 a_36608_29167# VGND 0.00165f
C34360 a_33728_29167# VGND 0.0017f
C34361 a_32800_29167# VGND 0.00146f
C34362 a_41160_29083# VGND 1.51502f
C34363 a_37584_29123# VGND 1.14318f
C34364 a_37291_29535# VGND 0.46556f
C34365 a_36284_29167# VGND 0.30255f
C34366 a_36656_29123# VGND 0.42298f
C34367 a_35728_29480# VGND 1.48795f
C34368 _362_.B VGND 4.98112f
C34369 a_29808_29167# VGND 0.0017f
C34370 a_28880_29167# VGND 0.00164f
C34371 a_33776_29123# VGND 1.11645f
C34372 a_33483_29535# VGND 0.4643f
C34373 a_32476_29167# VGND 0.29549f
C34374 a_32848_29123# VGND 0.41972f
C34375 a_31920_29480# VGND 1.47167f
C34376 a_25340_29167# VGND 0.00145f
C34377 a_29856_29123# VGND 0.8308f
C34378 a_29563_29535# VGND 0.46455f
C34379 a_28556_29167# VGND 0.30048f
C34380 a_28928_29123# VGND 0.42688f
C34381 a_28000_29480# VGND 1.48248f
C34382 _373_.ZN VGND 0.53671f
C34383 a_21287_29076# VGND 0.00801f
C34384 a_21103_29076# VGND 0.00667f
C34385 a_24952_29032# VGND 0.58068f
C34386 a_22996_29480# VGND 0.44904f
C34387 a_22548_29480# VGND 0.44364f
C34388 a_22100_29480# VGND 0.47356f
C34389 a_21652_29480# VGND 0.46346f
C34390 _378_.I VGND 1.03556f
C34391 _340_.ZN VGND 0.46424f
C34392 _343_.A2 VGND 1.36514f
C34393 a_23084_29383# VGND 0.27518f
C34394 a_22636_29383# VGND 0.28651f
C34395 a_22188_29383# VGND 0.28705f
C34396 a_21740_29383# VGND 0.2858f
C34397 _346_.B VGND 1.23455f
C34398 _375_.Z VGND 0.61478f
C34399 a_20191_29611# VGND 0.00135f
C34400 a_18472_29076# VGND 0.00531f
C34401 a_18264_29480# VGND 0.00372f
C34402 _467_.D VGND 0.90821f
C34403 a_17060_29480# VGND 0.47819f
C34404 a_16612_29480# VGND 0.4652f
C34405 a_16164_29480# VGND 0.47687f
C34406 a_15492_29480# VGND 0.46112f
C34407 a_15044_29480# VGND 0.45729f
C34408 a_14596_29480# VGND 0.45729f
C34409 a_14148_29480# VGND 0.47318f
C34410 a_13700_29480# VGND 0.47818f
C34411 a_13252_29480# VGND 0.47983f
C34412 a_12804_29480# VGND 0.48236f
C34413 a_12356_29480# VGND 0.52071f
C34414 a_11684_29480# VGND 0.48152f
C34415 a_11236_29480# VGND 0.47513f
C34416 a_10788_29480# VGND 0.47513f
C34417 a_10340_29480# VGND 0.47513f
C34418 a_9892_29480# VGND 0.47513f
C34419 a_9444_29480# VGND 0.47513f
C34420 a_8996_29480# VGND 0.47513f
C34421 a_8548_29480# VGND 0.48718f
C34422 a_7876_29480# VGND 0.47896f
C34423 a_7428_29480# VGND 0.47513f
C34424 a_6980_29480# VGND 0.47513f
C34425 a_6532_29480# VGND 0.47513f
C34426 a_6084_29480# VGND 0.47765f
C34427 a_5636_29480# VGND 0.47605f
C34428 a_5188_29480# VGND 0.47504f
C34429 a_4740_29480# VGND 0.49434f
C34430 a_4068_29480# VGND 0.44968f
C34431 a_3620_29480# VGND 0.43828f
C34432 a_3172_29480# VGND 0.43828f
C34433 a_2724_29480# VGND 0.43828f
C34434 a_2276_29480# VGND 0.43828f
C34435 a_1828_29480# VGND 0.43828f
C34436 a_1380_29480# VGND 0.43828f
C34437 a_932_29480# VGND 0.4664f
C34438 a_20003_29611# VGND 0.57259f
C34439 a_18760_29032# VGND 0.74f
C34440 _379_.Z VGND 0.71534f
C34441 a_17148_29383# VGND 0.26917f
C34442 a_16700_29383# VGND 0.28671f
C34443 a_16252_29383# VGND 0.2919f
C34444 a_15580_29383# VGND 0.28628f
C34445 a_15132_29383# VGND 0.2812f
C34446 a_14684_29383# VGND 0.2812f
C34447 a_14236_29383# VGND 0.2812f
C34448 a_13788_29383# VGND 0.28431f
C34449 a_13340_29383# VGND 0.28588f
C34450 a_12892_29383# VGND 0.28809f
C34451 a_12444_29383# VGND 0.30384f
C34452 a_11772_29383# VGND 0.29957f
C34453 a_11324_29383# VGND 0.28756f
C34454 a_10876_29383# VGND 0.28738f
C34455 a_10428_29383# VGND 0.28618f
C34456 a_9980_29383# VGND 0.28618f
C34457 a_9532_29383# VGND 0.28725f
C34458 a_9084_29383# VGND 0.28447f
C34459 a_8636_29383# VGND 0.28944f
C34460 a_7964_29383# VGND 0.29246f
C34461 a_7516_29383# VGND 0.28618f
C34462 a_7068_29383# VGND 0.28618f
C34463 a_6620_29383# VGND 0.28725f
C34464 a_6172_29383# VGND 0.28639f
C34465 a_5724_29383# VGND 0.28851f
C34466 a_5276_29383# VGND 0.29053f
C34467 a_4828_29383# VGND 0.29748f
C34468 a_4156_29383# VGND 0.2987f
C34469 a_3708_29383# VGND 0.2812f
C34470 a_3260_29383# VGND 0.2812f
C34471 a_2812_29383# VGND 0.2812f
C34472 a_2364_29383# VGND 0.2812f
C34473 a_1916_29383# VGND 0.2812f
C34474 a_1468_29383# VGND 0.2812f
C34475 a_1020_29383# VGND 0.29134f
C34476 _249_.A2 VGND 1.55143f
C34477 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.I VGND 1.41838f
C34478 a_65072_29860# VGND 1.52828f
C34479 vgaringosc.tapped_ring.c10_inv_array\[0\]_pdkinv_notouch_.ZN VGND 0.86383f
C34480 vgaringosc.tapped_ring.c09_inv_array\[2\]_pdkinv_notouch_.ZN VGND 0.95459f
C34481 a_64412_29816# VGND 0.27044f
C34482 vgaringosc.tapped_ring.c09_inv_array\[1\]_pdkinv_notouch_.I VGND 0.90746f
C34483 a_64324_29860# VGND 0.48317f
C34484 vgaringosc.tapped_ring.c08_inv_array\[7\]_pdkinv_notouch_.ZN VGND 1.36345f
C34485 vgaringosc.tapped_ring.c10_inv_array\[6\]_pdkinv_notouch_.ZN VGND 1.35188f
C34486 vgaringosc.tapped_ring.c10_inv_array\[4\]_pdkinv_notouch_.I VGND 1.21612f
C34487 vgaringosc.tapped_ring.c10_inv_array\[5\]_pdkinv_notouch_.ZN VGND 1.08876f
C34488 vgaringosc.tapped_ring.c10_inv_array\[2\]_pdkinv_notouch_.ZN VGND 1.21557f
C34489 a_61297_30300# VGND 0.53935f
C34490 _246_.B2 VGND 1.49108f
C34491 a_57220_29861# VGND 0.01496f
C34492 a_56596_29861# VGND 0.04006f
C34493 _324_.C VGND 9.29934f
C34494 _255_.I VGND 1.25156f
C34495 a_60401_30300# VGND 0.54345f
C34496 a_59332_29816# VGND 1.14039f
C34497 a_58116_30344# VGND 0.1535f
C34498 a_57500_30344# VGND 0.00491f
C34499 _228_.ZN VGND 0.50917f
C34500 _255_.ZN VGND 1.15532f
C34501 a_56804_30344# VGND 0.00209f
C34502 _274_.A2 VGND 1.04795f
C34503 _272_.A2 VGND 0.4678f
C34504 _258_.I VGND 0.8483f
C34505 _267_.A1 VGND 0.8356f
C34506 a_52640_29860# VGND 0.00125f
C34507 a_51457_29861# VGND 0.03073f
C34508 vgaringosc.ro_inv1.inv_array_notouch_\[3\].ZN VGND 0.68106f
C34509 vgaringosc.ro_inv4.inv_array_notouch_\[3\].I VGND 1.64466f
C34510 vgaringosc.ro_inv4.inv_array_notouch_\[4\].ZN VGND 0.6351f
C34511 _267_.A2 VGND 1.51824f
C34512 _274_.A1 VGND 1.6804f
C34513 _274_.A3 VGND 0.43106f
C34514 vgaringosc.ro_inv4.inv_array_notouch_\[1\].ZN VGND 1.70735f
C34515 a_53212_29816# VGND 1.4054f
C34516 a_52073_30344# VGND 0.00418f
C34517 a_51665_30344# VGND 0.00601f
C34518 a_50032_30345# VGND 0.00146f
C34519 a_49104_30345# VGND 0.0017f
C34520 _409_.ZN VGND 0.54725f
C34521 a_49496_30345# VGND 0.41533f
C34522 a_49600_30180# VGND 0.3041f
C34523 a_49112_29885# VGND 1.47748f
C34524 _416_.A1 VGND 4.68797f
C34525 _274_.ZN VGND 0.49998f
C34526 _275_.ZN VGND 0.64755f
C34527 a_48708_29816# VGND 0.46517f
C34528 _397_.A2 VGND 4.15354f
C34529 a_46336_30345# VGND 0.00146f
C34530 a_45408_30345# VGND 0.0017f
C34531 _393_.ZN VGND 0.80516f
C34532 a_45800_30345# VGND 0.423f
C34533 a_48104_30219# VGND 1.11958f
C34534 a_45904_30180# VGND 0.30336f
C34535 a_45416_29885# VGND 1.47287f
C34536 a_45012_29816# VGND 0.46755f
C34537 a_43916_29816# VGND 0.25701f
C34538 vgaringosc.workerclkbuff_notouch_.I VGND 3.61603f
C34539 a_35818_29860# VGND 0.00338f
C34540 a_40264_30320# VGND 0.43662f
C34541 a_44632_30206# VGND 0.84092f
C34542 a_43828_29860# VGND 0.49494f
C34543 a_38472_30169# VGND 1.53973f
C34544 _288_.ZN VGND 1.77115f
C34545 _460_.Q VGND 4.4009f
C34546 _461_.D VGND 0.65541f
C34547 _294_.ZN VGND 1.85184f
C34548 _362_.ZN VGND 0.7621f
C34549 a_31040_30345# VGND 0.0017f
C34550 a_30112_30345# VGND 0.00146f
C34551 a_30795_29977# VGND 0.46824f
C34552 a_31088_30301# VGND 0.85649f
C34553 a_29788_30345# VGND 0.30432f
C34554 a_30160_30301# VGND 0.42533f
C34555 _370_.ZN VGND 1.07535f
C34556 a_29232_29931# VGND 1.47796f
C34557 _349_.A4 VGND 2.27864f
C34558 a_26672_30345# VGND 0.0017f
C34559 a_25744_30345# VGND 0.00146f
C34560 a_28054_30196# VGND 0.73808f
C34561 a_26427_29977# VGND 0.45045f
C34562 a_26720_30301# VGND 0.85644f
C34563 a_25420_30345# VGND 0.29493f
C34564 a_25792_30301# VGND 0.42009f
C34565 _342_.ZN VGND 0.69478f
C34566 a_24864_29931# VGND 1.48059f
C34567 a_23644_29816# VGND 0.27271f
C34568 a_23196_29816# VGND 0.28921f
C34569 a_20624_30345# VGND 0.0017f
C34570 a_19696_30345# VGND 0.00171f
C34571 a_19372_30345# VGND 0.32566f
C34572 a_19744_30301# VGND 0.45598f
C34573 a_18816_29931# VGND 1.50222f
C34574 _459_.CLK VGND 12.66753f
C34575 a_23556_29860# VGND 0.48589f
C34576 a_23108_29860# VGND 0.46756f
C34577 a_22560_30288# VGND 0.37636f
C34578 a_20672_30301# VGND 1.69754f
C34579 a_20379_29977# VGND 0.66937f
C34580 a_18044_29816# VGND 0.24941f
C34581 a_17596_29816# VGND 0.28603f
C34582 a_17148_29816# VGND 0.2841f
C34583 a_16700_29816# VGND 0.28728f
C34584 a_17956_29860# VGND 0.47962f
C34585 a_17508_29860# VGND 0.47738f
C34586 a_17060_29860# VGND 0.47873f
C34587 a_16612_29860# VGND 0.48794f
C34588 a_16028_29816# VGND 0.2928f
C34589 a_15580_29816# VGND 0.28584f
C34590 a_15132_29816# VGND 0.28236f
C34591 a_14684_29816# VGND 0.28236f
C34592 a_14236_29816# VGND 0.28236f
C34593 a_13788_29816# VGND 0.28547f
C34594 a_13340_29816# VGND 0.28704f
C34595 a_12892_29816# VGND 0.28925f
C34596 a_12444_29816# VGND 0.30115f
C34597 a_11996_29816# VGND 0.31019f
C34598 a_11548_29816# VGND 0.28926f
C34599 a_11100_29816# VGND 0.28922f
C34600 a_10652_29816# VGND 0.28922f
C34601 a_10204_29816# VGND 0.28922f
C34602 a_9756_29816# VGND 0.28922f
C34603 a_9308_29816# VGND 0.28922f
C34604 a_8860_29816# VGND 0.29272f
C34605 a_15940_29860# VGND 0.48862f
C34606 a_15492_29860# VGND 0.45983f
C34607 a_15044_29860# VGND 0.47278f
C34608 a_14596_29860# VGND 0.47405f
C34609 a_14148_29860# VGND 0.4754f
C34610 a_13700_29860# VGND 0.47582f
C34611 a_13252_29860# VGND 0.46445f
C34612 a_12804_29860# VGND 0.46698f
C34613 a_12356_29860# VGND 0.50364f
C34614 a_11908_29860# VGND 0.48201f
C34615 a_11460_29860# VGND 0.44029f
C34616 a_11012_29860# VGND 0.45329f
C34617 a_10564_29860# VGND 0.45848f
C34618 a_10116_29860# VGND 0.45848f
C34619 a_9668_29860# VGND 0.45999f
C34620 a_9220_29860# VGND 0.47278f
C34621 a_8772_29860# VGND 0.48737f
C34622 a_8188_29816# VGND 0.29452f
C34623 a_7740_29816# VGND 0.2927f
C34624 a_7292_29816# VGND 0.28922f
C34625 a_6844_29816# VGND 0.28922f
C34626 a_6396_29816# VGND 0.28922f
C34627 a_5948_29816# VGND 0.29226f
C34628 a_5500_29816# VGND 0.29351f
C34629 a_5052_29816# VGND 0.29285f
C34630 a_4604_29816# VGND 0.31397f
C34631 a_4156_29816# VGND 0.29327f
C34632 a_3708_29816# VGND 0.28236f
C34633 a_3260_29816# VGND 0.28236f
C34634 a_2812_29816# VGND 0.28236f
C34635 a_2364_29816# VGND 0.28236f
C34636 a_1916_29816# VGND 0.28236f
C34637 a_1468_29816# VGND 0.28236f
C34638 a_1020_29816# VGND 0.29228f
C34639 a_8100_29860# VGND 0.48734f
C34640 a_7652_29860# VGND 0.45848f
C34641 a_7204_29860# VGND 0.45848f
C34642 a_6756_29860# VGND 0.45999f
C34643 a_6308_29860# VGND 0.47329f
C34644 a_5860_29860# VGND 0.47728f
C34645 a_5412_29860# VGND 0.47904f
C34646 a_4964_29860# VGND 0.48174f
C34647 a_4516_29860# VGND 0.5146f
C34648 a_4068_29860# VGND 0.44738f
C34649 a_3620_29860# VGND 0.44029f
C34650 a_3172_29860# VGND 0.44029f
C34651 a_2724_29860# VGND 0.44029f
C34652 a_2276_29860# VGND 0.44029f
C34653 a_1828_29860# VGND 0.44029f
C34654 a_1380_29860# VGND 0.44029f
C34655 a_932_29860# VGND 0.46832f
C34656 a_67861_30644# VGND 0.00314f
C34657 a_67237_30644# VGND 0.00265f
C34658 a_61029_30644# VGND 0.00298f
C34659 a_67741_30600# VGND 0.80997f
C34660 a_67117_30600# VGND 0.79307f
C34661 _256_.A2 VGND 3.48293f
C34662 vgaringosc.tapped_ring.c09_inv_array\[5\]_pdkinv_notouch_.I VGND 1.15169f
C34663 a_64996_31048# VGND 0.49416f
C34664 _229_.I VGND 3.90652f
C34665 _230_.I VGND 4.06822f
C34666 a_60405_30644# VGND 0.00254f
C34667 a_59163_30644# VGND 0.00277f
C34668 a_58539_30644# VGND 0.00322f
C34669 a_66787_30600# VGND 0.66757f
C34670 vgaringosc.tapped_ring.c09_inv_array\[3\]_pdkinv_notouch_.ZN VGND 1.28903f
C34671 a_65084_30951# VGND 0.31211f
C34672 a_63616_31128# VGND 1.56217f
C34673 a_62532_30736# VGND 0.3536f
C34674 a_61860_30736# VGND 0.38406f
C34675 a_60909_30600# VGND 0.79486f
C34676 a_60285_30600# VGND 0.78002f
C34677 _237_.A1 VGND 1.22584f
C34678 _270_.A2 VGND 0.90596f
C34679 a_52891_30644# VGND 0.0025f
C34680 a_52267_30644# VGND 0.00312f
C34681 a_59955_30600# VGND 0.64044f
C34682 a_58911_30644# VGND 0.68558f
C34683 a_58687_31220# VGND 0.8369f
C34684 _272_.B1 VGND 0.57638f
C34685 a_56260_31048# VGND 0.492f
C34686 _268_.A1 VGND 2.00293f
C34687 _276_.A2 VGND 0.81615f
C34688 a_41708_30644# VGND 0.73169f
C34689 a_41264_30669# VGND 0.0039f
C34690 a_58063_30644# VGND 0.80459f
C34691 _251_.A1 VGND 6.62074f
C34692 a_56348_30951# VGND 0.28278f
C34693 input9.Z VGND 0.80832f
C34694 a_54432_31128# VGND 1.51203f
C34695 _474_.CLK VGND 10.40479f
C34696 a_52639_30644# VGND 0.63592f
C34697 a_52415_31220# VGND 0.78214f
C34698 vgaringosc.ro_inv1.inv_array_notouch_\[1\].I VGND 0.80598f
C34699 _268_.A2 VGND 2.29026f
C34700 a_49764_31048# VGND 0.46627f
C34701 a_49316_31048# VGND 0.46224f
C34702 a_48868_31048# VGND 0.4608f
C34703 a_48420_31048# VGND 0.47027f
C34704 a_47972_31048# VGND 0.45013f
C34705 a_47524_31048# VGND 0.4688f
C34706 a_47076_31048# VGND 0.45983f
C34707 a_46628_31048# VGND 0.47121f
C34708 a_45956_31048# VGND 0.47172f
C34709 a_45508_31048# VGND 0.46114f
C34710 a_45060_31048# VGND 0.46735f
C34711 a_44612_31048# VGND 0.46405f
C34712 a_44164_31048# VGND 0.47274f
C34713 a_43716_31048# VGND 0.46484f
C34714 a_43268_31048# VGND 0.49546f
C34715 a_42820_31048# VGND 0.48584f
C34716 _495_.I VGND 0.70898f
C34717 _293_.A2 VGND 1.57639f
C34718 _462_.D VGND 0.49404f
C34719 a_36288_31048# VGND 0.00226f
C34720 a_35652_31048# VGND 0.50116f
C34721 a_35204_31048# VGND 0.48819f
C34722 a_32508_30644# VGND 0.00255f
C34723 a_29371_30644# VGND 0.00276f
C34724 _370_.B VGND 0.81169f
C34725 a_32240_31048# VGND 0.00492f
C34726 a_51791_30644# VGND 0.75327f
C34727 _275_.A2 VGND 1.33518f
C34728 a_50436_30689# VGND 0.4849f
C34729 a_49852_30951# VGND 0.30805f
C34730 a_49404_30951# VGND 0.30341f
C34731 a_48956_30951# VGND 0.30341f
C34732 a_48508_30951# VGND 0.30341f
C34733 a_48060_30951# VGND 0.30341f
C34734 a_47612_30951# VGND 0.30341f
C34735 a_47164_30951# VGND 0.30341f
C34736 a_46716_30951# VGND 0.30712f
C34737 a_46044_30951# VGND 0.30848f
C34738 a_45596_30951# VGND 0.30341f
C34739 a_45148_30951# VGND 0.30419f
C34740 a_44700_30951# VGND 0.30708f
C34741 a_44252_30951# VGND 0.30829f
C34742 a_43804_30951# VGND 0.31041f
C34743 a_43356_30951# VGND 0.3393f
C34744 a_42908_30951# VGND 0.31434f
C34745 _388_.B VGND 2.05944f
C34746 _304_.B VGND 9.07649f
C34747 a_41056_30669# VGND 0.67088f
C34748 _284_.ZN VGND 4.50574f
C34749 _296_.ZN VGND 1.71743f
C34750 _285_.Z VGND 1.81659f
C34751 _359_.B VGND 4.89034f
C34752 _365_.ZN VGND 0.74844f
C34753 a_35740_30951# VGND 0.31706f
C34754 a_35292_30951# VGND 0.32544f
C34755 _287_.A1 VGND 6.16895f
C34756 _290_.ZN VGND 1.74857f
C34757 _363_.Z VGND 2.24554f
C34758 _334_.A1 VGND 4.60375f
C34759 _223_.I VGND 2.3275f
C34760 a_31396_31048# VGND 0.49758f
C34761 _287_.A2 VGND 1.67657f
C34762 a_29716_31048# VGND 0.48587f
C34763 _340_.A2 VGND 1.79344f
C34764 a_31484_30951# VGND 0.27976f
C34765 _294_.A2 VGND 2.90134f
C34766 _459_.Q VGND 4.31976f
C34767 a_29804_30951# VGND 0.28664f
C34768 _350_.A2 VGND 2.71103f
C34769 _373_.A2 VGND 0.71793f
C34770 a_20853_30644# VGND 0.00294f
C34771 a_26916_31048# VGND 0.46887f
C34772 a_26468_31048# VGND 0.46845f
C34773 a_26020_31048# VGND 0.47588f
C34774 a_25012_31048# VGND 0.472f
C34775 a_24564_31048# VGND 0.4802f
C34776 a_22996_31048# VGND 0.47352f
C34777 a_22548_31048# VGND 0.46732f
C34778 a_22100_31048# VGND 0.4714f
C34779 a_21652_31048# VGND 0.45961f
C34780 a_21204_31048# VGND 0.46341f
C34781 _379_.A2 VGND 1.52606f
C34782 _350_.A1 VGND 4.69467f
C34783 _371_.ZN VGND 1.0407f
C34784 a_28124_30600# VGND 0.34009f
C34785 a_27668_31048# VGND 0.37272f
C34786 a_27004_30951# VGND 0.31255f
C34787 a_26556_30951# VGND 0.30891f
C34788 a_26108_30951# VGND 0.31004f
C34789 a_25652_31048# VGND 0.33763f
C34790 a_25100_30951# VGND 0.26751f
C34791 a_24652_30951# VGND 0.31004f
C34792 a_24196_31048# VGND 0.35072f
C34793 a_23084_30951# VGND 0.29723f
C34794 a_22636_30951# VGND 0.30848f
C34795 a_22188_30951# VGND 0.3063f
C34796 a_21740_30951# VGND 0.3063f
C34797 a_21292_30951# VGND 0.30623f
C34798 a_20250_31048# VGND 0.0041f
C34799 _465_.D VGND 0.79248f
C34800 a_19076_31048# VGND 0.47641f
C34801 a_18628_31048# VGND 0.46519f
C34802 a_18180_31048# VGND 0.47391f
C34803 a_17732_31048# VGND 0.47511f
C34804 a_17284_31048# VGND 0.48242f
C34805 a_16164_31048# VGND 0.49853f
C34806 a_14820_31048# VGND 0.48212f
C34807 a_14372_31048# VGND 0.48594f
C34808 a_13364_31048# VGND 0.47114f
C34809 a_12916_31048# VGND 0.47828f
C34810 a_11460_31048# VGND 0.46054f
C34811 a_10452_31048# VGND 0.46709f
C34812 a_10004_31048# VGND 0.47035f
C34813 a_8996_31048# VGND 0.48827f
C34814 a_7540_31048# VGND 0.46984f
C34815 a_7092_31048# VGND 0.47035f
C34816 a_6084_31048# VGND 0.47835f
C34817 a_5636_31048# VGND 0.47814f
C34818 a_5188_31048# VGND 0.48024f
C34819 a_4740_31048# VGND 0.49804f
C34820 a_4068_31048# VGND 0.44968f
C34821 a_3620_31048# VGND 0.43828f
C34822 a_3172_31048# VGND 0.43828f
C34823 a_2724_31048# VGND 0.43828f
C34824 a_2276_31048# VGND 0.43828f
C34825 a_1828_31048# VGND 0.43828f
C34826 a_1380_31048# VGND 0.43828f
C34827 a_932_31048# VGND 0.4664f
C34828 _355_.C VGND 7.46373f
C34829 a_19164_30951# VGND 0.29206f
C34830 a_18716_30951# VGND 0.30848f
C34831 a_18268_30951# VGND 0.3063f
C34832 a_17820_30951# VGND 0.3063f
C34833 a_17372_30951# VGND 0.30863f
C34834 a_16916_31048# VGND 0.34718f
C34835 a_16252_30951# VGND 0.2756f
C34836 a_15460_31048# VGND 0.33366f
C34837 a_14908_30951# VGND 0.26791f
C34838 a_14460_30951# VGND 0.31004f
C34839 a_14004_31048# VGND 0.34399f
C34840 a_13452_30951# VGND 0.27173f
C34841 a_13004_30951# VGND 0.31635f
C34842 a_12548_31048# VGND 0.35588f
C34843 a_11548_30951# VGND 0.29564f
C34844 a_11091_30644# VGND 0.44264f
C34845 a_10540_30951# VGND 0.26799f
C34846 a_10092_30951# VGND 0.31012f
C34847 a_9635_30644# VGND 0.44751f
C34848 a_9084_30951# VGND 0.27014f
C34849 a_8627_30644# VGND 0.49531f
C34850 a_7628_30951# VGND 0.28951f
C34851 a_7180_30951# VGND 0.31012f
C34852 a_6723_30644# VGND 0.44868f
C34853 a_6172_30951# VGND 0.26948f
C34854 a_5724_30951# VGND 0.31035f
C34855 a_5276_30951# VGND 0.31237f
C34856 a_4828_30951# VGND 0.31876f
C34857 a_4156_30951# VGND 0.3209f
C34858 a_3708_30951# VGND 0.30341f
C34859 a_3260_30951# VGND 0.30341f
C34860 a_2812_30951# VGND 0.30341f
C34861 a_2364_30951# VGND 0.30341f
C34862 a_1916_30951# VGND 0.30341f
C34863 a_1468_30951# VGND 0.30341f
C34864 a_1020_30951# VGND 0.31355f
C34865 a_45456_30301.t1 VGND 0.04768f
C34866 a_45456_30301.t2 VGND 0.04315f
C34867 a_45456_30301.t7 VGND 0.14451f
C34868 a_45456_30301.t6 VGND 0.12749f
C34869 a_45456_30301.n0 VGND 0.16514f
C34870 a_45456_30301.n1 VGND 0.05628f
C34871 a_45456_30301.n2 VGND 0.21301f
C34872 a_45456_30301.t3 VGND 0.02032f
C34873 a_45456_30301.t5 VGND 0.12779f
C34874 a_45456_30301.t4 VGND 0.40165f
C34875 a_45456_30301.n3 VGND 0.25796f
C34876 a_45456_30301.n4 VGND 0.59021f
C34877 a_45456_30301.t0 VGND 0.1048f
C34878 _268_.A2.t0 VGND 0.04193f
C34879 _268_.A2.t1 VGND 0.01565f
C34880 _268_.A2.t6 VGND 0.0328f
C34881 _268_.A2.t7 VGND 0.04195f
C34882 _268_.A2.n0 VGND 0.0514f
C34883 _268_.A2.t2 VGND 0.01427f
C34884 _268_.A2.t5 VGND 0.04728f
C34885 _268_.A2.n1 VGND 0.05662f
C34886 _268_.A2.n2 VGND 0.41031f
C34887 _268_.A2.t9 VGND 0.04474f
C34888 _268_.A2.t4 VGND 0.04181f
C34889 _268_.A2.n3 VGND 0.06045f
C34890 _268_.A2.n4 VGND 0.19046f
C34891 _268_.A2.t8 VGND 0.04337f
C34892 _268_.A2.t3 VGND 0.03238f
C34893 _268_.A2.n5 VGND 0.05396f
C34894 _268_.A2.n6 VGND 0.32398f
C34895 _268_.A2.n7 VGND 0.11942f
C34896 _256_.A2.t2 VGND 0.05652f
C34897 _256_.A2.t3 VGND 0.0721f
C34898 _256_.A2.n0 VGND 0.11847f
C34899 _256_.A2.t0 VGND 0.08037f
C34900 _256_.A2.t1 VGND 0.06379f
C34901 _256_.A2.n1 VGND 0.18102f
C34902 a_41028_28776.t6 VGND 0.04128f
C34903 a_41028_28776.t3 VGND 0.13823f
C34904 a_41028_28776.t2 VGND 0.12194f
C34905 a_41028_28776.n0 VGND 0.15796f
C34906 a_41028_28776.n1 VGND 0.05384f
C34907 a_41028_28776.t1 VGND 0.04561f
C34908 a_41028_28776.n2 VGND 0.20374f
C34909 a_41028_28776.t7 VGND 0.01944f
C34910 a_41028_28776.t4 VGND 0.12223f
C34911 a_41028_28776.t5 VGND 0.38419f
C34912 a_41028_28776.n3 VGND 0.24674f
C34913 a_41028_28776.n4 VGND 0.56455f
C34914 a_41028_28776.t0 VGND 0.10024f
C34915 a_42484_18183.t5 VGND 0.12223f
C34916 a_42484_18183.t7 VGND 0.38419f
C34917 a_42484_18183.t3 VGND 0.01944f
C34918 a_42484_18183.n0 VGND 0.24674f
C34919 a_42484_18183.t4 VGND 0.13823f
C34920 a_42484_18183.t2 VGND 0.12232f
C34921 a_42484_18183.n1 VGND 0.15759f
C34922 a_42484_18183.t6 VGND 0.04083f
C34923 a_42484_18183.n2 VGND 0.05429f
C34924 a_42484_18183.t1 VGND 0.04561f
C34925 a_42484_18183.n3 VGND 0.20374f
C34926 a_42484_18183.n4 VGND 0.56455f
C34927 a_42484_18183.t0 VGND 0.10024f
C34928 a_35316_29159.t4 VGND 0.12223f
C34929 a_35316_29159.t3 VGND 0.38419f
C34930 a_35316_29159.t6 VGND 0.01944f
C34931 a_35316_29159.n0 VGND 0.24674f
C34932 a_35316_29159.t2 VGND 0.13823f
C34933 a_35316_29159.t7 VGND 0.12232f
C34934 a_35316_29159.n1 VGND 0.15759f
C34935 a_35316_29159.t5 VGND 0.04083f
C34936 a_35316_29159.n2 VGND 0.05429f
C34937 a_35316_29159.t1 VGND 0.04561f
C34938 a_35316_29159.n3 VGND 0.20374f
C34939 a_35316_29159.n4 VGND 0.56455f
C34940 a_35316_29159.t0 VGND 0.10024f
C34941 _288_.ZN.t2 VGND 0.01309f
C34942 _288_.ZN.t1 VGND 0.01309f
C34943 _288_.ZN.n0 VGND 0.02836f
C34944 _288_.ZN.t4 VGND 0.05053f
C34945 _288_.ZN.t6 VGND 0.10149f
C34946 _288_.ZN.n1 VGND 0.12965f
C34947 _288_.ZN.n2 VGND 0.15927f
C34948 _288_.ZN.t8 VGND 0.05053f
C34949 _288_.ZN.t9 VGND 0.05053f
C34950 _288_.ZN.n3 VGND 0.06657f
C34951 _288_.ZN.t7 VGND 0.08315f
C34952 _288_.ZN.n4 VGND 0.08368f
C34953 _288_.ZN.t10 VGND 0.08315f
C34954 _288_.ZN.n5 VGND 0.08368f
C34955 _288_.ZN.n6 VGND 0.06657f
C34956 _288_.ZN.n7 VGND 0.08915f
C34957 _288_.ZN.t3 VGND 0.05053f
C34958 _288_.ZN.t5 VGND 0.10149f
C34959 _288_.ZN.n8 VGND 0.11908f
C34960 _288_.ZN.n9 VGND 0.17709f
C34961 _288_.ZN.n10 VGND 0.21067f
C34962 _288_.ZN.t0 VGND 0.0753f
C34963 a_23892_27208.t6 VGND 0.04128f
C34964 a_23892_27208.t5 VGND 0.13823f
C34965 a_23892_27208.t3 VGND 0.12194f
C34966 a_23892_27208.n0 VGND 0.15796f
C34967 a_23892_27208.n1 VGND 0.05384f
C34968 a_23892_27208.t1 VGND 0.04561f
C34969 a_23892_27208.n2 VGND 0.20374f
C34970 a_23892_27208.t2 VGND 0.01944f
C34971 a_23892_27208.t7 VGND 0.12223f
C34972 a_23892_27208.t4 VGND 0.38419f
C34973 a_23892_27208.n3 VGND 0.24674f
C34974 a_23892_27208.n4 VGND 0.56455f
C34975 a_23892_27208.t0 VGND 0.10024f
C34976 a_28820_30344.t7 VGND 0.04128f
C34977 a_28820_30344.t3 VGND 0.13823f
C34978 a_28820_30344.t6 VGND 0.12194f
C34979 a_28820_30344.n0 VGND 0.15796f
C34980 a_28820_30344.n1 VGND 0.05384f
C34981 a_28820_30344.t1 VGND 0.04561f
C34982 a_28820_30344.n2 VGND 0.20374f
C34983 a_28820_30344.t2 VGND 0.01944f
C34984 a_28820_30344.t5 VGND 0.12223f
C34985 a_28820_30344.t4 VGND 0.38419f
C34986 a_28820_30344.n3 VGND 0.24674f
C34987 a_28820_30344.n4 VGND 0.56455f
C34988 a_28820_30344.t0 VGND 0.10024f
C34989 a_52400_25987.t5 VGND 0.12223f
C34990 a_52400_25987.t7 VGND 0.38419f
C34991 a_52400_25987.t3 VGND 0.01944f
C34992 a_52400_25987.n0 VGND 0.24674f
C34993 a_52400_25987.t1 VGND 0.04561f
C34994 a_52400_25987.t6 VGND 0.13823f
C34995 a_52400_25987.t2 VGND 0.12232f
C34996 a_52400_25987.n1 VGND 0.15759f
C34997 a_52400_25987.t4 VGND 0.04083f
C34998 a_52400_25987.n2 VGND 0.05429f
C34999 a_52400_25987.n3 VGND 0.20374f
C35000 a_52400_25987.n4 VGND 0.56455f
C35001 a_52400_25987.t0 VGND 0.10024f
C35002 _311_.A2.t8 VGND 0.06059f
C35003 _311_.A2.t11 VGND 0.08082f
C35004 _311_.A2.n0 VGND 0.10031f
C35005 _311_.A2.t2 VGND 0.0266f
C35006 _311_.A2.t5 VGND 0.08811f
C35007 _311_.A2.n1 VGND 0.10637f
C35008 _311_.A2.n2 VGND 0.23979f
C35009 _311_.A2.t3 VGND 0.09098f
C35010 _311_.A2.t6 VGND 0.05398f
C35011 _311_.A2.n3 VGND 0.09897f
C35012 _311_.A2.t4 VGND 0.0647f
C35013 _311_.A2.t10 VGND 0.04682f
C35014 _311_.A2.n4 VGND 0.10194f
C35015 _311_.A2.n5 VGND 0.26472f
C35016 _311_.A2.t9 VGND 0.02265f
C35017 _311_.A2.t7 VGND 0.08855f
C35018 _311_.A2.n6 VGND 0.11175f
C35019 _311_.A2.n7 VGND 0.21593f
C35020 _311_.A2.n8 VGND 0.70096f
C35021 _311_.A2.n9 VGND 0.65228f
C35022 _311_.A2.n10 VGND 0.3909f
C35023 _311_.A2.t0 VGND 0.07012f
C35024 _311_.A2.n11 VGND 0.09251f
C35025 _311_.A2.t1 VGND 0.0545f
C35026 a_15828_27208.t6 VGND 0.04104f
C35027 a_15828_27208.t2 VGND 0.13745f
C35028 a_15828_27208.t5 VGND 0.12126f
C35029 a_15828_27208.n0 VGND 0.15708f
C35030 a_15828_27208.n1 VGND 0.05354f
C35031 a_15828_27208.t1 VGND 0.04536f
C35032 a_15828_27208.n2 VGND 0.19884f
C35033 a_15828_27208.t3 VGND 0.01933f
C35034 a_15828_27208.t4 VGND 0.12155f
C35035 a_15828_27208.t7 VGND 0.38204f
C35036 a_15828_27208.n3 VGND 0.24693f
C35037 a_15828_27208.n4 VGND 0.58092f
C35038 a_15828_27208.t0 VGND 0.09466f
C35039 a_29828_24455.t5 VGND 0.12223f
C35040 a_29828_24455.t6 VGND 0.38419f
C35041 a_29828_24455.t3 VGND 0.01944f
C35042 a_29828_24455.n0 VGND 0.24674f
C35043 a_29828_24455.t4 VGND 0.13823f
C35044 a_29828_24455.t7 VGND 0.12232f
C35045 a_29828_24455.n1 VGND 0.15759f
C35046 a_29828_24455.t2 VGND 0.04083f
C35047 a_29828_24455.n2 VGND 0.05429f
C35048 a_29828_24455.t1 VGND 0.04561f
C35049 a_29828_24455.n3 VGND 0.20374f
C35050 a_29828_24455.n4 VGND 0.56455f
C35051 a_29828_24455.t0 VGND 0.10024f
C35052 _325_.A2.t0 VGND 0.03552f
C35053 _325_.A2.t3 VGND 0.03725f
C35054 _325_.A2.t2 VGND 0.04046f
C35055 _325_.A2.n0 VGND 0.04677f
C35056 _325_.A2.n1 VGND 0.02387f
C35057 _325_.A2.t7 VGND 0.04193f
C35058 _325_.A2.t5 VGND 0.03412f
C35059 _325_.A2.n2 VGND 0.05384f
C35060 _325_.A2.n3 VGND 0.09588f
C35061 _325_.A2.t11 VGND 0.04046f
C35062 _325_.A2.t4 VGND 0.03714f
C35063 _325_.A2.n4 VGND 0.04688f
C35064 _325_.A2.n5 VGND 0.2846f
C35065 _325_.A2.t10 VGND 0.01076f
C35066 _325_.A2.t6 VGND 0.04208f
C35067 _325_.A2.n6 VGND 0.0531f
C35068 _325_.A2.n7 VGND 0.0369f
C35069 _325_.A2.n8 VGND 0.39274f
C35070 _325_.A2.t9 VGND 0.0384f
C35071 _325_.A2.t8 VGND 0.02867f
C35072 _325_.A2.n9 VGND 0.04744f
C35073 _325_.A2.n10 VGND 0.06256f
C35074 _325_.A2.n11 VGND 0.37581f
C35075 _325_.A2.t1 VGND 0.02497f
C35076 _325_.A2.n12 VGND 0.0614f
C35077 a_35204_24455.t4 VGND 0.12779f
C35078 a_35204_24455.t6 VGND 0.40165f
C35079 a_35204_24455.t7 VGND 0.02032f
C35080 a_35204_24455.n0 VGND 0.25796f
C35081 a_35204_24455.t2 VGND 0.14451f
C35082 a_35204_24455.t3 VGND 0.12788f
C35083 a_35204_24455.n1 VGND 0.16475f
C35084 a_35204_24455.t5 VGND 0.04268f
C35085 a_35204_24455.n2 VGND 0.05675f
C35086 a_35204_24455.t1 VGND 0.04768f
C35087 a_35204_24455.n3 VGND 0.21301f
C35088 a_35204_24455.n4 VGND 0.59021f
C35089 a_35204_24455.t0 VGND 0.1048f
C35090 _337_.A3.t1 VGND 0.07066f
C35091 _337_.A3.t0 VGND 0.10024f
C35092 _337_.A3.t3 VGND 0.08141f
C35093 _337_.A3.n0 VGND 0.06781f
C35094 _337_.A3.t8 VGND 0.08141f
C35095 _337_.A3.t13 VGND 0.09408f
C35096 _337_.A3.n1 VGND 0.11237f
C35097 _337_.A3.t9 VGND 0.09408f
C35098 _337_.A3.n2 VGND 0.11237f
C35099 _337_.A3.n3 VGND 0.06492f
C35100 _337_.A3.n4 VGND 0.15498f
C35101 _337_.A3.n5 VGND 0.11121f
C35102 _337_.A3.t11 VGND 0.08141f
C35103 _337_.A3.t14 VGND 0.09408f
C35104 _337_.A3.t6 VGND 0.08141f
C35105 _337_.A3.n6 VGND 0.06492f
C35106 _337_.A3.t15 VGND 0.09408f
C35107 _337_.A3.n7 VGND 0.11237f
C35108 _337_.A3.n8 VGND 0.11237f
C35109 _337_.A3.n9 VGND 0.06492f
C35110 _337_.A3.n10 VGND 0.05946f
C35111 _337_.A3.t4 VGND 0.09821f
C35112 _337_.A3.t12 VGND 0.09622f
C35113 _337_.A3.n11 VGND 0.13345f
C35114 _337_.A3.n12 VGND 0.72028f
C35115 _337_.A3.t10 VGND 0.09302f
C35116 _337_.A3.t7 VGND 0.10812f
C35117 _337_.A3.n13 VGND 0.12831f
C35118 _337_.A3.t2 VGND 0.0858f
C35119 _337_.A3.t5 VGND 0.11053f
C35120 _337_.A3.n14 VGND 0.12646f
C35121 _337_.A3.n15 VGND 0.3919f
C35122 _337_.A3.n16 VGND 0.52681f
C35123 a_52064_19715.t7 VGND 0.12223f
C35124 a_52064_19715.t5 VGND 0.38419f
C35125 a_52064_19715.t3 VGND 0.01944f
C35126 a_52064_19715.n0 VGND 0.24674f
C35127 a_52064_19715.t1 VGND 0.04561f
C35128 a_52064_19715.t2 VGND 0.13823f
C35129 a_52064_19715.t4 VGND 0.12232f
C35130 a_52064_19715.n1 VGND 0.15759f
C35131 a_52064_19715.t6 VGND 0.04083f
C35132 a_52064_19715.n2 VGND 0.05429f
C35133 a_52064_19715.n3 VGND 0.20374f
C35134 a_52064_19715.n4 VGND 0.56455f
C35135 a_52064_19715.t0 VGND 0.10024f
C35136 _451_.Q.t0 VGND 0.0669f
C35137 _451_.Q.t1 VGND 0.04716f
C35138 _451_.Q.t15 VGND 0.07016f
C35139 _451_.Q.t8 VGND 0.06068f
C35140 _451_.Q.n0 VGND 0.08237f
C35141 _451_.Q.t10 VGND 0.04521f
C35142 _451_.Q.t6 VGND 0.07586f
C35143 _451_.Q.n1 VGND 0.07993f
C35144 _451_.Q.n2 VGND 0.07207f
C35145 _451_.Q.n3 VGND 0.89422f
C35146 _451_.Q.t4 VGND 0.05395f
C35147 _451_.Q.t7 VGND 0.03904f
C35148 _451_.Q.n4 VGND 0.085f
C35149 _451_.Q.t2 VGND 0.05543f
C35150 _451_.Q.t9 VGND 0.07441f
C35151 _451_.Q.n5 VGND 0.0887f
C35152 _451_.Q.n6 VGND 0.28261f
C35153 _451_.Q.n7 VGND 0.82272f
C35154 _451_.Q.t17 VGND 0.07101f
C35155 _451_.Q.t14 VGND 0.06518f
C35156 _451_.Q.n8 VGND 0.08269f
C35157 _451_.Q.n9 VGND 0.07111f
C35158 _451_.Q.n10 VGND 0.3906f
C35159 _451_.Q.t13 VGND 0.0534f
C35160 _451_.Q.t11 VGND 0.04171f
C35161 _451_.Q.n11 VGND 0.08727f
C35162 _451_.Q.n12 VGND 0.16944f
C35163 _451_.Q.t5 VGND 0.07101f
C35164 _451_.Q.t12 VGND 0.06353f
C35165 _451_.Q.n13 VGND 0.08638f
C35166 _451_.Q.t16 VGND 0.04052f
C35167 _451_.Q.t3 VGND 0.05561f
C35168 _451_.Q.n14 VGND 0.09066f
C35169 _451_.Q.n15 VGND 0.06734f
C35170 _451_.Q.n16 VGND 0.2761f
C35171 _397_.A1.t0 VGND 0.02965f
C35172 _397_.A1.t1 VGND 0.0209f
C35173 _397_.A1.t10 VGND 0.01758f
C35174 _397_.A1.t12 VGND 0.03232f
C35175 _397_.A1.n0 VGND 0.03367f
C35176 _397_.A1.t7 VGND 0.01518f
C35177 _397_.A1.t13 VGND 0.03063f
C35178 _397_.A1.n1 VGND 0.0486f
C35179 _397_.A1.n2 VGND 0.13722f
C35180 _397_.A1.t15 VGND 0.03248f
C35181 _397_.A1.t17 VGND 0.02527f
C35182 _397_.A1.n3 VGND 0.03662f
C35183 _397_.A1.t11 VGND 0.0224f
C35184 _397_.A1.t4 VGND 0.03093f
C35185 _397_.A1.n4 VGND 0.0393f
C35186 _397_.A1.n5 VGND 0.25963f
C35187 _397_.A1.n6 VGND 0.37364f
C35188 _397_.A1.t5 VGND 0.02115f
C35189 _397_.A1.n7 VGND 0.01974f
C35190 _397_.A1.t8 VGND 0.02963f
C35191 _397_.A1.t14 VGND 0.02963f
C35192 _397_.A1.n8 VGND 0.025f
C35193 _397_.A1.n9 VGND 0.025f
C35194 _397_.A1.t6 VGND 0.02115f
C35195 _397_.A1.n10 VGND 0.01919f
C35196 _397_.A1.n11 VGND 0.0488f
C35197 _397_.A1.n12 VGND 0.14904f
C35198 _397_.A1.t3 VGND 0.03746f
C35199 _397_.A1.t16 VGND 0.02179f
C35200 _397_.A1.n13 VGND 0.03798f
C35201 _397_.A1.t2 VGND 0.02383f
C35202 _397_.A1.t9 VGND 0.02283f
C35203 _397_.A1.n14 VGND 0.04352f
C35204 _397_.A1.n15 VGND 0.02665f
C35205 _397_.A1.n16 VGND 0.06444f
C35206 _397_.A1.n17 VGND 0.2027f
C35207 a_53744_22851.t3 VGND 0.12223f
C35208 a_53744_22851.t6 VGND 0.38419f
C35209 a_53744_22851.t7 VGND 0.01944f
C35210 a_53744_22851.n0 VGND 0.24674f
C35211 a_53744_22851.t1 VGND 0.04561f
C35212 a_53744_22851.t4 VGND 0.13823f
C35213 a_53744_22851.t5 VGND 0.12232f
C35214 a_53744_22851.n1 VGND 0.15759f
C35215 a_53744_22851.t2 VGND 0.04083f
C35216 a_53744_22851.n2 VGND 0.05429f
C35217 a_53744_22851.n3 VGND 0.20374f
C35218 a_53744_22851.n4 VGND 0.56455f
C35219 a_53744_22851.t0 VGND 0.10024f
C35220 _284_.A2.t1 VGND 0.02927f
C35221 _284_.A2.t3 VGND 0.04721f
C35222 _284_.A2.t4 VGND 0.03937f
C35223 _284_.A2.n0 VGND 0.0669f
C35224 _284_.A2.n1 VGND 0.08992f
C35225 _284_.A2.t7 VGND 0.03188f
C35226 _284_.A2.t5 VGND 0.03937f
C35227 _284_.A2.n2 VGND 0.02824f
C35228 _284_.A2.n3 VGND 0.03984f
C35229 _284_.A2.t6 VGND 0.03188f
C35230 _284_.A2.n4 VGND 0.03984f
C35231 _284_.A2.t8 VGND 0.03937f
C35232 _284_.A2.n5 VGND 0.02824f
C35233 _284_.A2.n6 VGND 0.02542f
C35234 _284_.A2.t2 VGND 0.04497f
C35235 _284_.A2.t9 VGND 0.04095f
C35236 _284_.A2.n7 VGND 0.06652f
C35237 _284_.A2.t0 VGND 0.03766f
C35238 _284_.A2.n8 VGND 0.5649f
C35239 a_32180_25640.t7 VGND 0.04315f
C35240 a_32180_25640.t3 VGND 0.14451f
C35241 a_32180_25640.t2 VGND 0.12749f
C35242 a_32180_25640.n0 VGND 0.16514f
C35243 a_32180_25640.n1 VGND 0.05628f
C35244 a_32180_25640.t1 VGND 0.04768f
C35245 a_32180_25640.n2 VGND 0.21301f
C35246 a_32180_25640.t5 VGND 0.02032f
C35247 a_32180_25640.t4 VGND 0.12779f
C35248 a_32180_25640.t6 VGND 0.40165f
C35249 a_32180_25640.n3 VGND 0.25796f
C35250 a_32180_25640.n4 VGND 0.59021f
C35251 a_32180_25640.t0 VGND 0.1048f
C35252 a_28596_27916.t7 VGND 0.15904f
C35253 a_28596_27916.t4 VGND 0.05118f
C35254 a_28596_27916.t5 VGND 0.05118f
C35255 a_28596_27916.n0 VGND 0.10237f
C35256 a_28596_27916.n1 VGND 0.4343f
C35257 a_28596_27916.t1 VGND 0.05118f
C35258 a_28596_27916.t6 VGND 0.1063f
C35259 a_28596_27916.n2 VGND 0.15749f
C35260 a_28596_27916.n3 VGND 0.20525f
C35261 a_28596_27916.t10 VGND 0.05118f
C35262 a_28596_27916.t8 VGND 0.05118f
C35263 a_28596_27916.n4 VGND 0.10237f
C35264 a_28596_27916.n5 VGND 0.15394f
C35265 a_28596_27916.t0 VGND 0.05118f
C35266 a_28596_27916.t2 VGND 0.05118f
C35267 a_28596_27916.n6 VGND 0.10237f
C35268 a_28596_27916.n7 VGND 0.15394f
C35269 a_28596_27916.t9 VGND 0.05118f
C35270 a_28596_27916.t11 VGND 0.05118f
C35271 a_28596_27916.n8 VGND 0.10237f
C35272 a_28596_27916.n9 VGND 0.30161f
C35273 a_28596_27916.t3 VGND 0.15801f
C35274 _363_.Z.t1 VGND 0.02979f
C35275 _363_.Z.t0 VGND 0.04333f
C35276 _363_.Z.t3 VGND 0.0529f
C35277 _363_.Z.t6 VGND 0.03965f
C35278 _363_.Z.n0 VGND 0.06483f
C35279 _363_.Z.t9 VGND 0.03561f
C35280 _363_.Z.t5 VGND 0.03199f
C35281 _363_.Z.n1 VGND 0.06626f
C35282 _363_.Z.n2 VGND 0.13639f
C35283 _363_.Z.t7 VGND 0.04547f
C35284 _363_.Z.t2 VGND 0.04939f
C35285 _363_.Z.n3 VGND 0.0571f
C35286 _363_.Z.n4 VGND 0.05107f
C35287 _363_.Z.t8 VGND 0.03514f
C35288 _363_.Z.t4 VGND 0.04688f
C35289 _363_.Z.n5 VGND 0.05811f
C35290 _363_.Z.n6 VGND 0.05252f
C35291 _363_.Z.n7 VGND 0.40954f
C35292 _363_.Z.n8 VGND 0.50826f
C35293 a_33748_20936.t3 VGND 0.04315f
C35294 a_33748_20936.t6 VGND 0.14451f
C35295 a_33748_20936.t5 VGND 0.12749f
C35296 a_33748_20936.n0 VGND 0.16514f
C35297 a_33748_20936.n1 VGND 0.05628f
C35298 a_33748_20936.t1 VGND 0.04768f
C35299 a_33748_20936.n2 VGND 0.21301f
C35300 a_33748_20936.t4 VGND 0.02032f
C35301 a_33748_20936.t7 VGND 0.12779f
C35302 a_33748_20936.t2 VGND 0.40165f
C35303 a_33748_20936.n3 VGND 0.25796f
C35304 a_33748_20936.n4 VGND 0.59021f
C35305 a_33748_20936.t0 VGND 0.1048f
C35306 a_35092_19368.t4 VGND 0.04315f
C35307 a_35092_19368.t2 VGND 0.14451f
C35308 a_35092_19368.t6 VGND 0.12749f
C35309 a_35092_19368.n0 VGND 0.16514f
C35310 a_35092_19368.n1 VGND 0.05628f
C35311 a_35092_19368.t1 VGND 0.04768f
C35312 a_35092_19368.n2 VGND 0.21301f
C35313 a_35092_19368.t5 VGND 0.02032f
C35314 a_35092_19368.t3 VGND 0.12779f
C35315 a_35092_19368.t7 VGND 0.40165f
C35316 a_35092_19368.n3 VGND 0.25796f
C35317 a_35092_19368.n4 VGND 0.59021f
C35318 a_35092_19368.t0 VGND 0.1048f
C35319 a_31508_29159.t6 VGND 0.12223f
C35320 a_31508_29159.t3 VGND 0.38419f
C35321 a_31508_29159.t4 VGND 0.01944f
C35322 a_31508_29159.n0 VGND 0.24674f
C35323 a_31508_29159.t7 VGND 0.13823f
C35324 a_31508_29159.t5 VGND 0.12232f
C35325 a_31508_29159.n1 VGND 0.15759f
C35326 a_31508_29159.t2 VGND 0.04083f
C35327 a_31508_29159.n2 VGND 0.05429f
C35328 a_31508_29159.t1 VGND 0.04561f
C35329 a_31508_29159.n3 VGND 0.20374f
C35330 a_31508_29159.n4 VGND 0.56455f
C35331 a_31508_29159.t0 VGND 0.10024f
C35332 a_32740_22504.t4 VGND 0.04315f
C35333 a_32740_22504.t5 VGND 0.14451f
C35334 a_32740_22504.t2 VGND 0.12749f
C35335 a_32740_22504.n0 VGND 0.16514f
C35336 a_32740_22504.n1 VGND 0.05628f
C35337 a_32740_22504.t1 VGND 0.04768f
C35338 a_32740_22504.n2 VGND 0.21301f
C35339 a_32740_22504.t7 VGND 0.02032f
C35340 a_32740_22504.t6 VGND 0.12779f
C35341 a_32740_22504.t3 VGND 0.40165f
C35342 a_32740_22504.n3 VGND 0.25796f
C35343 a_32740_22504.n4 VGND 0.59021f
C35344 a_32740_22504.t0 VGND 0.1048f
C35345 a_21652_27591.t4 VGND 0.12223f
C35346 a_21652_27591.t7 VGND 0.38419f
C35347 a_21652_27591.t5 VGND 0.01944f
C35348 a_21652_27591.n0 VGND 0.24674f
C35349 a_21652_27591.t2 VGND 0.13823f
C35350 a_21652_27591.t3 VGND 0.12232f
C35351 a_21652_27591.n1 VGND 0.15759f
C35352 a_21652_27591.t6 VGND 0.04083f
C35353 a_21652_27591.n2 VGND 0.05429f
C35354 a_21652_27591.t1 VGND 0.04561f
C35355 a_21652_27591.n3 VGND 0.20374f
C35356 a_21652_27591.n4 VGND 0.56455f
C35357 a_21652_27591.t0 VGND 0.10024f
C35358 _294_.A2.t1 VGND 0.01414f
C35359 _294_.A2.t0 VGND 0.03714f
C35360 _294_.A2.t8 VGND 0.02577f
C35361 _294_.A2.t2 VGND 0.04324f
C35362 _294_.A2.n0 VGND 0.04693f
C35363 _294_.A2.t5 VGND 0.02577f
C35364 _294_.A2.t9 VGND 0.04324f
C35365 _294_.A2.n1 VGND 0.04556f
C35366 _294_.A2.n2 VGND 0.02851f
C35367 _294_.A2.t6 VGND 0.04324f
C35368 _294_.A2.t3 VGND 0.02565f
C35369 _294_.A2.n3 VGND 0.04567f
C35370 _294_.A2.n4 VGND 0.2012f
C35371 _294_.A2.n5 VGND 0.5202f
C35372 _294_.A2.t7 VGND 0.04324f
C35373 _294_.A2.t4 VGND 0.02565f
C35374 _294_.A2.n6 VGND 0.04567f
C35375 _294_.A2.n7 VGND 0.02966f
C35376 _294_.A2.n8 VGND 0.45692f
C35377 _294_.A2.n9 VGND 0.5596f
C35378 _411_.A2.t5 VGND 0.01165f
C35379 _411_.A2.t7 VGND 0.01165f
C35380 _411_.A2.n0 VGND 0.02683f
C35381 _411_.A2.t0 VGND 0.01165f
C35382 _411_.A2.t1 VGND 0.01165f
C35383 _411_.A2.n1 VGND 0.02329f
C35384 _411_.A2.n2 VGND 0.06711f
C35385 _411_.A2.t6 VGND 0.01165f
C35386 _411_.A2.t4 VGND 0.01165f
C35387 _411_.A2.n3 VGND 0.02329f
C35388 _411_.A2.n4 VGND 0.04994f
C35389 _411_.A2.t13 VGND 0.04013f
C35390 _411_.A2.t11 VGND 0.04414f
C35391 _411_.A2.n5 VGND 0.05184f
C35392 _411_.A2.t12 VGND 0.0332f
C35393 _411_.A2.t9 VGND 0.0318f
C35394 _411_.A2.n6 VGND 0.06103f
C35395 _411_.A2.n7 VGND 0.09154f
C35396 _411_.A2.t8 VGND 0.04525f
C35397 _411_.A2.t14 VGND 0.0352f
C35398 _411_.A2.n8 VGND 0.05102f
C35399 _411_.A2.n9 VGND 0.28628f
C35400 _411_.A2.t15 VGND 0.02791f
C35401 _411_.A2.t10 VGND 0.04684f
C35402 _411_.A2.n10 VGND 0.05084f
C35403 _411_.A2.n11 VGND 0.32283f
C35404 _411_.A2.n12 VGND 0.11716f
C35405 _411_.A2.t2 VGND 0.0097f
C35406 _411_.A2.t3 VGND 0.0097f
C35407 _411_.A2.n13 VGND 0.0217f
C35408 _281_.ZN.t3 VGND 0.01156f
C35409 _281_.ZN.t2 VGND 0.01156f
C35410 _281_.ZN.n0 VGND 0.02607f
C35411 _281_.ZN.t4 VGND 0.02771f
C35412 _281_.ZN.t9 VGND 0.0465f
C35413 _281_.ZN.n1 VGND 0.05047f
C35414 _281_.ZN.t6 VGND 0.03439f
C35415 _281_.ZN.t5 VGND 0.03273f
C35416 _281_.ZN.n2 VGND 0.06408f
C35417 _281_.ZN.n3 VGND 0.46949f
C35418 _281_.ZN.t8 VGND 0.03296f
C35419 _281_.ZN.t7 VGND 0.03542f
C35420 _281_.ZN.n4 VGND 0.06129f
C35421 _281_.ZN.n5 VGND 0.02621f
C35422 _281_.ZN.n6 VGND 0.44828f
C35423 _281_.ZN.t1 VGND 0.02705f
C35424 _281_.ZN.n7 VGND 0.34199f
C35425 _281_.ZN.t0 VGND 0.02801f
C35426 _281_.ZN.n8 VGND 0.06539f
C35427 a_49936_19325.t1 VGND 0.04768f
C35428 a_49936_19325.t6 VGND 0.04315f
C35429 a_49936_19325.t2 VGND 0.14451f
C35430 a_49936_19325.t7 VGND 0.12749f
C35431 a_49936_19325.n0 VGND 0.16514f
C35432 a_49936_19325.n1 VGND 0.05628f
C35433 a_49936_19325.n2 VGND 0.21301f
C35434 a_49936_19325.t4 VGND 0.02032f
C35435 a_49936_19325.t5 VGND 0.12779f
C35436 a_49936_19325.t3 VGND 0.40165f
C35437 a_49936_19325.n3 VGND 0.25796f
C35438 a_49936_19325.n4 VGND 0.59021f
C35439 a_49936_19325.t0 VGND 0.1048f
C35440 _417_.A2.t1 VGND 0.01311f
C35441 _417_.A2.t0 VGND 0.01311f
C35442 _417_.A2.n0 VGND 0.03192f
C35443 _417_.A2.t2 VGND 0.02783f
C35444 _417_.A2.t6 VGND 0.03627f
C35445 _417_.A2.t3 VGND 0.04457f
C35446 _417_.A2.n1 VGND 0.05701f
C35447 _417_.A2.n2 VGND 0.06973f
C35448 _417_.A2.t9 VGND 0.03234f
C35449 _417_.A2.t10 VGND 0.03399f
C35450 _417_.A2.n3 VGND 0.06296f
C35451 _417_.A2.n4 VGND 0.02878f
C35452 _417_.A2.n5 VGND 0.30062f
C35453 _417_.A2.t5 VGND 0.03937f
C35454 _417_.A2.t11 VGND 0.0433f
C35455 _417_.A2.n6 VGND 0.05205f
C35456 _417_.A2.t12 VGND 0.03257f
C35457 _417_.A2.t8 VGND 0.0312f
C35458 _417_.A2.n7 VGND 0.05987f
C35459 _417_.A2.n8 VGND 0.18035f
C35460 _417_.A2.n9 VGND 0.47757f
C35461 _417_.A2.t7 VGND 0.04595f
C35462 _417_.A2.t4 VGND 0.02726f
C35463 _417_.A2.n10 VGND 0.04888f
C35464 _417_.A2.n11 VGND 0.035f
C35465 _417_.A2.n12 VGND 0.31032f
C35466 a_18404_30344.t6 VGND 0.04291f
C35467 a_18404_30344.t4 VGND 0.1437f
C35468 a_18404_30344.t5 VGND 0.12677f
C35469 a_18404_30344.n0 VGND 0.16422f
C35470 a_18404_30344.n1 VGND 0.05597f
C35471 a_18404_30344.t1 VGND 0.04742f
C35472 a_18404_30344.n2 VGND 0.20788f
C35473 a_18404_30344.t3 VGND 0.02021f
C35474 a_18404_30344.t2 VGND 0.12707f
C35475 a_18404_30344.t7 VGND 0.39941f
C35476 a_18404_30344.n3 VGND 0.25815f
C35477 a_18404_30344.n4 VGND 0.60733f
C35478 a_18404_30344.t0 VGND 0.09896f
C35479 a_42596_27208.t4 VGND 0.04315f
C35480 a_42596_27208.t2 VGND 0.14451f
C35481 a_42596_27208.t7 VGND 0.12749f
C35482 a_42596_27208.n0 VGND 0.16514f
C35483 a_42596_27208.n1 VGND 0.05628f
C35484 a_42596_27208.t1 VGND 0.04768f
C35485 a_42596_27208.n2 VGND 0.21301f
C35486 a_42596_27208.t6 VGND 0.02032f
C35487 a_42596_27208.t3 VGND 0.12779f
C35488 a_42596_27208.t5 VGND 0.40165f
C35489 a_42596_27208.n3 VGND 0.25796f
C35490 a_42596_27208.n4 VGND 0.59021f
C35491 a_42596_27208.t0 VGND 0.1048f
C35492 _294_.ZN.t1 VGND 0.04914f
C35493 _294_.ZN.t10 VGND 0.03434f
C35494 _294_.ZN.t3 VGND 0.06897f
C35495 _294_.ZN.n0 VGND 0.08811f
C35496 _294_.ZN.n1 VGND 0.10824f
C35497 _294_.ZN.t6 VGND 0.03434f
C35498 _294_.ZN.t7 VGND 0.03434f
C35499 _294_.ZN.n2 VGND 0.04524f
C35500 _294_.ZN.t8 VGND 0.05651f
C35501 _294_.ZN.n3 VGND 0.05687f
C35502 _294_.ZN.t9 VGND 0.05651f
C35503 _294_.ZN.n4 VGND 0.05687f
C35504 _294_.ZN.n5 VGND 0.04524f
C35505 _294_.ZN.n6 VGND 0.06059f
C35506 _294_.ZN.t4 VGND 0.03434f
C35507 _294_.ZN.t5 VGND 0.06897f
C35508 _294_.ZN.n7 VGND 0.08093f
C35509 _294_.ZN.n8 VGND 0.44497f
C35510 _294_.ZN.n9 VGND 0.46755f
C35511 _294_.ZN.t2 VGND 0.0089f
C35512 _294_.ZN.t0 VGND 0.0089f
C35513 _294_.ZN.n10 VGND 0.02214f
C35514 a_32964_24072.t2 VGND 0.04315f
C35515 a_32964_24072.t5 VGND 0.14451f
C35516 a_32964_24072.t4 VGND 0.12749f
C35517 a_32964_24072.n0 VGND 0.16514f
C35518 a_32964_24072.n1 VGND 0.05628f
C35519 a_32964_24072.t1 VGND 0.04768f
C35520 a_32964_24072.n2 VGND 0.21301f
C35521 a_32964_24072.t3 VGND 0.02032f
C35522 a_32964_24072.t6 VGND 0.12779f
C35523 a_32964_24072.t7 VGND 0.40165f
C35524 a_32964_24072.n3 VGND 0.25796f
C35525 a_32964_24072.n4 VGND 0.59021f
C35526 a_32964_24072.t0 VGND 0.1048f
C35527 a_24452_30344.t4 VGND 0.04315f
C35528 a_24452_30344.t6 VGND 0.14451f
C35529 a_24452_30344.t3 VGND 0.12749f
C35530 a_24452_30344.n0 VGND 0.16514f
C35531 a_24452_30344.n1 VGND 0.05628f
C35532 a_24452_30344.t1 VGND 0.04768f
C35533 a_24452_30344.n2 VGND 0.21301f
C35534 a_24452_30344.t2 VGND 0.02032f
C35535 a_24452_30344.t7 VGND 0.12779f
C35536 a_24452_30344.t5 VGND 0.40165f
C35537 a_24452_30344.n3 VGND 0.25796f
C35538 a_24452_30344.n4 VGND 0.59021f
C35539 a_24452_30344.t0 VGND 0.1048f
C35540 a_41088_17757.t1 VGND 0.04768f
C35541 a_41088_17757.t5 VGND 0.04315f
C35542 a_41088_17757.t3 VGND 0.14451f
C35543 a_41088_17757.t6 VGND 0.12749f
C35544 a_41088_17757.n0 VGND 0.16514f
C35545 a_41088_17757.n1 VGND 0.05628f
C35546 a_41088_17757.n2 VGND 0.21301f
C35547 a_41088_17757.t4 VGND 0.02032f
C35548 a_41088_17757.t7 VGND 0.12779f
C35549 a_41088_17757.t2 VGND 0.40165f
C35550 a_41088_17757.n3 VGND 0.25796f
C35551 a_41088_17757.n4 VGND 0.59021f
C35552 a_41088_17757.t0 VGND 0.1048f
C35553 _336_.A2.t1 VGND 0.05803f
C35554 _336_.A2.t0 VGND 0.08232f
C35555 _336_.A2.t8 VGND 0.04828f
C35556 _336_.A2.t2 VGND 0.06639f
C35557 _336_.A2.n0 VGND 0.10357f
C35558 _336_.A2.n1 VGND 0.1701f
C35559 _336_.A2.t5 VGND 0.08737f
C35560 _336_.A2.t9 VGND 0.08021f
C35561 _336_.A2.n2 VGND 0.10124f
C35562 _336_.A2.n3 VGND 0.10349f
C35563 _336_.A2.t3 VGND 0.07636f
C35564 _336_.A2.t11 VGND 0.08434f
C35565 _336_.A2.n4 VGND 0.11167f
C35566 _336_.A2.t10 VGND 0.09403f
C35567 _336_.A2.t12 VGND 0.06377f
C35568 _336_.A2.n5 VGND 0.1073f
C35569 _336_.A2.n6 VGND 0.08859f
C35570 _336_.A2.n7 VGND 0.60973f
C35571 _336_.A2.n8 VGND 0.45417f
C35572 _336_.A2.t7 VGND 0.0784f
C35573 _336_.A2.t6 VGND 0.08737f
C35574 _336_.A2.n9 VGND 0.10607f
C35575 _336_.A2.t4 VGND 0.06843f
C35576 _336_.A2.t13 VGND 0.04986f
C35577 _336_.A2.n10 VGND 0.11155f
C35578 _336_.A2.n11 VGND 0.07696f
C35579 _336_.A2.n12 VGND 0.43618f
C35580 a_44784_25987.t7 VGND 0.12779f
C35581 a_44784_25987.t5 VGND 0.40165f
C35582 a_44784_25987.t4 VGND 0.02032f
C35583 a_44784_25987.n0 VGND 0.25796f
C35584 a_44784_25987.t1 VGND 0.04768f
C35585 a_44784_25987.t3 VGND 0.14451f
C35586 a_44784_25987.t2 VGND 0.12788f
C35587 a_44784_25987.n1 VGND 0.16475f
C35588 a_44784_25987.t6 VGND 0.04268f
C35589 a_44784_25987.n2 VGND 0.05675f
C35590 a_44784_25987.n3 VGND 0.21301f
C35591 a_44784_25987.n4 VGND 0.59021f
C35592 a_44784_25987.t0 VGND 0.1048f
C35593 uo_out[7].t1 VGND 0.01791f
C35594 uo_out[7].t0 VGND 0.01294f
C35595 uo_out[7].n0 VGND 0.03325f
C35596 uo_out[7].t3 VGND 0.00869f
C35597 uo_out[7].t5 VGND 0.00869f
C35598 uo_out[7].n1 VGND 0.02025f
C35599 uo_out[7].t4 VGND 0.02444f
C35600 uo_out[7].n2 VGND 0.65796f
C35601 uo_out[7].n3 VGND 0.0796f
C35602 uo_out[7].t2 VGND 0.03338f
C35603 uo_out[7].n4 VGND 0.10239f
C35604 _384_.A3.t6 VGND 0.06816f
C35605 _384_.A3.t9 VGND 0.02243f
C35606 _384_.A3.t4 VGND 0.02243f
C35607 _384_.A3.n0 VGND 0.04487f
C35608 _384_.A3.n1 VGND 0.26443f
C35609 _384_.A3.t1 VGND 0.02243f
C35610 _384_.A3.t0 VGND 0.02243f
C35611 _384_.A3.n2 VGND 0.04487f
C35612 _384_.A3.n3 VGND 0.09026f
C35613 _384_.A3.t2 VGND 0.02177f
C35614 _384_.A3.t3 VGND 0.02177f
C35615 _384_.A3.n4 VGND 0.08029f
C35616 _384_.A3.t7 VGND 0.06103f
C35617 _384_.A3.n5 VGND 0.43192f
C35618 _384_.A3.t5 VGND 0.02243f
C35619 _384_.A3.t8 VGND 0.02243f
C35620 _384_.A3.n6 VGND 0.04487f
C35621 _384_.A3.n7 VGND 0.09512f
C35622 _384_.A3.t12 VGND 0.05439f
C35623 _384_.A3.t10 VGND 0.0748f
C35624 _384_.A3.n8 VGND 0.11758f
C35625 _384_.A3.t15 VGND 0.08302f
C35626 _384_.A3.t17 VGND 0.10202f
C35627 _384_.A3.n9 VGND 0.13091f
C35628 _384_.A3.n10 VGND 0.94145f
C35629 _384_.A3.t11 VGND 0.07403f
C35630 _384_.A3.t13 VGND 0.07779f
C35631 _384_.A3.n11 VGND 0.14493f
C35632 _384_.A3.n12 VGND 0.203f
C35633 _384_.A3.t14 VGND 0.07004f
C35634 _384_.A3.t16 VGND 0.09343f
C35635 _384_.A3.n13 VGND 0.11509f
C35636 _384_.A3.n14 VGND 0.29366f
C35637 _384_.A3.n15 VGND 0.56343f
C35638 _384_.A3.n16 VGND 0.07317f
C35639 _424_.A2.t0 VGND 0.0151f
C35640 _424_.A2.t3 VGND 0.0151f
C35641 _424_.A2.n0 VGND 0.03075f
C35642 _424_.A2.t4 VGND 0.01096f
C35643 _424_.A2.t5 VGND 0.01096f
C35644 _424_.A2.n1 VGND 0.02571f
C35645 _424_.A2.t13 VGND 0.04393f
C35646 _424_.A2.t6 VGND 0.05017f
C35647 _424_.A2.n2 VGND 0.06262f
C35648 _424_.A2.n3 VGND 0.41105f
C35649 _424_.A2.t7 VGND 0.04578f
C35650 _424_.A2.t12 VGND 0.0482f
C35651 _424_.A2.n4 VGND 0.0648f
C35652 _424_.A2.n5 VGND 0.21063f
C35653 _424_.A2.t11 VGND 0.0482f
C35654 _424_.A2.t10 VGND 0.04578f
C35655 _424_.A2.n6 VGND 0.06511f
C35656 _424_.A2.t15 VGND 0.02737f
C35657 _424_.A2.t9 VGND 0.03764f
C35658 _424_.A2.n7 VGND 0.05872f
C35659 _424_.A2.n8 VGND 0.5784f
C35660 _424_.A2.n9 VGND 0.37205f
C35661 _424_.A2.t14 VGND 0.0482f
C35662 _424_.A2.t8 VGND 0.04578f
C35663 _424_.A2.n10 VGND 0.06511f
C35664 _424_.A2.n11 VGND 0.62608f
C35665 _424_.A2.n12 VGND 0.89028f
C35666 _424_.A2.n13 VGND 0.10996f
C35667 _424_.A2.n14 VGND 0.05582f
C35668 _424_.A2.t2 VGND 0.0151f
C35669 _424_.A2.t1 VGND 0.0151f
C35670 _424_.A2.n15 VGND 0.03944f
C35671 a_45508_20936.t6 VGND 0.04128f
C35672 a_45508_20936.t7 VGND 0.13823f
C35673 a_45508_20936.t4 VGND 0.12194f
C35674 a_45508_20936.n0 VGND 0.15796f
C35675 a_45508_20936.n1 VGND 0.05384f
C35676 a_45508_20936.t1 VGND 0.04561f
C35677 a_45508_20936.n2 VGND 0.20374f
C35678 a_45508_20936.t3 VGND 0.01944f
C35679 a_45508_20936.t5 VGND 0.12223f
C35680 a_45508_20936.t2 VGND 0.38419f
C35681 a_45508_20936.n3 VGND 0.24674f
C35682 a_45508_20936.n4 VGND 0.56455f
C35683 a_45508_20936.t0 VGND 0.10024f
C35684 _416_.A1.t2 VGND 0.00751f
C35685 _416_.A1.t3 VGND 0.00751f
C35686 _416_.A1.n0 VGND 0.01681f
C35687 _416_.A1.t7 VGND 0.04636f
C35688 _416_.A1.t10 VGND 0.06292f
C35689 _416_.A1.n1 VGND 0.06786f
C35690 _416_.A1.n2 VGND 0.16431f
C35691 _416_.A1.t14 VGND 0.06202f
C35692 _416_.A1.t4 VGND 0.03679f
C35693 _416_.A1.n3 VGND 0.06481f
C35694 _416_.A1.n4 VGND 0.80633f
C35695 _416_.A1.t9 VGND 0.0413f
C35696 _416_.A1.t15 VGND 0.05509f
C35697 _416_.A1.n5 VGND 0.06788f
C35698 _416_.A1.n6 VGND 0.15592f
C35699 _416_.A1.t13 VGND 0.0413f
C35700 _416_.A1.t5 VGND 0.05509f
C35701 _416_.A1.n7 VGND 0.06838f
C35702 _416_.A1.n8 VGND 0.52746f
C35703 _416_.A1.t8 VGND 0.05374f
C35704 _416_.A1.t11 VGND 0.04459f
C35705 _416_.A1.n9 VGND 0.06832f
C35706 _416_.A1.t6 VGND 0.0413f
C35707 _416_.A1.t12 VGND 0.05509f
C35708 _416_.A1.n10 VGND 0.06788f
C35709 _416_.A1.n11 VGND 0.11023f
C35710 _416_.A1.n12 VGND 0.97994f
C35711 _416_.A1.n13 VGND 1.17191f
C35712 _416_.A1.n14 VGND 1.00523f
C35713 _416_.A1.n15 VGND 0.08473f
C35714 _416_.A1.t0 VGND 0.02644f
C35715 _416_.A1.t1 VGND 0.0191f
C35716 _416_.A1.n16 VGND 0.0478f
C35717 _330_.A1.t0 VGND 0.03068f
C35718 _330_.A1.t1 VGND 0.02216f
C35719 _330_.A1.n0 VGND 0.05424f
C35720 _330_.A1.t2 VGND 0.01489f
C35721 _330_.A1.t3 VGND 0.01489f
C35722 _330_.A1.n1 VGND 0.03162f
C35723 _330_.A1.t11 VGND 0.06391f
C35724 _330_.A1.t4 VGND 0.04771f
C35725 _330_.A1.n2 VGND 0.07952f
C35726 _330_.A1.t17 VGND 0.06391f
C35727 _330_.A1.t9 VGND 0.04771f
C35728 _330_.A1.n3 VGND 0.07895f
C35729 _330_.A1.n4 VGND 0.03156f
C35730 _330_.A1.t12 VGND 0.06391f
C35731 _330_.A1.t23 VGND 0.04771f
C35732 _330_.A1.n5 VGND 0.07895f
C35733 _330_.A1.n6 VGND 0.0766f
C35734 _330_.A1.t8 VGND 0.06391f
C35735 _330_.A1.t16 VGND 0.04771f
C35736 _330_.A1.n7 VGND 0.07952f
C35737 _330_.A1.n8 VGND 0.40498f
C35738 _330_.A1.t14 VGND 0.04287f
C35739 _330_.A1.t15 VGND 0.07194f
C35740 _330_.A1.n9 VGND 0.075f
C35741 _330_.A1.n10 VGND 0.93588f
C35742 _330_.A1.n11 VGND 0.4449f
C35743 _330_.A1.t22 VGND 0.06391f
C35744 _330_.A1.t21 VGND 0.04771f
C35745 _330_.A1.n12 VGND 0.07895f
C35746 _330_.A1.n13 VGND 0.03156f
C35747 _330_.A1.n14 VGND 0.41648f
C35748 _330_.A1.n15 VGND 0.40418f
C35749 _330_.A1.t5 VGND 0.06391f
C35750 _330_.A1.t20 VGND 0.04771f
C35751 _330_.A1.n16 VGND 0.07952f
C35752 _330_.A1.n17 VGND 0.75814f
C35753 _330_.A1.t13 VGND 0.04287f
C35754 _330_.A1.t7 VGND 0.07194f
C35755 _330_.A1.n18 VGND 0.0758f
C35756 _330_.A1.n19 VGND 0.03912f
C35757 _330_.A1.n20 VGND 1.29323f
C35758 _330_.A1.t10 VGND 0.06199f
C35759 _330_.A1.t6 VGND 0.06601f
C35760 _330_.A1.n21 VGND 0.07743f
C35761 _330_.A1.n22 VGND 0.98887f
C35762 _330_.A1.t18 VGND 0.06551f
C35763 _330_.A1.t19 VGND 0.06223f
C35764 _330_.A1.n23 VGND 0.0885f
C35765 _330_.A1.n24 VGND 0.80638f
C35766 _330_.A1.n25 VGND 0.09875f
C35767 a_39124_27208.t2 VGND 0.04128f
C35768 a_39124_27208.t5 VGND 0.13823f
C35769 a_39124_27208.t6 VGND 0.12194f
C35770 a_39124_27208.n0 VGND 0.15796f
C35771 a_39124_27208.n1 VGND 0.05384f
C35772 a_39124_27208.t1 VGND 0.04561f
C35773 a_39124_27208.n2 VGND 0.20374f
C35774 a_39124_27208.t3 VGND 0.01944f
C35775 a_39124_27208.t7 VGND 0.12223f
C35776 a_39124_27208.t4 VGND 0.38419f
C35777 a_39124_27208.n3 VGND 0.24674f
C35778 a_39124_27208.n4 VGND 0.56455f
C35779 a_39124_27208.t0 VGND 0.10024f
C35780 _325_.A1.t0 VGND 0.02f
C35781 _325_.A1.t1 VGND 0.02f
C35782 _325_.A1.n0 VGND 0.04039f
C35783 _325_.A1.t3 VGND 0.01344f
C35784 _325_.A1.t2 VGND 0.01344f
C35785 _325_.A1.n1 VGND 0.02707f
C35786 _325_.A1.t20 VGND 0.05595f
C35787 _325_.A1.t10 VGND 0.06077f
C35788 _325_.A1.n2 VGND 0.07026f
C35789 _325_.A1.n3 VGND 0.1068f
C35790 _325_.A1.t17 VGND 0.06299f
C35791 _325_.A1.t9 VGND 0.05125f
C35792 _325_.A1.n4 VGND 0.08082f
C35793 _325_.A1.t7 VGND 0.06077f
C35794 _325_.A1.t19 VGND 0.05579f
C35795 _325_.A1.n5 VGND 0.07077f
C35796 _325_.A1.n6 VGND 0.11237f
C35797 _325_.A1.n7 VGND 0.32997f
C35798 _325_.A1.n8 VGND 0.29099f
C35799 _325_.A1.t8 VGND 0.06273f
C35800 _325_.A1.t6 VGND 0.04879f
C35801 _325_.A1.n9 VGND 0.07072f
C35802 _325_.A1.n10 VGND 0.15599f
C35803 _325_.A1.t21 VGND 0.06014f
C35804 _325_.A1.t14 VGND 0.0524f
C35805 _325_.A1.n11 VGND 0.08226f
C35806 _325_.A1.n12 VGND 0.11274f
C35807 _325_.A1.t5 VGND 0.04325f
C35808 _325_.A1.t4 VGND 0.05973f
C35809 _325_.A1.n13 VGND 0.07589f
C35810 _325_.A1.n14 VGND 0.23458f
C35811 _325_.A1.t15 VGND 0.05973f
C35812 _325_.A1.t18 VGND 0.04325f
C35813 _325_.A1.n15 VGND 0.07546f
C35814 _325_.A1.n16 VGND 0.05024f
C35815 _325_.A1.n17 VGND 0.23418f
C35816 _325_.A1.t11 VGND 0.03394f
C35817 _325_.A1.t12 VGND 0.06241f
C35818 _325_.A1.n18 VGND 0.06478f
C35819 _325_.A1.n19 VGND 0.03611f
C35820 _325_.A1.n20 VGND 0.46141f
C35821 _325_.A1.t13 VGND 0.0357f
C35822 _325_.A1.t16 VGND 0.04555f
C35823 _325_.A1.n21 VGND 0.07486f
C35824 _325_.A1.n22 VGND 0.17174f
C35825 _325_.A1.n23 VGND 0.1588f
C35826 _325_.A1.n24 VGND 0.1036f
C35827 clk.t11 VGND 0.1054f
C35828 clk.t2 VGND 0.06956f
C35829 clk.t8 VGND 0.03867f
C35830 clk.n0 VGND 0.19171f
C35831 clk.t5 VGND 0.06956f
C35832 clk.t10 VGND 0.03867f
C35833 clk.n1 VGND 0.13541f
C35834 clk.t0 VGND 0.1007f
C35835 clk.t12 VGND 0.06956f
C35836 clk.t1 VGND 0.03867f
C35837 clk.n2 VGND 0.19042f
C35838 clk.t13 VGND 0.06956f
C35839 clk.t3 VGND 0.03867f
C35840 clk.n3 VGND 0.13541f
C35841 clk.t7 VGND 0.06956f
C35842 clk.t6 VGND 0.03867f
C35843 clk.n4 VGND 0.13541f
C35844 clk.t4 VGND 0.06956f
C35845 clk.t9 VGND 0.03867f
C35846 clk.n5 VGND 0.16087f
C35847 _455_.Q.t0 VGND 0.08744f
C35848 _455_.Q.t1 VGND 0.06164f
C35849 _455_.Q.t5 VGND 0.09616f
C35850 _455_.Q.t6 VGND 0.07388f
C35851 _455_.Q.n0 VGND 0.12718f
C35852 _455_.Q.n1 VGND 0.09114f
C35853 _455_.Q.t9 VGND 0.08722f
C35854 _455_.Q.t3 VGND 0.07388f
C35855 _455_.Q.n2 VGND 0.06281f
C35856 _455_.Q.n3 VGND 0.07408f
C35857 _455_.Q.t7 VGND 0.08722f
C35858 _455_.Q.n4 VGND 0.07408f
C35859 _455_.Q.t8 VGND 0.07388f
C35860 _455_.Q.n5 VGND 0.06281f
C35861 _455_.Q.n6 VGND 0.09893f
C35862 _455_.Q.t14 VGND 0.09621f
C35863 _455_.Q.t4 VGND 0.07388f
C35864 _455_.Q.n7 VGND 0.1167f
C35865 _455_.Q.n8 VGND 0.32375f
C35866 _455_.Q.t10 VGND 0.08543f
C35867 _455_.Q.t12 VGND 0.0928f
C35868 _455_.Q.n9 VGND 0.10783f
C35869 _455_.Q.n10 VGND 1.02485f
C35870 _455_.Q.t11 VGND 0.09618f
C35871 _455_.Q.t13 VGND 0.07826f
C35872 _455_.Q.n11 VGND 0.12354f
C35873 _455_.Q.t2 VGND 0.0928f
C35874 _455_.Q.t15 VGND 0.08519f
C35875 _455_.Q.n12 VGND 0.10807f
C35876 _455_.Q.n13 VGND 0.10709f
C35877 _455_.Q.n14 VGND 0.54005f
C35878 _455_.Q.n15 VGND 0.53498f
C35879 _437_.A1.t0 VGND 0.04194f
C35880 _437_.A1.t1 VGND 0.02957f
C35881 _437_.A1.t2 VGND 0.04482f
C35882 _437_.A1.t5 VGND 0.04075f
C35883 _437_.A1.n0 VGND 0.05131f
C35884 _437_.A1.t15 VGND 0.03229f
C35885 _437_.A1.t10 VGND 0.03371f
C35886 _437_.A1.n1 VGND 0.06197f
C35887 _437_.A1.n2 VGND 0.06819f
C35888 _437_.A1.t14 VGND 0.04756f
C35889 _437_.A1.t6 VGND 0.02822f
C35890 _437_.A1.n3 VGND 0.05024f
C35891 _437_.A1.n4 VGND 0.03025f
C35892 _437_.A1.t4 VGND 0.03382f
C35893 _437_.A1.t7 VGND 0.02448f
C35894 _437_.A1.n5 VGND 0.05289f
C35895 _437_.A1.n6 VGND 0.06809f
C35896 _437_.A1.t13 VGND 0.03168f
C35897 _437_.A1.t12 VGND 0.04375f
C35898 _437_.A1.n7 VGND 0.05527f
C35899 _437_.A1.n8 VGND 0.0184f
C35900 _437_.A1.n9 VGND 0.24275f
C35901 _437_.A1.t9 VGND 0.04756f
C35902 _437_.A1.t3 VGND 0.02822f
C35903 _437_.A1.n10 VGND 0.05024f
C35904 _437_.A1.n11 VGND 0.11441f
C35905 _437_.A1.n12 VGND 0.33228f
C35906 _437_.A1.n13 VGND 0.34656f
C35907 _437_.A1.t8 VGND 0.02834f
C35908 _437_.A1.t11 VGND 0.04756f
C35909 _437_.A1.n14 VGND 0.04958f
C35910 _437_.A1.n15 VGND 0.24755f
C35911 _437_.A1.n16 VGND 0.18218f
C35912 a_27588_29159.t2 VGND 0.12779f
C35913 a_27588_29159.t4 VGND 0.40165f
C35914 a_27588_29159.t5 VGND 0.02032f
C35915 a_27588_29159.n0 VGND 0.25796f
C35916 a_27588_29159.t7 VGND 0.14451f
C35917 a_27588_29159.t6 VGND 0.12788f
C35918 a_27588_29159.n1 VGND 0.16475f
C35919 a_27588_29159.t3 VGND 0.04268f
C35920 a_27588_29159.n2 VGND 0.05675f
C35921 a_27588_29159.t1 VGND 0.04768f
C35922 a_27588_29159.n3 VGND 0.21301f
C35923 a_27588_29159.n4 VGND 0.59021f
C35924 a_27588_29159.t0 VGND 0.1048f
C35925 _229_.I.t0 VGND 0.06688f
C35926 _229_.I.t1 VGND 0.04508f
C35927 _229_.I.t14 VGND 0.06672f
C35928 _229_.I.t2 VGND 0.06435f
C35929 _229_.I.n0 VGND 0.08154f
C35930 _229_.I.t10 VGND 0.05676f
C35931 _229_.I.t7 VGND 0.04136f
C35932 _229_.I.n1 VGND 0.09327f
C35933 _229_.I.t9 VGND 0.06502f
C35934 _229_.I.t8 VGND 0.07247f
C35935 _229_.I.n2 VGND 0.08798f
C35936 _229_.I.n3 VGND 0.06207f
C35937 _229_.I.t5 VGND 0.07125f
C35938 _229_.I.t4 VGND 0.06653f
C35939 _229_.I.n4 VGND 0.08338f
C35940 _229_.I.n5 VGND 0.01147f
C35941 _229_.I.t15 VGND 0.04047f
C35942 _229_.I.t3 VGND 0.07442f
C35943 _229_.I.n6 VGND 0.07753f
C35944 _229_.I.t12 VGND 0.05818f
C35945 _229_.I.t13 VGND 0.0748f
C35946 _229_.I.n7 VGND 0.08433f
C35947 _229_.I.n8 VGND 0.4003f
C35948 _229_.I.t6 VGND 0.06797f
C35949 _229_.I.t11 VGND 0.04567f
C35950 _229_.I.n9 VGND 0.10443f
C35951 _229_.I.n10 VGND 0.21044f
C35952 _229_.I.n11 VGND 0.44527f
C35953 _229_.I.n12 VGND 0.22244f
C35954 _229_.I.n13 VGND 0.16356f
C35955 _229_.I.n14 VGND 0.28927f
C35956 _229_.I.n15 VGND 0.20981f
C35957 _448_.Q.t1 VGND 0.04844f
C35958 _448_.Q.t0 VGND 0.06872f
C35959 _448_.Q.t5 VGND 0.07792f
C35960 _448_.Q.t2 VGND 0.04623f
C35961 _448_.Q.n0 VGND 0.08143f
C35962 _448_.Q.t4 VGND 0.05693f
C35963 _448_.Q.t9 VGND 0.07643f
C35964 _448_.Q.n1 VGND 0.09111f
C35965 _448_.Q.t8 VGND 0.07206f
C35966 _448_.Q.t7 VGND 0.06232f
C35967 _448_.Q.n2 VGND 0.0846f
C35968 _448_.Q.t12 VGND 0.07217f
C35969 _448_.Q.t14 VGND 0.06288f
C35970 _448_.Q.n3 VGND 0.09875f
C35971 _448_.Q.n4 VGND 0.80077f
C35972 _448_.Q.t11 VGND 0.07981f
C35973 _448_.Q.t10 VGND 0.04979f
C35974 _448_.Q.n5 VGND 0.09478f
C35975 _448_.Q.n6 VGND 0.09398f
C35976 _448_.Q.n7 VGND 0.51145f
C35977 _448_.Q.n8 VGND 0.30289f
C35978 _448_.Q.t6 VGND 0.07489f
C35979 _448_.Q.t15 VGND 0.04073f
C35980 _448_.Q.n9 VGND 0.07802f
C35981 _448_.Q.n10 VGND 0.18206f
C35982 _448_.Q.t3 VGND 0.05541f
C35983 _448_.Q.t13 VGND 0.0401f
C35984 _448_.Q.n11 VGND 0.08665f
C35985 _448_.Q.n12 VGND 0.20671f
C35986 _448_.Q.n13 VGND 0.33329f
C35987 a_17060_28776.t6 VGND 0.04104f
C35988 a_17060_28776.t2 VGND 0.13745f
C35989 a_17060_28776.t4 VGND 0.12126f
C35990 a_17060_28776.n0 VGND 0.15708f
C35991 a_17060_28776.n1 VGND 0.05354f
C35992 a_17060_28776.t1 VGND 0.04536f
C35993 a_17060_28776.n2 VGND 0.19884f
C35994 a_17060_28776.t7 VGND 0.01933f
C35995 a_17060_28776.t3 VGND 0.12155f
C35996 a_17060_28776.t5 VGND 0.38204f
C35997 a_17060_28776.n3 VGND 0.24693f
C35998 a_17060_28776.n4 VGND 0.58092f
C35999 a_17060_28776.t0 VGND 0.09466f
C36000 a_42392_22825.t4 VGND 0.05796f
C36001 a_42392_22825.t3 VGND 0.04186f
C36002 a_42392_22825.t5 VGND 0.05796f
C36003 a_42392_22825.n0 VGND 0.12446f
C36004 a_42392_22825.t6 VGND 0.04186f
C36005 a_42392_22825.t1 VGND 0.05796f
C36006 a_42392_22825.n1 VGND 0.10102f
C36007 a_42392_22825.t0 VGND 0.04186f
C36008 a_42392_22825.t2 VGND 0.05796f
C36009 a_42392_22825.n2 VGND 0.10102f
C36010 a_42392_22825.t12 VGND 0.05137f
C36011 a_42392_22825.t11 VGND 0.02067f
C36012 a_42392_22825.t13 VGND 0.02067f
C36013 a_42392_22825.n3 VGND 0.04203f
C36014 a_42392_22825.t10 VGND 0.02067f
C36015 a_42392_22825.t8 VGND 0.02067f
C36016 a_42392_22825.n4 VGND 0.04203f
C36017 a_42392_22825.t9 VGND 0.06511f
C36018 a_42392_22825.n5 VGND 0.41377f
C36019 a_42392_22825.n6 VGND 0.2495f
C36020 a_42392_22825.n7 VGND 0.2072f
C36021 a_42392_22825.t32 VGND 0.18155f
C36022 a_42392_22825.t37 VGND 0.11957f
C36023 a_42392_22825.n8 VGND 0.26772f
C36024 a_42392_22825.t34 VGND 0.18155f
C36025 a_42392_22825.t40 VGND 0.11957f
C36026 a_42392_22825.n9 VGND 0.30447f
C36027 a_42392_22825.t30 VGND 0.18155f
C36028 a_42392_22825.t36 VGND 0.11957f
C36029 a_42392_22825.n10 VGND 0.30447f
C36030 a_42392_22825.t20 VGND 0.18155f
C36031 a_42392_22825.t22 VGND 0.18155f
C36032 a_42392_22825.t17 VGND 0.11957f
C36033 a_42392_22825.n11 VGND 0.26772f
C36034 a_42392_22825.t28 VGND 0.18155f
C36035 a_42392_22825.t33 VGND 0.11957f
C36036 a_42392_22825.n12 VGND 0.30447f
C36037 a_42392_22825.t23 VGND 0.18155f
C36038 a_42392_22825.t29 VGND 0.11957f
C36039 a_42392_22825.n13 VGND 0.30447f
C36040 a_42392_22825.t24 VGND 0.18155f
C36041 a_42392_22825.t31 VGND 0.11957f
C36042 a_42392_22825.n14 VGND -0.56964f
C36043 a_42392_22825.t41 VGND 0.18155f
C36044 a_42392_22825.t35 VGND 0.11957f
C36045 a_42392_22825.n15 VGND 0.30447f
C36046 a_42392_22825.t38 VGND 0.18155f
C36047 a_42392_22825.t43 VGND 0.11957f
C36048 a_42392_22825.n16 VGND 0.30447f
C36049 a_42392_22825.t42 VGND 0.18155f
C36050 a_42392_22825.t14 VGND 0.11957f
C36051 a_42392_22825.n17 VGND 0.30447f
C36052 a_42392_22825.t39 VGND 0.18155f
C36053 a_42392_22825.t44 VGND 0.11957f
C36054 a_42392_22825.n18 VGND 0.30447f
C36055 a_42392_22825.t15 VGND 0.18155f
C36056 a_42392_22825.t45 VGND 0.11957f
C36057 a_42392_22825.n19 VGND 0.30447f
C36058 a_42392_22825.t19 VGND 0.18155f
C36059 a_42392_22825.t26 VGND 0.11957f
C36060 a_42392_22825.n20 VGND 0.30447f
C36061 a_42392_22825.t16 VGND 0.18155f
C36062 a_42392_22825.n21 VGND 0.15345f
C36063 a_42392_22825.t21 VGND 0.11898f
C36064 a_42392_22825.n22 VGND 0.15264f
C36065 a_42392_22825.t27 VGND 0.11898f
C36066 a_42392_22825.n23 VGND 0.15264f
C36067 a_42392_22825.n24 VGND 0.15345f
C36068 a_42392_22825.t25 VGND 0.18155f
C36069 a_42392_22825.t18 VGND 0.11957f
C36070 a_42392_22825.n25 VGND 0.83236f
C36071 a_42392_22825.n26 VGND 0.57691f
C36072 a_42392_22825.n27 VGND 0.21092f
C36073 a_42392_22825.n28 VGND 0.25801f
C36074 a_42392_22825.n29 VGND 0.40181f
C36075 a_42392_22825.n30 VGND 0.10102f
C36076 a_42392_22825.t7 VGND 0.04186f
C36077 a_36996_18183.t3 VGND 0.12779f
C36078 a_36996_18183.t4 VGND 0.40165f
C36079 a_36996_18183.t5 VGND 0.02032f
C36080 a_36996_18183.n0 VGND 0.25796f
C36081 a_36996_18183.t2 VGND 0.14451f
C36082 a_36996_18183.t7 VGND 0.12788f
C36083 a_36996_18183.n1 VGND 0.16475f
C36084 a_36996_18183.t6 VGND 0.04268f
C36085 a_36996_18183.n2 VGND 0.05675f
C36086 a_36996_18183.t1 VGND 0.04768f
C36087 a_36996_18183.n3 VGND 0.21301f
C36088 a_36996_18183.n4 VGND 0.59021f
C36089 a_36996_18183.t0 VGND 0.1048f
C36090 a_49152_30301.t1 VGND 0.04561f
C36091 a_49152_30301.t4 VGND 0.04128f
C36092 a_49152_30301.t6 VGND 0.13823f
C36093 a_49152_30301.t7 VGND 0.12194f
C36094 a_49152_30301.n0 VGND 0.15796f
C36095 a_49152_30301.n1 VGND 0.05384f
C36096 a_49152_30301.n2 VGND 0.20374f
C36097 a_49152_30301.t5 VGND 0.01944f
C36098 a_49152_30301.t3 VGND 0.12223f
C36099 a_49152_30301.t2 VGND 0.38419f
C36100 a_49152_30301.n3 VGND 0.24674f
C36101 a_49152_30301.n4 VGND 0.56455f
C36102 a_49152_30301.t0 VGND 0.10024f
C36103 _452_.Q.t4 VGND 0.05557f
C36104 _452_.Q.t18 VGND 0.07113f
C36105 _452_.Q.n0 VGND 0.11108f
C36106 _452_.Q.t14 VGND 0.09135f
C36107 _452_.Q.t7 VGND 0.04513f
C36108 _452_.Q.n1 VGND 0.13704f
C36109 _452_.Q.n2 VGND 0.06383f
C36110 _452_.Q.t16 VGND 0.06937f
C36111 _452_.Q.t10 VGND 0.08171f
C36112 _452_.Q.n3 VGND 0.1144f
C36113 _452_.Q.t20 VGND 0.07692f
C36114 _452_.Q.t5 VGND 0.07636f
C36115 _452_.Q.n4 VGND 0.1122f
C36116 _452_.Q.n5 VGND 0.24041f
C36117 _452_.Q.n6 VGND 0.4149f
C36118 _452_.Q.n7 VGND 0.47593f
C36119 _452_.Q.t13 VGND 0.06527f
C36120 _452_.Q.t9 VGND 0.08706f
C36121 _452_.Q.n8 VGND 0.10896f
C36122 _452_.Q.n9 VGND 0.30339f
C36123 _452_.Q.t6 VGND 0.0854f
C36124 _452_.Q.t8 VGND 0.08085f
C36125 _452_.Q.n10 VGND 0.11626f
C36126 _452_.Q.t12 VGND 0.09016f
C36127 _452_.Q.t17 VGND 0.06528f
C36128 _452_.Q.n11 VGND 0.11389f
C36129 _452_.Q.n12 VGND 0.03586f
C36130 _452_.Q.n13 VGND 0.80282f
C36131 _452_.Q.n14 VGND 0.4837f
C36132 _452_.Q.t19 VGND 0.08297f
C36133 _452_.Q.t15 VGND 0.08445f
C36134 _452_.Q.n15 VGND 0.1153f
C36135 _452_.Q.n16 VGND 0.80949f
C36136 _452_.Q.t11 VGND 0.06899f
C36137 _452_.Q.t21 VGND 0.05389f
C36138 _452_.Q.n17 VGND 0.11272f
C36139 _452_.Q.n18 VGND 0.49104f
C36140 _452_.Q.t0 VGND 0.03018f
C36141 _452_.Q.t1 VGND 0.03018f
C36142 _452_.Q.n19 VGND 0.06036f
C36143 _452_.Q.n20 VGND 0.04473f
C36144 _452_.Q.t2 VGND 0.02029f
C36145 _452_.Q.t3 VGND 0.02029f
C36146 _452_.Q.n21 VGND 0.04857f
C36147 _459_.Q.t0 VGND 0.05876f
C36148 _459_.Q.t1 VGND 0.04142f
C36149 _459_.Q.t14 VGND 0.04258f
C36150 _459_.Q.n0 VGND 0.04016f
C36151 _459_.Q.t8 VGND 0.04258f
C36152 _459_.Q.t3 VGND 0.05515f
C36153 _459_.Q.n1 VGND 0.06337f
C36154 _459_.Q.t12 VGND 0.05515f
C36155 _459_.Q.n2 VGND 0.06337f
C36156 _459_.Q.n3 VGND 0.03916f
C36157 _459_.Q.n4 VGND 0.06561f
C36158 _459_.Q.t13 VGND 0.04258f
C36159 _459_.Q.n5 VGND 0.04009f
C36160 _459_.Q.t9 VGND 0.04258f
C36161 _459_.Q.t17 VGND 0.05515f
C36162 _459_.Q.t15 VGND 0.05515f
C36163 _459_.Q.n6 VGND 0.06337f
C36164 _459_.Q.n7 VGND 0.06337f
C36165 _459_.Q.n8 VGND 0.03916f
C36166 _459_.Q.n9 VGND 0.04456f
C36167 _459_.Q.n10 VGND 0.48307f
C36168 _459_.Q.t16 VGND 0.05122f
C36169 _459_.Q.t10 VGND 0.05887f
C36170 _459_.Q.n11 VGND 0.07257f
C36171 _459_.Q.t11 VGND 0.06663f
C36172 _459_.Q.t5 VGND 0.03953f
C36173 _459_.Q.n12 VGND 0.06963f
C36174 _459_.Q.n13 VGND 0.58004f
C36175 _459_.Q.t6 VGND 0.05758f
C36176 _459_.Q.t4 VGND 0.05641f
C36177 _459_.Q.n14 VGND 0.07823f
C36178 _459_.Q.t7 VGND 0.0469f
C36179 _459_.Q.t2 VGND 0.03664f
C36180 _459_.Q.n15 VGND 0.07665f
C36181 _459_.Q.n16 VGND 0.46095f
C36182 _459_.Q.n17 VGND 0.95368f
C36183 _352_.A2.t3 VGND 0.02494f
C36184 _352_.A2.t9 VGND 0.02494f
C36185 _352_.A2.n0 VGND 0.05604f
C36186 _352_.A2.t11 VGND 0.02494f
C36187 _352_.A2.t0 VGND 0.02494f
C36188 _352_.A2.n1 VGND 0.04989f
C36189 _352_.A2.n2 VGND 0.19268f
C36190 _352_.A2.t2 VGND 0.02494f
C36191 _352_.A2.t10 VGND 0.02494f
C36192 _352_.A2.n3 VGND 0.04989f
C36193 _352_.A2.n4 VGND 0.12127f
C36194 _352_.A2.t14 VGND 0.01704f
C36195 _352_.A2.t13 VGND 0.01704f
C36196 _352_.A2.n5 VGND 0.05075f
C36197 _352_.A2.t12 VGND 0.01704f
C36198 _352_.A2.t15 VGND 0.01704f
C36199 _352_.A2.n6 VGND 0.03409f
C36200 _352_.A2.n7 VGND 0.19058f
C36201 _352_.A2.t5 VGND 0.0106f
C36202 _352_.A2.t6 VGND 0.0106f
C36203 _352_.A2.n8 VGND 0.02148f
C36204 _352_.A2.t24 VGND 0.07395f
C36205 _352_.A2.t27 VGND 0.06462f
C36206 _352_.A2.n9 VGND 0.08656f
C36207 _352_.A2.n10 VGND 0.09185f
C36208 _352_.A2.t26 VGND 0.07315f
C36209 _352_.A2.t29 VGND 0.05461f
C36210 _352_.A2.n11 VGND 0.09033f
C36211 _352_.A2.n12 VGND 0.25389f
C36212 _352_.A2.t28 VGND 0.05556f
C36213 _352_.A2.t16 VGND 0.04992f
C36214 _352_.A2.n13 VGND 0.10123f
C36215 _352_.A2.t22 VGND 0.08254f
C36216 _352_.A2.t25 VGND 0.06187f
C36217 _352_.A2.n14 VGND 0.10117f
C36218 _352_.A2.n15 VGND 0.18655f
C36219 _352_.A2.n16 VGND 0.66952f
C36220 _352_.A2.n17 VGND 0.38502f
C36221 _352_.A2.t20 VGND 0.08034f
C36222 _352_.A2.t23 VGND 0.0205f
C36223 _352_.A2.n18 VGND 0.1015f
C36224 _352_.A2.t19 VGND 0.07095f
C36225 _352_.A2.t31 VGND 0.07707f
C36226 _352_.A2.n19 VGND 0.0891f
C36227 _352_.A2.n20 VGND 0.03788f
C36228 _352_.A2.t17 VGND 0.05415f
C36229 _352_.A2.t30 VGND 0.08354f
C36230 _352_.A2.n21 VGND 0.08662f
C36231 _352_.A2.n22 VGND 0.42533f
C36232 _352_.A2.n23 VGND 0.54196f
C36233 _352_.A2.n24 VGND 0.32802f
C36234 _352_.A2.t21 VGND 0.07707f
C36235 _352_.A2.t18 VGND 0.07075f
C36236 _352_.A2.n25 VGND 0.0893f
C36237 _352_.A2.n26 VGND 0.22536f
C36238 _352_.A2.t4 VGND 0.0106f
C36239 _352_.A2.t7 VGND 0.0106f
C36240 _352_.A2.n27 VGND 0.0212f
C36241 _352_.A2.n28 VGND 0.09486f
C36242 _352_.A2.n29 VGND 0.112f
C36243 _352_.A2.n30 VGND 0.12525f
C36244 _352_.A2.t8 VGND 0.02494f
C36245 _352_.A2.t1 VGND 0.02494f
C36246 _352_.A2.n31 VGND 0.04989f
C36247 _352_.A2.n32 VGND 0.06649f
C36248 _381_.A2.t4 VGND 0.03949f
C36249 _381_.A2.t7 VGND 0.04244f
C36250 _381_.A2.n0 VGND 0.07387f
C36251 _381_.A2.t3 VGND 0.04355f
C36252 _381_.A2.t2 VGND 0.05591f
C36253 _381_.A2.n1 VGND 0.06975f
C36254 _381_.A2.t5 VGND 0.04659f
C36255 _381_.A2.t6 VGND 0.05161f
C36256 _381_.A2.n2 VGND 0.08294f
C36257 _381_.A2.n3 VGND 0.09277f
C36258 _381_.A2.n4 VGND 0.71082f
C36259 _381_.A2.t1 VGND 0.03243f
C36260 _381_.A2.n5 VGND 0.19231f
C36261 _381_.A2.t0 VGND 0.04403f
C36262 _335_.ZN.t2 VGND 0.024f
C36263 _335_.ZN.t15 VGND 0.024f
C36264 _335_.ZN.n0 VGND 0.04868f
C36265 _335_.ZN.t13 VGND 0.024f
C36266 _335_.ZN.t1 VGND 0.024f
C36267 _335_.ZN.n1 VGND 0.04868f
C36268 _335_.ZN.t4 VGND 0.04299f
C36269 _335_.ZN.t7 VGND 0.04299f
C36270 _335_.ZN.n2 VGND 0.10302f
C36271 _335_.ZN.t6 VGND 0.04299f
C36272 _335_.ZN.t5 VGND 0.04299f
C36273 _335_.ZN.n3 VGND 0.07615f
C36274 _335_.ZN.n4 VGND 0.3294f
C36275 _335_.ZN.n5 VGND 0.25354f
C36276 _335_.ZN.n6 VGND 0.16799f
C36277 _335_.ZN.t12 VGND 0.024f
C36278 _335_.ZN.t3 VGND 0.024f
C36279 _335_.ZN.n7 VGND 0.04868f
C36280 _335_.ZN.n8 VGND 0.16018f
C36281 _335_.ZN.t0 VGND 0.024f
C36282 _335_.ZN.t14 VGND 0.024f
C36283 _335_.ZN.n9 VGND 0.04868f
C36284 _335_.ZN.t9 VGND 0.024f
C36285 _335_.ZN.t16 VGND 0.024f
C36286 _335_.ZN.n10 VGND 0.04868f
C36287 _335_.ZN.t17 VGND 0.024f
C36288 _335_.ZN.t11 VGND 0.024f
C36289 _335_.ZN.n11 VGND 0.04868f
C36290 _335_.ZN.t10 VGND 0.024f
C36291 _335_.ZN.t19 VGND 0.024f
C36292 _335_.ZN.n12 VGND 0.04868f
C36293 _335_.ZN.t18 VGND 0.024f
C36294 _335_.ZN.t8 VGND 0.024f
C36295 _335_.ZN.n13 VGND 0.04873f
C36296 _335_.ZN.t20 VGND 0.07012f
C36297 _335_.ZN.t23 VGND 0.11788f
C36298 _335_.ZN.n14 VGND 0.15816f
C36299 _335_.ZN.t25 VGND 0.10354f
C36300 _335_.ZN.t26 VGND 0.09129f
C36301 _335_.ZN.n15 VGND 0.15892f
C36302 _335_.ZN.n16 VGND 0.04903f
C36303 _335_.ZN.t27 VGND 0.07012f
C36304 _335_.ZN.t24 VGND 0.09539f
C36305 _335_.ZN.t21 VGND 0.07012f
C36306 _335_.ZN.n17 VGND 0.07307f
C36307 _335_.ZN.t22 VGND 0.09539f
C36308 _335_.ZN.n18 VGND 0.115f
C36309 _335_.ZN.n19 VGND 0.115f
C36310 _335_.ZN.n20 VGND 0.07307f
C36311 _335_.ZN.n21 VGND 0.05342f
C36312 _335_.ZN.n22 VGND 0.39608f
C36313 _335_.ZN.n23 VGND 0.31271f
C36314 _335_.ZN.n24 VGND 0.15417f
C36315 _335_.ZN.n25 VGND 0.15477f
C36316 _335_.ZN.n26 VGND 0.15477f
C36317 _335_.ZN.n27 VGND 0.1013f
C36318 uo_out[1].t1 VGND 0.03335f
C36319 uo_out[1].t0 VGND 0.03335f
C36320 uo_out[1].n0 VGND 0.06745f
C36321 uo_out[1].t11 VGND 0.01115f
C36322 uo_out[1].t5 VGND 0.01115f
C36323 uo_out[1].n1 VGND 0.0224f
C36324 uo_out[1].t2 VGND 0.01115f
C36325 uo_out[1].t9 VGND 0.01115f
C36326 uo_out[1].n2 VGND 0.0224f
C36327 uo_out[1].t10 VGND 0.01115f
C36328 uo_out[1].t3 VGND 0.01115f
C36329 uo_out[1].n3 VGND 0.0224f
C36330 uo_out[1].t4 VGND 0.01115f
C36331 uo_out[1].t8 VGND 0.01115f
C36332 uo_out[1].n4 VGND 0.02919f
C36333 uo_out[1].n5 VGND 0.14113f
C36334 uo_out[1].n6 VGND 0.08985f
C36335 uo_out[1].n7 VGND 0.146f
C36336 uo_out[1].n8 VGND 0.17283f
C36337 uo_out[1].t6 VGND 0.03335f
C36338 uo_out[1].t7 VGND 0.03335f
C36339 uo_out[1].n9 VGND 0.0667f
C36340 uo_out[1].n10 VGND 0.36414f
C36341 a_20084_26023.t3 VGND 0.12223f
C36342 a_20084_26023.t6 VGND 0.38419f
C36343 a_20084_26023.t5 VGND 0.01944f
C36344 a_20084_26023.n0 VGND 0.24674f
C36345 a_20084_26023.t2 VGND 0.13823f
C36346 a_20084_26023.t7 VGND 0.12232f
C36347 a_20084_26023.n1 VGND 0.15759f
C36348 a_20084_26023.t4 VGND 0.04083f
C36349 a_20084_26023.n2 VGND 0.05429f
C36350 a_20084_26023.t1 VGND 0.04561f
C36351 a_20084_26023.n3 VGND 0.20374f
C36352 a_20084_26023.n4 VGND 0.56455f
C36353 a_20084_26023.t0 VGND 0.10024f
C36354 _251_.A1.t1 VGND 0.02244f
C36355 _251_.A1.t0 VGND 0.01621f
C36356 _251_.A1.n0 VGND 0.03905f
C36357 _251_.A1.t5 VGND 0.00604f
C36358 _251_.A1.t4 VGND 0.00604f
C36359 _251_.A1.n1 VGND 0.01231f
C36360 _251_.A1.t6 VGND 0.00604f
C36361 _251_.A1.t7 VGND 0.00604f
C36362 _251_.A1.n2 VGND 0.01741f
C36363 _251_.A1.n3 VGND 0.10478f
C36364 _251_.A1.n4 VGND 0.05772f
C36365 _251_.A1.t2 VGND 0.01621f
C36366 _251_.A1.t3 VGND 0.02244f
C36367 _251_.A1.n5 VGND 0.03943f
C36368 _251_.A1.t24 VGND 0.02751f
C36369 _251_.A1.t18 VGND 0.05058f
C36370 _251_.A1.n6 VGND 0.05269f
C36371 _251_.A1.t30 VGND 0.05262f
C36372 _251_.A1.t25 VGND 0.03122f
C36373 _251_.A1.n7 VGND 0.05499f
C36374 _251_.A1.t23 VGND 0.04991f
C36375 _251_.A1.t9 VGND 0.04445f
C36376 _251_.A1.t16 VGND 0.05118f
C36377 _251_.A1.n8 VGND 0.06055f
C36378 _251_.A1.t15 VGND 0.05483f
C36379 _251_.A1.n9 VGND 0.09479f
C36380 _251_.A1.n10 VGND 0.09027f
C36381 _251_.A1.t20 VGND 0.05021f
C36382 _251_.A1.t19 VGND 0.05118f
C36383 _251_.A1.t33 VGND 0.04445f
C36384 _251_.A1.n11 VGND 0.06055f
C36385 _251_.A1.t29 VGND 0.05483f
C36386 _251_.A1.n12 VGND 0.09479f
C36387 _251_.A1.n13 VGND 0.07162f
C36388 _251_.A1.n14 VGND 0.37932f
C36389 _251_.A1.n15 VGND 0.45394f
C36390 _251_.A1.n16 VGND 0.33026f
C36391 _251_.A1.t13 VGND 0.03136f
C36392 _251_.A1.t14 VGND 0.05262f
C36393 _251_.A1.n17 VGND 0.05486f
C36394 _251_.A1.t22 VGND 0.05352f
C36395 _251_.A1.t34 VGND 0.03461f
C36396 _251_.A1.n18 VGND 0.05509f
C36397 _251_.A1.n19 VGND 0.06792f
C36398 _251_.A1.n20 VGND 0.17404f
C36399 _251_.A1.t11 VGND 0.05021f
C36400 _251_.A1.t32 VGND 0.05118f
C36401 _251_.A1.t27 VGND 0.04445f
C36402 _251_.A1.n21 VGND 0.06055f
C36403 _251_.A1.t10 VGND 0.05483f
C36404 _251_.A1.n22 VGND 0.09479f
C36405 _251_.A1.n23 VGND 0.07905f
C36406 _251_.A1.n24 VGND 0.3101f
C36407 _251_.A1.t28 VGND 0.05118f
C36408 _251_.A1.t35 VGND 0.04445f
C36409 _251_.A1.n25 VGND 0.06055f
C36410 _251_.A1.t31 VGND 0.05483f
C36411 _251_.A1.n26 VGND 0.09479f
C36412 _251_.A1.t26 VGND 0.05021f
C36413 _251_.A1.n27 VGND 0.07162f
C36414 _251_.A1.n28 VGND 0.31302f
C36415 _251_.A1.t8 VGND 0.03461f
C36416 _251_.A1.t12 VGND 0.05339f
C36417 _251_.A1.n29 VGND 0.05522f
C36418 _251_.A1.n30 VGND 0.02261f
C36419 _251_.A1.n31 VGND 0.3412f
C36420 _251_.A1.n32 VGND 0.56858f
C36421 _251_.A1.t21 VGND 0.04534f
C36422 _251_.A1.t17 VGND 0.03523f
C36423 _251_.A1.n33 VGND 0.05541f
C36424 _251_.A1.n34 VGND 0.24563f
C36425 _251_.A1.n35 VGND 0.09824f
C36426 a_23668_25640.t2 VGND 0.04128f
C36427 a_23668_25640.t5 VGND 0.13823f
C36428 a_23668_25640.t3 VGND 0.12194f
C36429 a_23668_25640.n0 VGND 0.15796f
C36430 a_23668_25640.n1 VGND 0.05384f
C36431 a_23668_25640.t1 VGND 0.04561f
C36432 a_23668_25640.n2 VGND 0.20374f
C36433 a_23668_25640.t4 VGND 0.01944f
C36434 a_23668_25640.t6 VGND 0.12223f
C36435 a_23668_25640.t7 VGND 0.38419f
C36436 a_23668_25640.n3 VGND 0.24674f
C36437 a_23668_25640.n4 VGND 0.56455f
C36438 a_23668_25640.t0 VGND 0.10024f
C36439 a_45284_19751.t6 VGND 0.12223f
C36440 a_45284_19751.t7 VGND 0.38419f
C36441 a_45284_19751.t3 VGND 0.01944f
C36442 a_45284_19751.n0 VGND 0.24674f
C36443 a_45284_19751.t5 VGND 0.13823f
C36444 a_45284_19751.t4 VGND 0.12232f
C36445 a_45284_19751.n1 VGND 0.15759f
C36446 a_45284_19751.t2 VGND 0.04083f
C36447 a_45284_19751.n2 VGND 0.05429f
C36448 a_45284_19751.t1 VGND 0.04561f
C36449 a_45284_19751.n3 VGND 0.20374f
C36450 a_45284_19751.n4 VGND 0.56455f
C36451 a_45284_19751.t0 VGND 0.10024f
C36452 _459_.CLK.t9 VGND 0.00961f
C36453 _459_.CLK.t10 VGND 0.00961f
C36454 _459_.CLK.n0 VGND 0.01953f
C36455 _459_.CLK.t12 VGND 0.00961f
C36456 _459_.CLK.t11 VGND 0.00961f
C36457 _459_.CLK.n1 VGND 0.02754f
C36458 _459_.CLK.n2 VGND 0.16648f
C36459 _459_.CLK.t14 VGND 0.00961f
C36460 _459_.CLK.t15 VGND 0.00961f
C36461 _459_.CLK.n3 VGND 0.01953f
C36462 _459_.CLK.t13 VGND 0.00961f
C36463 _459_.CLK.t8 VGND 0.00961f
C36464 _459_.CLK.n4 VGND 0.02754f
C36465 _459_.CLK.n5 VGND 0.18144f
C36466 _459_.CLK.n6 VGND 0.0753f
C36467 _459_.CLK.t5 VGND 0.03777f
C36468 _459_.CLK.t2 VGND 0.03777f
C36469 _459_.CLK.n7 VGND 0.07648f
C36470 _459_.CLK.t6 VGND 0.03777f
C36471 _459_.CLK.t3 VGND 0.03777f
C36472 _459_.CLK.n8 VGND 0.07755f
C36473 _459_.CLK.t47 VGND 0.05003f
C36474 _459_.CLK.t51 VGND 0.05332f
C36475 _459_.CLK.n9 VGND 0.07887f
C36476 _459_.CLK.t44 VGND 0.05353f
C36477 _459_.CLK.t25 VGND 0.04981f
C36478 _459_.CLK.n10 VGND 0.07888f
C36479 _459_.CLK.t49 VGND 0.04179f
C36480 _459_.CLK.t50 VGND 0.06541f
C36481 _459_.CLK.n11 VGND 0.11319f
C36482 _459_.CLK.n12 VGND 0.26581f
C36483 _459_.CLK.t19 VGND 0.05003f
C36484 _459_.CLK.t33 VGND 0.05332f
C36485 _459_.CLK.n13 VGND 0.07878f
C36486 _459_.CLK.n14 VGND 0.04632f
C36487 _459_.CLK.n15 VGND 0.39794f
C36488 _459_.CLK.t23 VGND 0.05003f
C36489 _459_.CLK.t37 VGND 0.05332f
C36490 _459_.CLK.n16 VGND 0.07878f
C36491 _459_.CLK.n17 VGND 0.04632f
C36492 _459_.CLK.t24 VGND 0.05003f
C36493 _459_.CLK.t16 VGND 0.05332f
C36494 _459_.CLK.n18 VGND 0.07878f
C36495 _459_.CLK.n19 VGND 0.13118f
C36496 _459_.CLK.n20 VGND 0.45258f
C36497 _459_.CLK.t31 VGND 0.05353f
C36498 _459_.CLK.t29 VGND 0.04981f
C36499 _459_.CLK.n21 VGND 0.07879f
C36500 _459_.CLK.n22 VGND 0.04632f
C36501 _459_.CLK.t43 VGND 0.05003f
C36502 _459_.CLK.t21 VGND 0.05332f
C36503 _459_.CLK.n23 VGND 0.07878f
C36504 _459_.CLK.n24 VGND 0.09826f
C36505 _459_.CLK.t18 VGND 0.05003f
C36506 _459_.CLK.t42 VGND 0.05332f
C36507 _459_.CLK.n25 VGND 0.07887f
C36508 _459_.CLK.t39 VGND 0.05003f
C36509 _459_.CLK.t45 VGND 0.05332f
C36510 _459_.CLK.n26 VGND 0.07878f
C36511 _459_.CLK.n27 VGND 0.04384f
C36512 _459_.CLK.n28 VGND 0.86155f
C36513 _459_.CLK.n29 VGND 0.95978f
C36514 _459_.CLK.t28 VGND 0.05353f
C36515 _459_.CLK.t17 VGND 0.04981f
C36516 _459_.CLK.n30 VGND 0.07879f
C36517 _459_.CLK.n31 VGND 0.04632f
C36518 _459_.CLK.n32 VGND 0.6002f
C36519 _459_.CLK.n33 VGND 0.81274f
C36520 _459_.CLK.n34 VGND 0.64432f
C36521 _459_.CLK.n35 VGND 0.54199f
C36522 _459_.CLK.t27 VGND 0.05353f
C36523 _459_.CLK.t48 VGND 0.04981f
C36524 _459_.CLK.n36 VGND 0.07879f
C36525 _459_.CLK.n37 VGND 0.41739f
C36526 _459_.CLK.t34 VGND 0.05003f
C36527 _459_.CLK.t30 VGND 0.05332f
C36528 _459_.CLK.n38 VGND 0.07878f
C36529 _459_.CLK.n39 VGND 0.05083f
C36530 _459_.CLK.n40 VGND 1.22035f
C36531 _459_.CLK.n41 VGND 0.82849f
C36532 _459_.CLK.t32 VGND 0.05353f
C36533 _459_.CLK.t46 VGND 0.04981f
C36534 _459_.CLK.n42 VGND 0.07879f
C36535 _459_.CLK.n43 VGND 0.05904f
C36536 _459_.CLK.n44 VGND 0.20183f
C36537 _459_.CLK.t22 VGND 0.05003f
C36538 _459_.CLK.t36 VGND 0.05332f
C36539 _459_.CLK.n45 VGND 0.07878f
C36540 _459_.CLK.n46 VGND 0.14908f
C36541 _459_.CLK.n47 VGND 0.57697f
C36542 _459_.CLK.t38 VGND 0.05353f
C36543 _459_.CLK.t41 VGND 0.04981f
C36544 _459_.CLK.n48 VGND 0.07879f
C36545 _459_.CLK.n49 VGND 0.05904f
C36546 _459_.CLK.n50 VGND 0.37711f
C36547 _459_.CLK.t20 VGND 0.05003f
C36548 _459_.CLK.t40 VGND 0.05332f
C36549 _459_.CLK.n51 VGND 0.07887f
C36550 _459_.CLK.n52 VGND 0.94986f
C36551 _459_.CLK.t26 VGND 0.05353f
C36552 _459_.CLK.t35 VGND 0.04981f
C36553 _459_.CLK.n53 VGND 0.07888f
C36554 _459_.CLK.n54 VGND 1.10469f
C36555 _459_.CLK.n55 VGND 1.08325f
C36556 _459_.CLK.n56 VGND 0.34499f
C36557 _459_.CLK.n57 VGND 0.12218f
C36558 _459_.CLK.n58 VGND 0.09896f
C36559 _459_.CLK.t1 VGND 0.03777f
C36560 _459_.CLK.t0 VGND 0.03777f
C36561 _459_.CLK.n59 VGND 0.09439f
C36562 _459_.CLK.t4 VGND 0.03777f
C36563 _459_.CLK.t7 VGND 0.03777f
C36564 _459_.CLK.n60 VGND 0.07648f
C36565 _459_.CLK.n61 VGND 0.19982f
C36566 _459_.CLK.n62 VGND 0.07994f
C36567 a_43440_19325.t1 VGND 0.04354f
C36568 a_43440_19325.t6 VGND 0.0394f
C36569 a_43440_19325.t3 VGND 0.13194f
C36570 a_43440_19325.t7 VGND 0.1164f
C36571 a_43440_19325.n0 VGND 0.15078f
C36572 a_43440_19325.n1 VGND 0.05139f
C36573 a_43440_19325.n2 VGND 0.19448f
C36574 a_43440_19325.t5 VGND 0.01856f
C36575 a_43440_19325.t2 VGND 0.11668f
C36576 a_43440_19325.t4 VGND 0.36673f
C36577 a_43440_19325.n3 VGND 0.23553f
C36578 a_43440_19325.n4 VGND 0.53889f
C36579 a_43440_19325.t0 VGND 0.09569f
C36580 _284_.ZN.t32 VGND 0.09925f
C36581 _284_.ZN.n0 VGND 0.06508f
C36582 _284_.ZN.t20 VGND 0.09925f
C36583 _284_.ZN.t37 VGND 0.09124f
C36584 _284_.ZN.n1 VGND 0.10079f
C36585 _284_.ZN.t35 VGND 0.09124f
C36586 _284_.ZN.n2 VGND 0.10079f
C36587 _284_.ZN.n3 VGND 0.06236f
C36588 _284_.ZN.n4 VGND 0.1628f
C36589 _284_.ZN.t13 VGND 0.0316f
C36590 _284_.ZN.t14 VGND 0.0316f
C36591 _284_.ZN.n5 VGND 0.13363f
C36592 _284_.ZN.t12 VGND 0.0316f
C36593 _284_.ZN.t15 VGND 0.0316f
C36594 _284_.ZN.n6 VGND 0.0632f
C36595 _284_.ZN.n7 VGND 0.34613f
C36596 _284_.ZN.t1 VGND 0.04306f
C36597 _284_.ZN.t8 VGND 0.01289f
C36598 _284_.ZN.n8 VGND 0.08964f
C36599 _284_.ZN.t9 VGND 0.02367f
C36600 _284_.ZN.t3 VGND 0.02367f
C36601 _284_.ZN.n9 VGND 0.04733f
C36602 _284_.ZN.n10 VGND 0.17265f
C36603 _284_.ZN.t2 VGND 0.02367f
C36604 _284_.ZN.t10 VGND 0.02367f
C36605 _284_.ZN.n11 VGND 0.04733f
C36606 _284_.ZN.n12 VGND 0.11437f
C36607 _284_.ZN.t11 VGND 0.01289f
C36608 _284_.ZN.n13 VGND 0.00844f
C36609 _284_.ZN.t0 VGND 0.00278f
C36610 _284_.ZN.n14 VGND 0.05235f
C36611 _284_.ZN.n15 VGND 0.06103f
C36612 _284_.ZN.n16 VGND 0.14164f
C36613 _284_.ZN.n17 VGND 0.16273f
C36614 _284_.ZN.t5 VGND 0.02843f
C36615 _284_.ZN.t17 VGND 0.02843f
C36616 _284_.ZN.n18 VGND 0.06876f
C36617 _284_.ZN.t19 VGND 0.02843f
C36618 _284_.ZN.t6 VGND 0.02843f
C36619 _284_.ZN.n19 VGND 0.05685f
C36620 _284_.ZN.n20 VGND 0.2831f
C36621 _284_.ZN.t4 VGND 0.02843f
C36622 _284_.ZN.t18 VGND 0.02843f
C36623 _284_.ZN.n21 VGND 0.05685f
C36624 _284_.ZN.n22 VGND 0.16703f
C36625 _284_.ZN.t16 VGND 0.02843f
C36626 _284_.ZN.t7 VGND 0.02843f
C36627 _284_.ZN.n23 VGND 0.05685f
C36628 _284_.ZN.n24 VGND 0.1092f
C36629 _284_.ZN.n25 VGND 1.20891f
C36630 _284_.ZN.t21 VGND 0.09925f
C36631 _284_.ZN.n26 VGND 0.06508f
C36632 _284_.ZN.t30 VGND 0.09925f
C36633 _284_.ZN.t22 VGND 0.09124f
C36634 _284_.ZN.n27 VGND 0.10079f
C36635 _284_.ZN.t36 VGND 0.09124f
C36636 _284_.ZN.n28 VGND 0.10079f
C36637 _284_.ZN.n29 VGND 0.06236f
C36638 _284_.ZN.n30 VGND 0.12302f
C36639 _284_.ZN.t33 VGND 0.09925f
C36640 _284_.ZN.n31 VGND 0.06619f
C36641 _284_.ZN.t28 VGND 0.09925f
C36642 _284_.ZN.t29 VGND 0.09124f
C36643 _284_.ZN.t24 VGND 0.09124f
C36644 _284_.ZN.n32 VGND 0.10079f
C36645 _284_.ZN.n33 VGND 0.10079f
C36646 _284_.ZN.n34 VGND 0.06236f
C36647 _284_.ZN.n35 VGND 0.19438f
C36648 _284_.ZN.n36 VGND 0.05541f
C36649 _284_.ZN.n37 VGND 1.51446f
C36650 _284_.ZN.t25 VGND 0.08491f
C36651 _284_.ZN.t34 VGND 0.09283f
C36652 _284_.ZN.n38 VGND 0.15381f
C36653 _284_.ZN.t31 VGND 0.13114f
C36654 _284_.ZN.n39 VGND 0.09614f
C36655 _284_.ZN.n40 VGND 0.50835f
C36656 _284_.ZN.n41 VGND 0.12771f
C36657 _284_.ZN.t38 VGND 0.09925f
C36658 _284_.ZN.t27 VGND 0.09925f
C36659 _284_.ZN.n42 VGND 0.06263f
C36660 _284_.ZN.t23 VGND 0.09124f
C36661 _284_.ZN.n43 VGND 0.10079f
C36662 _284_.ZN.t26 VGND 0.09124f
C36663 _284_.ZN.n44 VGND 0.10079f
C36664 _284_.ZN.n45 VGND 0.06236f
C36665 _284_.ZN.n46 VGND 0.09946f
C36666 _397_.A2.t1 VGND 0.01144f
C36667 _397_.A2.t0 VGND 0.01144f
C36668 _397_.A2.n0 VGND 0.0231f
C36669 _397_.A2.t2 VGND 0.00769f
C36670 _397_.A2.t3 VGND 0.00769f
C36671 _397_.A2.n1 VGND 0.01548f
C36672 _397_.A2.t12 VGND 0.03416f
C36673 _397_.A2.t10 VGND 0.02474f
C36674 _397_.A2.n2 VGND 0.04316f
C36675 _397_.A2.n3 VGND 0.02983f
C36676 _397_.A2.t7 VGND 0.01941f
C36677 _397_.A2.t19 VGND 0.0357f
C36678 _397_.A2.n4 VGND 0.03705f
C36679 _397_.A2.n5 VGND 0.0351f
C36680 _397_.A2.t20 VGND 0.02791f
C36681 _397_.A2.t11 VGND 0.03588f
C36682 _397_.A2.n6 VGND 0.04045f
C36683 _397_.A2.n7 VGND 0.1468f
C36684 _397_.A2.t18 VGND 0.02374f
C36685 _397_.A2.n8 VGND 0.0182f
C36686 _397_.A2.t15 VGND 0.03488f
C36687 _397_.A2.n9 VGND 0.0325f
C36688 _397_.A2.t6 VGND 0.03488f
C36689 _397_.A2.n10 VGND 0.0325f
C36690 _397_.A2.t14 VGND 0.02374f
C36691 _397_.A2.n11 VGND 0.01855f
C36692 _397_.A2.t5 VGND 0.02747f
C36693 _397_.A2.t21 VGND 0.02614f
C36694 _397_.A2.n12 VGND 0.05088f
C36695 _397_.A2.n13 VGND 0.14699f
C36696 _397_.A2.t13 VGND 0.02903f
C36697 _397_.A2.t9 VGND 0.02915f
C36698 _397_.A2.n14 VGND 0.05017f
C36699 _397_.A2.t16 VGND 0.03105f
C36700 _397_.A2.t4 VGND 0.02628f
C36701 _397_.A2.n15 VGND 0.04326f
C36702 _397_.A2.n16 VGND 0.02288f
C36703 _397_.A2.n17 VGND 0.34067f
C36704 _397_.A2.n18 VGND 0.18723f
C36705 _397_.A2.n19 VGND 0.10227f
C36706 _397_.A2.t8 VGND 0.02474f
C36707 _397_.A2.t17 VGND 0.03416f
C36708 _397_.A2.n20 VGND 0.0434f
C36709 _397_.A2.n21 VGND 0.11838f
C36710 _397_.A2.n22 VGND 0.2545f
C36711 _397_.A2.n23 VGND 0.08896f
C36712 _371_.A1.t2 VGND 0.01526f
C36713 _371_.A1.t3 VGND 0.01526f
C36714 _371_.A1.n0 VGND 0.03416f
C36715 _371_.A1.t5 VGND 0.01833f
C36716 _371_.A1.t6 VGND 0.01833f
C36717 _371_.A1.n1 VGND 0.04222f
C36718 _371_.A1.t1 VGND 0.01833f
C36719 _371_.A1.t0 VGND 0.01833f
C36720 _371_.A1.n2 VGND 0.03667f
C36721 _371_.A1.n3 VGND 0.10564f
C36722 _371_.A1.t7 VGND 0.01833f
C36723 _371_.A1.t4 VGND 0.01833f
C36724 _371_.A1.n4 VGND 0.03667f
C36725 _371_.A1.n5 VGND 0.10897f
C36726 _371_.A1.t17 VGND 0.0655f
C36727 _371_.A1.t8 VGND 0.0489f
C36728 _371_.A1.n6 VGND 0.08091f
C36729 _371_.A1.n7 VGND 0.23471f
C36730 _371_.A1.t14 VGND 0.04393f
C36731 _371_.A1.t13 VGND 0.07373f
C36732 _371_.A1.n8 VGND 0.07686f
C36733 _371_.A1.n9 VGND 0.50601f
C36734 _371_.A1.t9 VGND 0.0618f
C36735 _371_.A1.n10 VGND 0.04472f
C36736 _371_.A1.t19 VGND 0.03522f
C36737 _371_.A1.n11 VGND 0.04399f
C36738 _371_.A1.t10 VGND 0.03522f
C36739 _371_.A1.t11 VGND 0.06449f
C36740 _371_.A1.n12 VGND 0.06802f
C36741 _371_.A1.t18 VGND 0.06449f
C36742 _371_.A1.n13 VGND 0.06802f
C36743 _371_.A1.n14 VGND 0.04252f
C36744 _371_.A1.n15 VGND 0.10235f
C36745 _371_.A1.t15 VGND 0.0481f
C36746 _371_.A1.n16 VGND 0.05678f
C36747 _371_.A1.t12 VGND 0.0481f
C36748 _371_.A1.n17 VGND 0.05678f
C36749 _371_.A1.t16 VGND 0.0618f
C36750 _371_.A1.n18 VGND 0.04357f
C36751 _371_.A1.n19 VGND 0.07624f
C36752 _371_.A1.n20 VGND 0.90908f
C36753 _371_.A1.n21 VGND 0.29973f
C36754 a_42820_29159.t4 VGND 0.12779f
C36755 a_42820_29159.t7 VGND 0.40165f
C36756 a_42820_29159.t5 VGND 0.02032f
C36757 a_42820_29159.n0 VGND 0.25796f
C36758 a_42820_29159.t1 VGND 0.1048f
C36759 a_42820_29159.n1 VGND 0.59021f
C36760 a_42820_29159.t2 VGND 0.14451f
C36761 a_42820_29159.t6 VGND 0.12788f
C36762 a_42820_29159.n2 VGND 0.16475f
C36763 a_42820_29159.t3 VGND 0.04268f
C36764 a_42820_29159.n3 VGND 0.05675f
C36765 a_42820_29159.n4 VGND 0.21301f
C36766 a_42820_29159.t0 VGND 0.04768f
C36767 _362_.B.t2 VGND 0.03697f
C36768 _362_.B.t3 VGND 0.03697f
C36769 _362_.B.n0 VGND 0.07446f
C36770 _362_.B.t5 VGND 0.17321f
C36771 _362_.B.t13 VGND 0.13307f
C36772 _362_.B.n1 VGND 0.22906f
C36773 _362_.B.n2 VGND 0.16416f
C36774 _362_.B.t16 VGND 0.15709f
C36775 _362_.B.t10 VGND 0.13307f
C36776 _362_.B.n3 VGND 0.11313f
C36777 _362_.B.n4 VGND 0.13342f
C36778 _362_.B.t8 VGND 0.15709f
C36779 _362_.B.n5 VGND 0.13342f
C36780 _362_.B.t15 VGND 0.13307f
C36781 _362_.B.n6 VGND 0.11313f
C36782 _362_.B.n7 VGND 0.17819f
C36783 _362_.B.t18 VGND 0.17328f
C36784 _362_.B.t12 VGND 0.13307f
C36785 _362_.B.n8 VGND 0.21019f
C36786 _362_.B.n9 VGND 0.3723f
C36787 _362_.B.t19 VGND 0.0982f
C36788 _362_.B.t4 VGND 0.12527f
C36789 _362_.B.n10 VGND 0.20587f
C36790 _362_.B.n11 VGND 0.86217f
C36791 _362_.B.t11 VGND 0.15118f
C36792 _362_.B.t6 VGND 0.15388f
C36793 _362_.B.n12 VGND 0.2101f
C36794 _362_.B.n13 VGND 1.18499f
C36795 _362_.B.t21 VGND 0.16133f
C36796 _362_.B.t9 VGND 0.14564f
C36797 _362_.B.n14 VGND 0.21407f
C36798 _362_.B.t20 VGND 0.12192f
C36799 _362_.B.t17 VGND 0.17945f
C36800 _362_.B.n15 VGND 0.20577f
C36801 _362_.B.n16 VGND 0.16722f
C36802 _362_.B.n17 VGND 0.1387f
C36803 _362_.B.t14 VGND 0.17858f
C36804 _362_.B.t7 VGND 0.10595f
C36805 _362_.B.n18 VGND 0.18662f
C36806 _362_.B.n19 VGND 0.8014f
C36807 _362_.B.n20 VGND 0.37849f
C36808 _362_.B.t1 VGND 0.055f
C36809 _362_.B.t0 VGND 0.055f
C36810 _362_.B.n21 VGND 0.11108f
C36811 a_48272_25156.t6 VGND 0.05842f
C36812 a_48272_25156.t3 VGND 0.05842f
C36813 a_48272_25156.t5 VGND 0.04219f
C36814 a_48272_25156.n0 VGND 0.10181f
C36815 a_48272_25156.t4 VGND 0.05842f
C36816 a_48272_25156.t2 VGND 0.04219f
C36817 a_48272_25156.n1 VGND 0.10181f
C36818 a_48272_25156.t1 VGND 0.05842f
C36819 a_48272_25156.t0 VGND 0.04219f
C36820 a_48272_25156.n2 VGND 0.10181f
C36821 a_48272_25156.t9 VGND 0.05178f
C36822 a_48272_25156.t12 VGND 0.02084f
C36823 a_48272_25156.t10 VGND 0.02084f
C36824 a_48272_25156.n3 VGND 0.04236f
C36825 a_48272_25156.t11 VGND 0.02084f
C36826 a_48272_25156.t13 VGND 0.02084f
C36827 a_48272_25156.n4 VGND 0.04236f
C36828 a_48272_25156.t8 VGND 0.06562f
C36829 a_48272_25156.n5 VGND 0.41703f
C36830 a_48272_25156.n6 VGND 0.25146f
C36831 a_48272_25156.n7 VGND 0.20883f
C36832 a_48272_25156.t37 VGND 0.12051f
C36833 a_48272_25156.t31 VGND 0.12111f
C36834 a_48272_25156.t17 VGND 0.18298f
C36835 a_48272_25156.n8 VGND 0.26923f
C36836 a_48272_25156.t36 VGND 0.12111f
C36837 a_48272_25156.t23 VGND 0.18298f
C36838 a_48272_25156.n9 VGND 0.30628f
C36839 a_48272_25156.t35 VGND 0.12111f
C36840 a_48272_25156.t20 VGND 0.18298f
C36841 a_48272_25156.n10 VGND 0.30628f
C36842 a_48272_25156.t26 VGND 0.12111f
C36843 a_48272_25156.t45 VGND 0.18298f
C36844 a_48272_25156.n11 VGND -0.57472f
C36845 a_48272_25156.t22 VGND 0.12111f
C36846 a_48272_25156.t42 VGND 0.18298f
C36847 a_48272_25156.n12 VGND 0.30628f
C36848 a_48272_25156.t16 VGND 0.12111f
C36849 a_48272_25156.t38 VGND 0.18298f
C36850 a_48272_25156.n13 VGND 0.30628f
C36851 a_48272_25156.t21 VGND 0.12111f
C36852 a_48272_25156.t40 VGND 0.18298f
C36853 a_48272_25156.n14 VGND 0.30628f
C36854 a_48272_25156.t41 VGND 0.12111f
C36855 a_48272_25156.t30 VGND 0.18298f
C36856 a_48272_25156.n15 VGND 0.30628f
C36857 a_48272_25156.t44 VGND 0.12111f
C36858 a_48272_25156.t34 VGND 0.18298f
C36859 a_48272_25156.n16 VGND 0.30628f
C36860 a_48272_25156.t39 VGND 0.12111f
C36861 a_48272_25156.t29 VGND 0.18298f
C36862 a_48272_25156.n17 VGND 0.30628f
C36863 a_48272_25156.t25 VGND 0.18298f
C36864 a_48272_25156.n18 VGND 0.15465f
C36865 a_48272_25156.n19 VGND 0.15324f
C36866 a_48272_25156.t33 VGND 0.12051f
C36867 a_48272_25156.n20 VGND 0.15324f
C36868 a_48272_25156.t19 VGND 0.18298f
C36869 a_48272_25156.n21 VGND 0.15465f
C36870 a_48272_25156.t24 VGND 0.12111f
C36871 a_48272_25156.t43 VGND 0.18298f
C36872 a_48272_25156.n22 VGND 0.26923f
C36873 a_48272_25156.t27 VGND 0.12111f
C36874 a_48272_25156.t14 VGND 0.18298f
C36875 a_48272_25156.n23 VGND 0.30628f
C36876 a_48272_25156.t32 VGND 0.12111f
C36877 a_48272_25156.t18 VGND 0.18298f
C36878 a_48272_25156.n24 VGND 0.30628f
C36879 a_48272_25156.t28 VGND 0.12111f
C36880 a_48272_25156.t15 VGND 0.18298f
C36881 a_48272_25156.n25 VGND 0.83832f
C36882 a_48272_25156.n26 VGND 0.58145f
C36883 a_48272_25156.n27 VGND 0.21258f
C36884 a_48272_25156.n28 VGND 0.26004f
C36885 a_48272_25156.n29 VGND 0.40497f
C36886 a_48272_25156.n30 VGND 0.12544f
C36887 a_48272_25156.t7 VGND 0.04219f
C36888 _350_.A2.t15 VGND 0.01857f
C36889 _350_.A2.t7 VGND 0.06204f
C36890 _350_.A2.n0 VGND 0.12915f
C36891 _350_.A2.t4 VGND 0.0341f
C36892 _350_.A2.t9 VGND 0.0341f
C36893 _350_.A2.n1 VGND 0.06819f
C36894 _350_.A2.n2 VGND 0.24875f
C36895 _350_.A2.t11 VGND 0.0341f
C36896 _350_.A2.t6 VGND 0.0341f
C36897 _350_.A2.n3 VGND 0.06819f
C36898 _350_.A2.n4 VGND 0.16479f
C36899 _350_.A2.t5 VGND 0.06204f
C36900 _350_.A2.t12 VGND 0.01857f
C36901 _350_.A2.n5 VGND 0.11747f
C36902 _350_.A2.n6 VGND 0.20407f
C36903 _350_.A2.t17 VGND 0.04096f
C36904 _350_.A2.t0 VGND 0.04096f
C36905 _350_.A2.n7 VGND 0.09907f
C36906 _350_.A2.t2 VGND 0.04096f
C36907 _350_.A2.t18 VGND 0.04096f
C36908 _350_.A2.n8 VGND 0.08192f
C36909 _350_.A2.n9 VGND 0.40789f
C36910 _350_.A2.t16 VGND 0.04096f
C36911 _350_.A2.t1 VGND 0.04096f
C36912 _350_.A2.n10 VGND 0.08192f
C36913 _350_.A2.n11 VGND 0.24066f
C36914 _350_.A2.t3 VGND 0.04096f
C36915 _350_.A2.t19 VGND 0.04096f
C36916 _350_.A2.n12 VGND 0.08192f
C36917 _350_.A2.n13 VGND 0.19205f
C36918 _350_.A2.n14 VGND 0.26451f
C36919 _350_.A2.t14 VGND 0.04553f
C36920 _350_.A2.t10 VGND 0.04553f
C36921 _350_.A2.n15 VGND 0.09247f
C36922 _350_.A2.t26 VGND 0.15233f
C36923 _350_.A2.t28 VGND 0.13176f
C36924 _350_.A2.n16 VGND 0.17886f
C36925 _350_.A2.t21 VGND 0.18203f
C36926 _350_.A2.t20 VGND 0.10316f
C36927 _350_.A2.n17 VGND 0.22116f
C36928 _350_.A2.n18 VGND 0.07718f
C36929 _350_.A2.t25 VGND 0.16593f
C36930 _350_.A2.t29 VGND 0.1113f
C36931 _350_.A2.n19 VGND 0.07054f
C36932 _350_.A2.n20 VGND 0.13685f
C36933 _350_.A2.t22 VGND 0.16516f
C36934 _350_.A2.n21 VGND 0.13982f
C36935 _350_.A2.t27 VGND 0.10316f
C36936 _350_.A2.n22 VGND 0.0878f
C36937 _350_.A2.n23 VGND 0.17183f
C36938 _350_.A2.t23 VGND 0.14234f
C36939 _350_.A2.t24 VGND 0.15321f
C36940 _350_.A2.n24 VGND 0.17786f
C36941 _350_.A2.n25 VGND 0.21734f
C36942 _350_.A2.n26 VGND 1.54464f
C36943 _350_.A2.n27 VGND 0.57327f
C36944 _350_.A2.t8 VGND 0.04553f
C36945 _350_.A2.t13 VGND 0.04553f
C36946 _350_.A2.n28 VGND 0.09106f
C36947 _350_.A2.n29 VGND 0.28527f
C36948 _447_.Q.t1 VGND 0.04265f
C36949 _447_.Q.t0 VGND 0.06051f
C36950 _447_.Q.t14 VGND 0.06628f
C36951 _447_.Q.t12 VGND 0.05156f
C36952 _447_.Q.n0 VGND 0.07473f
C36953 _447_.Q.t2 VGND 0.05156f
C36954 _447_.Q.t5 VGND 0.06628f
C36955 _447_.Q.n1 VGND 0.07473f
C36956 _447_.Q.n2 VGND 0.99284f
C36957 _447_.Q.t4 VGND 0.05416f
C36958 _447_.Q.t11 VGND 0.06656f
C36959 _447_.Q.n3 VGND 0.08513f
C36960 _447_.Q.n4 VGND 0.03573f
C36961 _447_.Q.n5 VGND 0.12666f
C36962 _447_.Q.t16 VGND 0.03943f
C36963 _447_.Q.t10 VGND 0.0493f
C36964 _447_.Q.n6 VGND 0.07755f
C36965 _447_.Q.n7 VGND 0.06364f
C36966 _447_.Q.n8 VGND 0.18924f
C36967 _447_.Q.t13 VGND 0.06861f
C36968 _447_.Q.t6 VGND 0.04071f
C36969 _447_.Q.n9 VGND 0.07247f
C36970 _447_.Q.n10 VGND 0.11564f
C36971 _447_.Q.t17 VGND 0.07028f
C36972 _447_.Q.t9 VGND 0.04384f
C36973 _447_.Q.n11 VGND 0.08351f
C36974 _447_.Q.n12 VGND 0.28713f
C36975 _447_.Q.n13 VGND 0.18513f
C36976 _447_.Q.t7 VGND 0.04088f
C36977 _447_.Q.t8 VGND 0.06861f
C36978 _447_.Q.n14 VGND 0.07153f
C36979 _447_.Q.n15 VGND 0.2346f
C36980 _447_.Q.t15 VGND 0.0488f
C36981 _447_.Q.t3 VGND 0.03531f
C36982 _447_.Q.n16 VGND 0.0763f
C36983 _447_.Q.n17 VGND 0.36518f
C36984 a_54864_22461.t1 VGND 0.04561f
C36985 a_54864_22461.t3 VGND 0.04128f
C36986 a_54864_22461.t6 VGND 0.13823f
C36987 a_54864_22461.t4 VGND 0.12194f
C36988 a_54864_22461.n0 VGND 0.15796f
C36989 a_54864_22461.n1 VGND 0.05384f
C36990 a_54864_22461.n2 VGND 0.20374f
C36991 a_54864_22461.t7 VGND 0.01944f
C36992 a_54864_22461.t5 VGND 0.12223f
C36993 a_54864_22461.t2 VGND 0.38419f
C36994 a_54864_22461.n3 VGND 0.24674f
C36995 a_54864_22461.n4 VGND 0.56455f
C36996 a_54864_22461.t0 VGND 0.10024f
C36997 _304_.A1.t1 VGND 0.04602f
C36998 _304_.A1.t0 VGND 0.06528f
C36999 _304_.A1.t6 VGND 0.07402f
C37000 _304_.A1.t4 VGND 0.04392f
C37001 _304_.A1.n0 VGND 0.07735f
C37002 _304_.A1.t15 VGND 0.05264f
C37003 _304_.A1.t14 VGND 0.0381f
C37004 _304_.A1.n1 VGND 0.08231f
C37005 _304_.A1.n2 VGND 0.32783f
C37006 _304_.A1.t12 VGND 0.04657f
C37007 _304_.A1.n3 VGND 0.04347f
C37008 _304_.A1.t11 VGND 0.04657f
C37009 _304_.A1.t10 VGND 0.06506f
C37010 _304_.A1.n4 VGND 0.05522f
C37011 _304_.A1.t17 VGND 0.06506f
C37012 _304_.A1.n5 VGND 0.05522f
C37013 _304_.A1.n6 VGND 0.04226f
C37014 _304_.A1.n7 VGND 0.10744f
C37015 _304_.A1.t3 VGND 0.04254f
C37016 _304_.A1.t7 VGND 0.05318f
C37017 _304_.A1.n8 VGND 0.08444f
C37018 _304_.A1.n9 VGND 0.67002f
C37019 _304_.A1.t5 VGND 0.07402f
C37020 _304_.A1.t13 VGND 0.04392f
C37021 _304_.A1.n10 VGND 0.08052f
C37022 _304_.A1.n11 VGND 0.35577f
C37023 _304_.A1.t9 VGND 0.07582f
C37024 _304_.A1.t2 VGND 0.0473f
C37025 _304_.A1.n12 VGND 0.09004f
C37026 _304_.A1.n13 VGND 0.05591f
C37027 _304_.A1.n14 VGND 0.27872f
C37028 _304_.A1.t8 VGND 0.0407f
C37029 _304_.A1.t16 VGND 0.05192f
C37030 _304_.A1.n15 VGND 0.08531f
C37031 _304_.A1.n16 VGND 0.39688f
C37032 _304_.A1.n17 VGND 0.21642f
C37033 _424_.B1.t4 VGND 0.01646f
C37034 _424_.B1.t5 VGND 0.01646f
C37035 _424_.B1.n0 VGND 0.05291f
C37036 _424_.B1.t1 VGND 0.02268f
C37037 _424_.B1.t2 VGND 0.02268f
C37038 _424_.B1.n1 VGND 0.04619f
C37039 _424_.B1.n2 VGND 0.23476f
C37040 _424_.B1.t8 VGND 0.05597f
C37041 _424_.B1.t10 VGND 0.05881f
C37042 _424_.B1.n3 VGND 0.10894f
C37043 _424_.B1.n4 VGND 0.05005f
C37044 _424_.B1.t13 VGND 0.06878f
C37045 _424_.B1.t14 VGND 0.07241f
C37046 _424_.B1.n5 VGND 0.09739f
C37047 _424_.B1.t15 VGND 0.07241f
C37048 _424_.B1.t7 VGND 0.06878f
C37049 _424_.B1.n6 VGND 0.09739f
C37050 _424_.B1.n7 VGND 0.8962f
C37051 _424_.B1.n8 VGND 0.44283f
C37052 _424_.B1.t11 VGND 0.07241f
C37053 _424_.B1.t6 VGND 0.06878f
C37054 _424_.B1.n9 VGND 0.09739f
C37055 _424_.B1.t9 VGND 0.07241f
C37056 _424_.B1.t12 VGND 0.06878f
C37057 _424_.B1.n10 VGND 0.09739f
C37058 _424_.B1.n11 VGND 1.02392f
C37059 _424_.B1.n12 VGND 0.41013f
C37060 _424_.B1.t3 VGND 0.02268f
C37061 _424_.B1.t0 VGND 0.02268f
C37062 _424_.B1.n13 VGND 0.04683f
C37063 _424_.B1.n14 VGND 0.10311f
C37064 a_36548_27591.t6 VGND 0.12779f
C37065 a_36548_27591.t2 VGND 0.40165f
C37066 a_36548_27591.t5 VGND 0.02032f
C37067 a_36548_27591.n0 VGND 0.25796f
C37068 a_36548_27591.t4 VGND 0.14451f
C37069 a_36548_27591.t3 VGND 0.12788f
C37070 a_36548_27591.n1 VGND 0.16475f
C37071 a_36548_27591.t7 VGND 0.04268f
C37072 a_36548_27591.n2 VGND 0.05675f
C37073 a_36548_27591.t1 VGND 0.04768f
C37074 a_36548_27591.n3 VGND 0.21301f
C37075 a_36548_27591.n4 VGND 0.59021f
C37076 a_36548_27591.t0 VGND 0.1048f
C37077 _452_.CLK.t14 VGND 0.02766f
C37078 _452_.CLK.t8 VGND 0.0383f
C37079 _452_.CLK.n0 VGND 0.07886f
C37080 _452_.CLK.t10 VGND 0.02766f
C37081 _452_.CLK.t9 VGND 0.0383f
C37082 _452_.CLK.n1 VGND 0.06597f
C37083 _452_.CLK.n2 VGND 0.30738f
C37084 _452_.CLK.t24 VGND 0.02766f
C37085 _452_.CLK.t27 VGND 0.0383f
C37086 _452_.CLK.n3 VGND 0.06597f
C37087 _452_.CLK.n4 VGND 0.21097f
C37088 _452_.CLK.t25 VGND 0.02766f
C37089 _452_.CLK.t28 VGND 0.0383f
C37090 _452_.CLK.n5 VGND 0.06597f
C37091 _452_.CLK.n6 VGND 0.12776f
C37092 _452_.CLK.t18 VGND 0.0383f
C37093 _452_.CLK.t20 VGND 0.02766f
C37094 _452_.CLK.n7 VGND 0.07778f
C37095 _452_.CLK.t16 VGND 0.02766f
C37096 _452_.CLK.t11 VGND 0.0383f
C37097 _452_.CLK.n8 VGND 0.06597f
C37098 _452_.CLK.n9 VGND 0.29835f
C37099 _452_.CLK.t6 VGND 0.02766f
C37100 _452_.CLK.t2 VGND 0.0383f
C37101 _452_.CLK.n10 VGND 0.06597f
C37102 _452_.CLK.n11 VGND 0.21097f
C37103 _452_.CLK.t5 VGND 0.02766f
C37104 _452_.CLK.t1 VGND 0.0383f
C37105 _452_.CLK.n12 VGND 0.06597f
C37106 _452_.CLK.n13 VGND 0.13535f
C37107 _452_.CLK.n14 VGND 0.17218f
C37108 _452_.CLK.t12 VGND 0.011f
C37109 _452_.CLK.t31 VGND 0.011f
C37110 _452_.CLK.n15 VGND 0.02229f
C37111 _452_.CLK.t13 VGND 0.011f
C37112 _452_.CLK.t7 VGND 0.011f
C37113 _452_.CLK.n16 VGND 0.02229f
C37114 _452_.CLK.t22 VGND 0.011f
C37115 _452_.CLK.t4 VGND 0.011f
C37116 _452_.CLK.n17 VGND 0.02229f
C37117 _452_.CLK.t23 VGND 0.011f
C37118 _452_.CLK.t26 VGND 0.011f
C37119 _452_.CLK.n18 VGND 0.02415f
C37120 _452_.CLK.t59 VGND 0.05075f
C37121 _452_.CLK.t50 VGND 0.05407f
C37122 _452_.CLK.n19 VGND 0.0799f
C37123 _452_.CLK.n20 VGND 0.04698f
C37124 _452_.CLK.t53 VGND 0.05075f
C37125 _452_.CLK.t42 VGND 0.05407f
C37126 _452_.CLK.n21 VGND 0.07999f
C37127 _452_.CLK.t34 VGND 0.05075f
C37128 _452_.CLK.t41 VGND 0.05407f
C37129 _452_.CLK.n22 VGND 0.0799f
C37130 _452_.CLK.n23 VGND 0.05988f
C37131 _452_.CLK.n24 VGND 1.00819f
C37132 _452_.CLK.t38 VGND 0.05429f
C37133 _452_.CLK.t32 VGND 0.05052f
C37134 _452_.CLK.n25 VGND 0.07991f
C37135 _452_.CLK.n26 VGND 0.1512f
C37136 _452_.CLK.n27 VGND 0.83003f
C37137 _452_.CLK.t55 VGND 0.05429f
C37138 _452_.CLK.t39 VGND 0.05052f
C37139 _452_.CLK.n28 VGND 0.07991f
C37140 _452_.CLK.n29 VGND 0.04698f
C37141 _452_.CLK.n30 VGND 0.96119f
C37142 _452_.CLK.n31 VGND 0.53183f
C37143 _452_.CLK.t47 VGND 0.05075f
C37144 _452_.CLK.t56 VGND 0.05407f
C37145 _452_.CLK.n32 VGND 0.0799f
C37146 _452_.CLK.n33 VGND 0.04698f
C37147 _452_.CLK.n34 VGND 0.52042f
C37148 _452_.CLK.t45 VGND 0.05075f
C37149 _452_.CLK.t46 VGND 0.05407f
C37150 _452_.CLK.n35 VGND 0.07999f
C37151 _452_.CLK.n36 VGND 0.60594f
C37152 _452_.CLK.t52 VGND 0.05075f
C37153 _452_.CLK.t36 VGND 0.05407f
C37154 _452_.CLK.n37 VGND 0.0799f
C37155 _452_.CLK.n38 VGND 0.04759f
C37156 _452_.CLK.n39 VGND 0.82345f
C37157 _452_.CLK.t43 VGND 0.05429f
C37158 _452_.CLK.t58 VGND 0.05052f
C37159 _452_.CLK.n40 VGND 0.08f
C37160 _452_.CLK.n41 VGND 0.85006f
C37161 _452_.CLK.t51 VGND 0.05429f
C37162 _452_.CLK.t49 VGND 0.05052f
C37163 _452_.CLK.n42 VGND 0.08f
C37164 _452_.CLK.n43 VGND 0.96701f
C37165 _452_.CLK.t48 VGND 0.05075f
C37166 _452_.CLK.t35 VGND 0.05407f
C37167 _452_.CLK.n44 VGND 0.0799f
C37168 _452_.CLK.n45 VGND 0.1512f
C37169 _452_.CLK.n46 VGND 0.64129f
C37170 _452_.CLK.t54 VGND 0.05075f
C37171 _452_.CLK.t40 VGND 0.05407f
C37172 _452_.CLK.n47 VGND 0.0799f
C37173 _452_.CLK.n48 VGND 0.04698f
C37174 _452_.CLK.n49 VGND 0.39739f
C37175 _452_.CLK.t33 VGND 0.05429f
C37176 _452_.CLK.t37 VGND 0.05052f
C37177 _452_.CLK.n50 VGND 0.08f
C37178 _452_.CLK.n51 VGND 0.21817f
C37179 _452_.CLK.t44 VGND 0.05075f
C37180 _452_.CLK.t57 VGND 0.05407f
C37181 _452_.CLK.n52 VGND 0.07999f
C37182 _452_.CLK.n53 VGND 0.57283f
C37183 _452_.CLK.n54 VGND 0.24491f
C37184 _452_.CLK.n55 VGND 0.1218f
C37185 _452_.CLK.n56 VGND 0.1458f
C37186 _452_.CLK.n57 VGND 0.10128f
C37187 _452_.CLK.t29 VGND 0.011f
C37188 _452_.CLK.t21 VGND 0.011f
C37189 _452_.CLK.n58 VGND 0.02229f
C37190 _452_.CLK.t17 VGND 0.011f
C37191 _452_.CLK.t15 VGND 0.011f
C37192 _452_.CLK.n59 VGND 0.02229f
C37193 _452_.CLK.t19 VGND 0.011f
C37194 _452_.CLK.t3 VGND 0.011f
C37195 _452_.CLK.n60 VGND 0.03029f
C37196 _452_.CLK.n61 VGND 0.2275f
C37197 _452_.CLK.n62 VGND 0.1458f
C37198 _452_.CLK.t30 VGND 0.011f
C37199 _452_.CLK.t0 VGND 0.011f
C37200 _452_.CLK.n63 VGND 0.02229f
C37201 _452_.CLK.n64 VGND 0.10268f
C37202 _452_.CLK.n65 VGND 0.10843f
C37203 _350_.A1.t0 VGND 0.03087f
C37204 _350_.A1.t1 VGND 0.02176f
C37205 _350_.A1.t5 VGND 0.035f
C37206 _350_.A1.t9 VGND 0.02077f
C37207 _350_.A1.n0 VGND 0.03658f
C37208 _350_.A1.t15 VGND 0.03381f
C37209 _350_.A1.t11 VGND 0.0263f
C37210 _350_.A1.n1 VGND 0.03812f
C37211 _350_.A1.n2 VGND 0.1785f
C37212 _350_.A1.t2 VGND 0.035f
C37213 _350_.A1.t12 VGND 0.02077f
C37214 _350_.A1.n3 VGND 0.03658f
C37215 _350_.A1.n4 VGND 0.4898f
C37216 _350_.A1.t8 VGND 0.03016f
C37217 _350_.A1.n5 VGND 0.02047f
C37218 _350_.A1.t7 VGND 0.03016f
C37219 _350_.A1.t14 VGND 0.03488f
C37220 _350_.A1.t10 VGND 0.03564f
C37221 _350_.A1.t4 VGND 0.02641f
C37222 _350_.A1.n6 VGND 0.04321f
C37223 _350_.A1.n7 VGND 0.02184f
C37224 _350_.A1.n8 VGND 0.02308f
C37225 _350_.A1.t6 VGND 0.03014f
C37226 _350_.A1.t13 VGND 0.03068f
C37227 _350_.A1.n9 VGND 0.02296f
C37228 _350_.A1.t3 VGND 0.03057f
C37229 _350_.A1.n10 VGND 0.02689f
C37230 _350_.A1.n11 VGND 0.0193f
C37231 _350_.A1.n12 VGND 0.00609f
C37232 _350_.A1.n13 VGND 0.08421f
C37233 _350_.A1.n14 VGND 0.18011f
C37234 _230_.I.t0 VGND 0.06294f
C37235 _230_.I.t1 VGND 0.04243f
C37236 _230_.I.t8 VGND 0.06279f
C37237 _230_.I.t11 VGND 0.06057f
C37238 _230_.I.n0 VGND 0.07672f
C37239 _230_.I.t12 VGND 0.05447f
C37240 _230_.I.t10 VGND 0.07393f
C37241 _230_.I.n1 VGND 0.07974f
C37242 _230_.I.n2 VGND 0.11321f
C37243 _230_.I.n3 VGND 0.40032f
C37244 _230_.I.t2 VGND 0.05828f
C37245 _230_.I.t13 VGND 0.06739f
C37246 _230_.I.n4 VGND 0.07912f
C37247 _230_.I.t15 VGND 0.03809f
C37248 _230_.I.t7 VGND 0.07004f
C37249 _230_.I.n5 VGND 0.0727f
C37250 _230_.I.n6 VGND 0.37077f
C37251 _230_.I.n7 VGND 0.41962f
C37252 _230_.I.t6 VGND 0.06572f
C37253 _230_.I.t5 VGND 0.04156f
C37254 _230_.I.n8 VGND 0.09824f
C37255 _230_.I.n9 VGND 0.40006f
C37256 _230_.I.n10 VGND 0.20443f
C37257 _230_.I.t3 VGND 0.04917f
C37258 _230_.I.t4 VGND 0.04418f
C37259 _230_.I.n11 VGND 0.09377f
C37260 _230_.I.t9 VGND 0.07305f
C37261 _230_.I.t14 VGND 0.05476f
C37262 _230_.I.n12 VGND 0.08335f
C37263 _230_.I.n13 VGND 0.07898f
C37264 _230_.I.n14 VGND 0.26898f
C37265 _230_.I.n15 VGND 0.10685f
C37266 a_42168_25640.t11 VGND 0.02949f
C37267 a_42168_25640.t1 VGND 0.09397f
C37268 a_42168_25640.t4 VGND 0.02949f
C37269 a_42168_25640.t5 VGND 0.02949f
C37270 a_42168_25640.n0 VGND 0.05898f
C37271 a_42168_25640.n1 VGND 0.24509f
C37272 a_42168_25640.t3 VGND 0.02949f
C37273 a_42168_25640.t2 VGND 0.02949f
C37274 a_42168_25640.n2 VGND 0.05898f
C37275 a_42168_25640.n3 VGND 0.14253f
C37276 a_42168_25640.t6 VGND 0.02949f
C37277 a_42168_25640.t7 VGND 0.02949f
C37278 a_42168_25640.n4 VGND 0.05898f
C37279 a_42168_25640.n5 VGND 0.14953f
C37280 a_42168_25640.t10 VGND 0.11041f
C37281 a_42168_25640.t8 VGND 0.02949f
C37282 a_42168_25640.t9 VGND 0.02949f
C37283 a_42168_25640.n6 VGND 0.05898f
C37284 a_42168_25640.n7 VGND 0.43444f
C37285 a_42168_25640.n8 VGND 0.23422f
C37286 a_42168_25640.n9 VGND 0.05898f
C37287 a_42168_25640.t0 VGND 0.02949f
C37288 _355_.C.t0 VGND 0.02489f
C37289 _355_.C.t1 VGND 0.01798f
C37290 _355_.C.n0 VGND 0.04402f
C37291 _355_.C.t2 VGND 0.01208f
C37292 _355_.C.t3 VGND 0.01208f
C37293 _355_.C.n1 VGND 0.02762f
C37294 _355_.C.t19 VGND 0.05186f
C37295 _355_.C.t21 VGND 0.03872f
C37296 _355_.C.n2 VGND 0.06406f
C37297 _355_.C.n3 VGND 0.10708f
C37298 _355_.C.t14 VGND 0.05838f
C37299 _355_.C.t23 VGND 0.03464f
C37300 _355_.C.n4 VGND 0.06166f
C37301 _355_.C.n5 VGND 0.05002f
C37302 _355_.C.t10 VGND 0.03888f
C37303 _355_.C.t15 VGND 0.05186f
C37304 _355_.C.n6 VGND 0.06437f
C37305 _355_.C.t17 VGND 0.05059f
C37306 _355_.C.t6 VGND 0.04197f
C37307 _355_.C.n7 VGND 0.06431f
C37308 _355_.C.n8 VGND 0.68078f
C37309 _355_.C.t13 VGND 0.05838f
C37310 _355_.C.t18 VGND 0.03464f
C37311 _355_.C.n9 VGND 0.06101f
C37312 _355_.C.t11 VGND 0.05838f
C37313 _355_.C.t12 VGND 0.03464f
C37314 _355_.C.n10 VGND 0.06166f
C37315 _355_.C.n11 VGND 0.2286f
C37316 _355_.C.n12 VGND 0.71976f
C37317 _355_.C.t4 VGND 0.03052f
C37318 _355_.C.t5 VGND 0.05611f
C37319 _355_.C.n13 VGND 0.05846f
C37320 _355_.C.n14 VGND 0.36667f
C37321 _355_.C.t22 VGND 0.03888f
C37322 _355_.C.t8 VGND 0.05186f
C37323 _355_.C.n15 VGND 0.06437f
C37324 _355_.C.n16 VGND 0.45042f
C37325 _355_.C.t20 VGND 0.05186f
C37326 _355_.C.t9 VGND 0.03872f
C37327 _355_.C.n17 VGND 0.06406f
C37328 _355_.C.n18 VGND 0.03387f
C37329 _355_.C.n19 VGND 0.48748f
C37330 _355_.C.t16 VGND 0.05838f
C37331 _355_.C.t7 VGND 0.03464f
C37332 _355_.C.n20 VGND 0.06166f
C37333 _355_.C.n21 VGND 0.04719f
C37334 _355_.C.n22 VGND 0.4682f
C37335 _355_.C.n23 VGND 0.29065f
C37336 _355_.C.n24 VGND 0.5916f
C37337 _355_.C.n25 VGND 0.20625f
C37338 a_41048_29816.t1 VGND 0.02319f
C37339 a_41048_29816.t2 VGND 0.02319f
C37340 a_41048_29816.t0 VGND 0.02319f
C37341 a_41048_29816.n0 VGND 0.04686f
C37342 a_41048_29816.t4 VGND 0.02055f
C37343 a_41048_29816.t5 VGND 0.00827f
C37344 a_41048_29816.t6 VGND 0.00827f
C37345 a_41048_29816.n1 VGND 0.02443f
C37346 a_41048_29816.n2 VGND 0.14305f
C37347 a_41048_29816.t12 VGND 0.04454f
C37348 a_41048_29816.t20 VGND 0.07341f
C37349 a_41048_29816.n3 VGND 0.10696f
C37350 a_41048_29816.t21 VGND 0.04454f
C37351 a_41048_29816.t22 VGND 0.07341f
C37352 a_41048_29816.n4 VGND 0.10993f
C37353 a_41048_29816.t15 VGND 0.04454f
C37354 a_41048_29816.t16 VGND 0.07341f
C37355 a_41048_29816.n5 VGND 0.10696f
C37356 a_41048_29816.t13 VGND 0.04454f
C37357 a_41048_29816.t9 VGND 0.07341f
C37358 a_41048_29816.n6 VGND -0.02869f
C37359 a_41048_29816.t17 VGND 0.04454f
C37360 a_41048_29816.t18 VGND 0.07341f
C37361 a_41048_29816.n7 VGND 0.12166f
C37362 a_41048_29816.t19 VGND 0.04454f
C37363 a_41048_29816.t11 VGND 0.07341f
C37364 a_41048_29816.n8 VGND 0.12166f
C37365 a_41048_29816.t7 VGND 0.04454f
C37366 a_41048_29816.t8 VGND 0.07341f
C37367 a_41048_29816.n9 VGND 0.12166f
C37368 a_41048_29816.t10 VGND 0.04454f
C37369 a_41048_29816.t14 VGND 0.07341f
C37370 a_41048_29816.n10 VGND 0.11869f
C37371 a_41048_29816.n11 VGND 0.07137f
C37372 a_41048_29816.n12 VGND 0.15897f
C37373 a_41048_29816.n13 VGND 0.1468f
C37374 a_41048_29816.n14 VGND 0.05624f
C37375 a_41048_29816.t3 VGND 0.02319f
C37376 vgaringosc.workerclkbuff_notouch_.I.t0 VGND 0.01068f
C37377 vgaringosc.workerclkbuff_notouch_.I.t2 VGND 0.01068f
C37378 vgaringosc.workerclkbuff_notouch_.I.n0 VGND 0.02263f
C37379 vgaringosc.workerclkbuff_notouch_.I.t3 VGND 0.01592f
C37380 vgaringosc.workerclkbuff_notouch_.I.t1 VGND 0.01592f
C37381 vgaringosc.workerclkbuff_notouch_.I.n1 VGND 0.03443f
C37382 vgaringosc.workerclkbuff_notouch_.I.t6 VGND 0.02373f
C37383 vgaringosc.workerclkbuff_notouch_.I.t8 VGND 0.04202f
C37384 vgaringosc.workerclkbuff_notouch_.I.n2 VGND 0.07248f
C37385 vgaringosc.workerclkbuff_notouch_.I.t5 VGND 0.02373f
C37386 vgaringosc.workerclkbuff_notouch_.I.t4 VGND 0.04202f
C37387 vgaringosc.workerclkbuff_notouch_.I.n3 VGND 0.0761f
C37388 vgaringosc.workerclkbuff_notouch_.I.t9 VGND 0.06373f
C37389 vgaringosc.workerclkbuff_notouch_.I.t10 VGND 0.02373f
C37390 vgaringosc.workerclkbuff_notouch_.I.t7 VGND 0.04202f
C37391 vgaringosc.workerclkbuff_notouch_.I.n4 VGND 0.11227f
C37392 vgaringosc.workerclkbuff_notouch_.I.n5 VGND 0.00969f
C37393 _324_.B.t4 VGND 0.01496f
C37394 _324_.B.t5 VGND 0.01496f
C37395 _324_.B.n0 VGND 0.03037f
C37396 _324_.B.t26 VGND 0.02828f
C37397 _324_.B.t20 VGND 0.052f
C37398 _324_.B.n1 VGND 0.05418f
C37399 _324_.B.t32 VGND 0.05411f
C37400 _324_.B.t21 VGND 0.0321f
C37401 _324_.B.n2 VGND 0.05654f
C37402 _324_.B.t27 VGND 0.04662f
C37403 _324_.B.t25 VGND 0.06251f
C37404 _324_.B.t28 VGND 0.02722f
C37405 _324_.B.n3 VGND 0.06847f
C37406 _324_.B.t30 VGND 0.02647f
C37407 _324_.B.n4 VGND 0.04671f
C37408 _324_.B.n5 VGND 0.04196f
C37409 _324_.B.n6 VGND 0.10555f
C37410 _324_.B.n7 VGND 0.32548f
C37411 _324_.B.n8 VGND 0.34462f
C37412 _324_.B.t22 VGND 0.04379f
C37413 _324_.B.t23 VGND 0.05011f
C37414 _324_.B.n9 VGND 0.06844f
C37415 _324_.B.t33 VGND 0.04544f
C37416 _324_.B.t31 VGND 0.05064f
C37417 _324_.B.n10 VGND 0.06073f
C37418 _324_.B.t24 VGND 0.04531f
C37419 _324_.B.t29 VGND 0.05078f
C37420 _324_.B.n11 VGND 0.05977f
C37421 _324_.B.n12 VGND 0.04473f
C37422 _324_.B.n13 VGND 0.35004f
C37423 _324_.B.n14 VGND 0.10571f
C37424 _324_.B.n15 VGND 0.10297f
C37425 _324_.B.t10 VGND 0.01496f
C37426 _324_.B.t11 VGND 0.01496f
C37427 _324_.B.n16 VGND 0.02991f
C37428 _324_.B.n17 VGND 0.0937f
C37429 _324_.B.t19 VGND 0.01345f
C37430 _324_.B.t12 VGND 0.01345f
C37431 _324_.B.n18 VGND 0.03254f
C37432 _324_.B.t14 VGND 0.01345f
C37433 _324_.B.t16 VGND 0.01345f
C37434 _324_.B.n19 VGND 0.02691f
C37435 _324_.B.n20 VGND 0.13397f
C37436 _324_.B.t18 VGND 0.01345f
C37437 _324_.B.t13 VGND 0.01345f
C37438 _324_.B.n21 VGND 0.02691f
C37439 _324_.B.n22 VGND 0.07905f
C37440 _324_.B.t15 VGND 0.01345f
C37441 _324_.B.t17 VGND 0.01345f
C37442 _324_.B.n23 VGND 0.02691f
C37443 _324_.B.n24 VGND 0.06308f
C37444 _324_.B.t1 VGND 0.02038f
C37445 _324_.B.t6 VGND 0.0061f
C37446 _324_.B.n25 VGND 0.04242f
C37447 _324_.B.t7 VGND 0.0112f
C37448 _324_.B.t3 VGND 0.0112f
C37449 _324_.B.n26 VGND 0.0224f
C37450 _324_.B.n27 VGND 0.0817f
C37451 _324_.B.t0 VGND 0.0112f
C37452 _324_.B.t8 VGND 0.0112f
C37453 _324_.B.n28 VGND 0.0224f
C37454 _324_.B.n29 VGND 0.05413f
C37455 _324_.B.t9 VGND 0.0061f
C37456 _324_.B.t2 VGND 0.02038f
C37457 _324_.B.n30 VGND 0.03858f
C37458 _324_.B.n31 VGND 0.06703f
C37459 _324_.B.n32 VGND 0.08688f
C37460 _402_.A1.t0 VGND 0.01602f
C37461 _402_.A1.t1 VGND 0.01602f
C37462 _402_.A1.n0 VGND 0.03236f
C37463 _402_.A1.t3 VGND 0.01077f
C37464 _402_.A1.t2 VGND 0.01077f
C37465 _402_.A1.n1 VGND 0.02578f
C37466 _402_.A1.t23 VGND 0.03372f
C37467 _402_.A1.t17 VGND 0.05795f
C37468 _402_.A1.n2 VGND 0.05875f
C37469 _402_.A1.t5 VGND 0.03532f
C37470 _402_.A1.t7 VGND 0.03687f
C37471 _402_.A1.n3 VGND 0.0682f
C37472 _402_.A1.t4 VGND 0.03962f
C37473 _402_.A1.t20 VGND 0.03687f
C37474 _402_.A1.n4 VGND 0.06856f
C37475 _402_.A1.n5 VGND 0.10021f
C37476 _402_.A1.t14 VGND 0.05f
C37477 _402_.A1.t13 VGND 0.02719f
C37478 _402_.A1.n6 VGND 0.05209f
C37479 _402_.A1.t18 VGND 0.04257f
C37480 _402_.A1.t12 VGND 0.04948f
C37481 _402_.A1.n7 VGND 0.04392f
C37482 _402_.A1.t8 VGND 0.03927f
C37483 _402_.A1.t9 VGND 0.05058f
C37484 _402_.A1.n8 VGND 0.05787f
C37485 _402_.A1.n9 VGND 0.08598f
C37486 _402_.A1.n10 VGND 0.23759f
C37487 _402_.A1.n11 VGND 0.40449f
C37488 _402_.A1.t15 VGND 0.05025f
C37489 _402_.A1.t10 VGND 0.03909f
C37490 _402_.A1.n12 VGND 0.05666f
C37491 _402_.A1.n13 VGND 0.29031f
C37492 _402_.A1.t11 VGND 0.04161f
C37493 _402_.A1.t16 VGND 0.04811f
C37494 _402_.A1.n14 VGND 0.05604f
C37495 _402_.A1.n15 VGND 0.06015f
C37496 _402_.A1.n16 VGND 0.0928f
C37497 _402_.A1.t21 VGND 0.04869f
C37498 _402_.A1.t19 VGND 0.0447f
C37499 _402_.A1.n17 VGND 0.05642f
C37500 _402_.A1.n18 VGND 0.08739f
C37501 _402_.A1.t6 VGND 0.04106f
C37502 _402_.A1.t22 VGND 0.05046f
C37503 _402_.A1.n19 VGND 0.06482f
C37504 _402_.A1.n20 VGND 0.51836f
C37505 _402_.A1.n21 VGND 0.41343f
C37506 _402_.A1.n22 VGND 0.75184f
C37507 _474_.CLK.t30 VGND 0.0105f
C37508 _474_.CLK.t25 VGND 0.0105f
C37509 _474_.CLK.n0 VGND 0.02129f
C37510 _474_.CLK.t23 VGND 0.0105f
C37511 _474_.CLK.t19 VGND 0.0105f
C37512 _474_.CLK.n1 VGND 0.02129f
C37513 _474_.CLK.t14 VGND 0.0105f
C37514 _474_.CLK.t18 VGND 0.0105f
C37515 _474_.CLK.n2 VGND 0.02129f
C37516 _474_.CLK.t13 VGND 0.0105f
C37517 _474_.CLK.t10 VGND 0.0105f
C37518 _474_.CLK.n3 VGND 0.02892f
C37519 _474_.CLK.n4 VGND 0.21723f
C37520 _474_.CLK.n5 VGND 0.13922f
C37521 _474_.CLK.n6 VGND 0.09671f
C37522 _474_.CLK.t7 VGND 0.0105f
C37523 _474_.CLK.t27 VGND 0.0105f
C37524 _474_.CLK.n7 VGND 0.02129f
C37525 _474_.CLK.t8 VGND 0.0105f
C37526 _474_.CLK.t2 VGND 0.0105f
C37527 _474_.CLK.n8 VGND 0.02129f
C37528 _474_.CLK.t21 VGND 0.0105f
C37529 _474_.CLK.t12 VGND 0.0105f
C37530 _474_.CLK.n9 VGND 0.02129f
C37531 _474_.CLK.t17 VGND 0.0105f
C37532 _474_.CLK.t22 VGND 0.0105f
C37533 _474_.CLK.n10 VGND 0.02892f
C37534 _474_.CLK.n11 VGND 0.21723f
C37535 _474_.CLK.n12 VGND 0.13922f
C37536 _474_.CLK.n13 VGND 0.09805f
C37537 _474_.CLK.n14 VGND 0.10354f
C37538 _474_.CLK.t3 VGND 0.03658f
C37539 _474_.CLK.t9 VGND 0.02642f
C37540 _474_.CLK.n15 VGND 0.06303f
C37541 _474_.CLK.t53 VGND 0.05184f
C37542 _474_.CLK.t39 VGND 0.04824f
C37543 _474_.CLK.n16 VGND 0.07631f
C37544 _474_.CLK.n17 VGND 0.04486f
C37545 _474_.CLK.t35 VGND 0.04846f
C37546 _474_.CLK.t47 VGND 0.05163f
C37547 _474_.CLK.n18 VGND 0.07638f
C37548 _474_.CLK.n19 VGND 0.79265f
C37549 _474_.CLK.t37 VGND 0.04846f
C37550 _474_.CLK.t33 VGND 0.05163f
C37551 _474_.CLK.n20 VGND 0.0763f
C37552 _474_.CLK.n21 VGND 0.09093f
C37553 _474_.CLK.n22 VGND 1.01423f
C37554 _474_.CLK.t36 VGND 0.05184f
C37555 _474_.CLK.t43 VGND 0.04824f
C37556 _474_.CLK.n23 VGND 0.07631f
C37557 _474_.CLK.n24 VGND 0.04486f
C37558 _474_.CLK.n25 VGND 0.5471f
C37559 _474_.CLK.t54 VGND 0.08578f
C37560 _474_.CLK.t40 VGND 0.05089f
C37561 _474_.CLK.n26 VGND 0.0906f
C37562 _474_.CLK.n27 VGND 0.18911f
C37563 _474_.CLK.t38 VGND 0.08245f
C37564 _474_.CLK.t45 VGND 0.04484f
C37565 _474_.CLK.n28 VGND 0.08558f
C37566 _474_.CLK.n29 VGND 0.06187f
C37567 _474_.CLK.n30 VGND 0.68494f
C37568 _474_.CLK.t49 VGND 0.04846f
C37569 _474_.CLK.t48 VGND 0.05163f
C37570 _474_.CLK.n31 VGND 0.07638f
C37571 _474_.CLK.t55 VGND 0.05184f
C37572 _474_.CLK.t34 VGND 0.04824f
C37573 _474_.CLK.n32 VGND 0.07639f
C37574 _474_.CLK.t32 VGND 0.09813f
C37575 _474_.CLK.t56 VGND 0.05347f
C37576 _474_.CLK.t44 VGND 0.06944f
C37577 _474_.CLK.n33 VGND 0.10996f
C37578 _474_.CLK.n34 VGND 0.07299f
C37579 _474_.CLK.n35 VGND 0.89527f
C37580 _474_.CLK.n36 VGND 0.73366f
C37581 _474_.CLK.t42 VGND 0.04846f
C37582 _474_.CLK.t41 VGND 0.05163f
C37583 _474_.CLK.n37 VGND 0.07638f
C37584 _474_.CLK.n38 VGND 0.52492f
C37585 _474_.CLK.t52 VGND 0.05111f
C37586 _474_.CLK.t51 VGND 0.08578f
C37587 _474_.CLK.n39 VGND 0.09102f
C37588 _474_.CLK.n40 VGND 0.06533f
C37589 _474_.CLK.n41 VGND 0.47775f
C37590 _474_.CLK.n42 VGND 0.70183f
C37591 _474_.CLK.t46 VGND 0.05184f
C37592 _474_.CLK.t50 VGND 0.04824f
C37593 _474_.CLK.n43 VGND 0.07631f
C37594 _474_.CLK.n44 VGND 0.04486f
C37595 _474_.CLK.n45 VGND 0.69143f
C37596 _474_.CLK.n46 VGND 0.66652f
C37597 _474_.CLK.n47 VGND 0.14755f
C37598 _474_.CLK.t6 VGND 0.03658f
C37599 _474_.CLK.t31 VGND 0.02642f
C37600 _474_.CLK.n48 VGND 0.06299f
C37601 _474_.CLK.n49 VGND 0.19373f
C37602 _474_.CLK.t28 VGND 0.03658f
C37603 _474_.CLK.t24 VGND 0.02642f
C37604 _474_.CLK.n50 VGND 0.06299f
C37605 _474_.CLK.n51 VGND 0.20145f
C37606 _474_.CLK.t26 VGND 0.03658f
C37607 _474_.CLK.t16 VGND 0.02642f
C37608 _474_.CLK.n52 VGND 0.06299f
C37609 _474_.CLK.n53 VGND 0.122f
C37610 _474_.CLK.t0 VGND 0.02642f
C37611 _474_.CLK.t29 VGND 0.03658f
C37612 _474_.CLK.n54 VGND 0.07427f
C37613 _474_.CLK.t1 VGND 0.03658f
C37614 _474_.CLK.t4 VGND 0.02642f
C37615 _474_.CLK.n55 VGND 0.06299f
C37616 _474_.CLK.n56 VGND 0.28489f
C37617 _474_.CLK.t11 VGND 0.03658f
C37618 _474_.CLK.t5 VGND 0.02642f
C37619 _474_.CLK.n57 VGND 0.06299f
C37620 _474_.CLK.n58 VGND 0.20145f
C37621 _474_.CLK.t20 VGND 0.03658f
C37622 _474_.CLK.t15 VGND 0.02642f
C37623 _474_.CLK.n59 VGND 0.06299f
C37624 _474_.CLK.n60 VGND 0.12924f
C37625 _474_.CLK.n61 VGND 0.16441f
C37626 _268_.A1.t0 VGND 0.04954f
C37627 _268_.A1.t9 VGND 0.03572f
C37628 _268_.A1.t7 VGND 0.05994f
C37629 _268_.A1.n0 VGND 0.06315f
C37630 _268_.A1.n1 VGND 0.04972f
C37631 _268_.A1.t4 VGND 0.05493f
C37632 _268_.A1.t5 VGND 0.05133f
C37633 _268_.A1.n2 VGND 0.07391f
C37634 _268_.A1.n3 VGND 0.02055f
C37635 _268_.A1.t3 VGND 0.05325f
C37636 _268_.A1.t8 VGND 0.03975f
C37637 _268_.A1.n4 VGND 0.06577f
C37638 _268_.A1.n5 VGND 0.08678f
C37639 _268_.A1.n6 VGND 0.16666f
C37640 _268_.A1.n7 VGND 0.12752f
C37641 _268_.A1.t6 VGND 0.03445f
C37642 _268_.A1.t2 VGND 0.04306f
C37643 _268_.A1.n8 VGND 0.06838f
C37644 _268_.A1.n9 VGND 0.49979f
C37645 _268_.A1.t1 VGND 0.0185f
C37646 _268_.A1.n10 VGND 0.14937f
C37647 _287_.A1.t1 VGND 0.03408f
C37648 _287_.A1.t2 VGND 0.02461f
C37649 _287_.A1.n0 VGND 0.06382f
C37650 _287_.A1.t6 VGND 0.00918f
C37651 _287_.A1.t7 VGND 0.00918f
C37652 _287_.A1.n1 VGND 0.0187f
C37653 _287_.A1.t4 VGND 0.00918f
C37654 _287_.A1.t5 VGND 0.00918f
C37655 _287_.A1.n2 VGND 0.02644f
C37656 _287_.A1.n3 VGND 0.13679f
C37657 _287_.A1.t38 VGND 0.06938f
C37658 _287_.A1.n4 VGND 0.0455f
C37659 _287_.A1.t19 VGND 0.06938f
C37660 _287_.A1.t8 VGND 0.06378f
C37661 _287_.A1.n5 VGND 0.07046f
C37662 _287_.A1.t33 VGND 0.06378f
C37663 _287_.A1.n6 VGND 0.07046f
C37664 _287_.A1.n7 VGND 0.04359f
C37665 _287_.A1.n8 VGND 0.0999f
C37666 _287_.A1.t10 VGND 0.06938f
C37667 _287_.A1.n9 VGND 0.04627f
C37668 _287_.A1.t21 VGND 0.06938f
C37669 _287_.A1.t24 VGND 0.06378f
C37670 _287_.A1.t28 VGND 0.06378f
C37671 _287_.A1.n10 VGND 0.07046f
C37672 _287_.A1.n11 VGND 0.07046f
C37673 _287_.A1.n12 VGND 0.04359f
C37674 _287_.A1.n13 VGND 0.13588f
C37675 _287_.A1.n14 VGND 0.32697f
C37676 _287_.A1.t25 VGND 0.06938f
C37677 _287_.A1.n15 VGND 0.04627f
C37678 _287_.A1.t26 VGND 0.06938f
C37679 _287_.A1.t23 VGND 0.06378f
C37680 _287_.A1.n16 VGND 0.07046f
C37681 _287_.A1.t20 VGND 0.06378f
C37682 _287_.A1.n17 VGND 0.07046f
C37683 _287_.A1.n18 VGND 0.04359f
C37684 _287_.A1.n19 VGND 0.12197f
C37685 _287_.A1.t18 VGND 0.06938f
C37686 _287_.A1.n20 VGND 0.0455f
C37687 _287_.A1.t17 VGND 0.06938f
C37688 _287_.A1.t11 VGND 0.06378f
C37689 _287_.A1.n21 VGND 0.07046f
C37690 _287_.A1.t15 VGND 0.06378f
C37691 _287_.A1.n22 VGND 0.07046f
C37692 _287_.A1.n23 VGND 0.04359f
C37693 _287_.A1.n24 VGND 0.11381f
C37694 _287_.A1.n25 VGND 0.06339f
C37695 _287_.A1.t30 VGND 0.06938f
C37696 _287_.A1.n26 VGND 0.0455f
C37697 _287_.A1.t39 VGND 0.06402f
C37698 _287_.A1.n27 VGND 0.07022f
C37699 _287_.A1.t37 VGND 0.06402f
C37700 _287_.A1.n28 VGND 0.07022f
C37701 _287_.A1.t13 VGND 0.06938f
C37702 _287_.A1.n29 VGND 0.04359f
C37703 _287_.A1.n30 VGND 0.11381f
C37704 _287_.A1.n31 VGND 0.073f
C37705 _287_.A1.t22 VGND 0.06402f
C37706 _287_.A1.t14 VGND 0.06938f
C37707 _287_.A1.n32 VGND 0.04359f
C37708 _287_.A1.n33 VGND 0.07022f
C37709 _287_.A1.t29 VGND 0.06402f
C37710 _287_.A1.n34 VGND 0.07022f
C37711 _287_.A1.t35 VGND 0.06938f
C37712 _287_.A1.n35 VGND 0.04359f
C37713 _287_.A1.n36 VGND 0.06491f
C37714 _287_.A1.n37 VGND 0.1906f
C37715 _287_.A1.n38 VGND 0.77977f
C37716 _287_.A1.t32 VGND 0.06938f
C37717 _287_.A1.n39 VGND 0.0455f
C37718 _287_.A1.t12 VGND 0.06402f
C37719 _287_.A1.n40 VGND 0.07022f
C37720 _287_.A1.t9 VGND 0.06402f
C37721 _287_.A1.n41 VGND 0.07022f
C37722 _287_.A1.t16 VGND 0.06938f
C37723 _287_.A1.n42 VGND 0.04359f
C37724 _287_.A1.n43 VGND 0.11381f
C37725 _287_.A1.t36 VGND 0.06938f
C37726 _287_.A1.n44 VGND 0.04627f
C37727 _287_.A1.t34 VGND 0.06402f
C37728 _287_.A1.t31 VGND 0.06402f
C37729 _287_.A1.n45 VGND 0.07022f
C37730 _287_.A1.n46 VGND 0.07022f
C37731 _287_.A1.t27 VGND 0.06938f
C37732 _287_.A1.n47 VGND 0.04359f
C37733 _287_.A1.n48 VGND 0.12197f
C37734 _287_.A1.n49 VGND 0.05426f
C37735 _287_.A1.n50 VGND 0.67945f
C37736 _287_.A1.n51 VGND 0.09154f
C37737 _287_.A1.t0 VGND 0.02461f
C37738 _287_.A1.t3 VGND 0.03408f
C37739 _287_.A1.n52 VGND 0.05931f
C37740 _287_.A1.n53 VGND 0.06645f
C37741 a_26916_25640.t7 VGND 0.04128f
C37742 a_26916_25640.t6 VGND 0.13823f
C37743 a_26916_25640.t2 VGND 0.12194f
C37744 a_26916_25640.n0 VGND 0.15796f
C37745 a_26916_25640.n1 VGND 0.05384f
C37746 a_26916_25640.t1 VGND 0.04561f
C37747 a_26916_25640.n2 VGND 0.20374f
C37748 a_26916_25640.t5 VGND 0.01944f
C37749 a_26916_25640.t4 VGND 0.12223f
C37750 a_26916_25640.t3 VGND 0.38419f
C37751 a_26916_25640.n3 VGND 0.24674f
C37752 a_26916_25640.n4 VGND 0.56455f
C37753 a_26916_25640.t0 VGND 0.10024f
C37754 _359_.B.t0 VGND 0.09387f
C37755 _359_.B.t1 VGND 0.06617f
C37756 _359_.B.t2 VGND 0.08836f
C37757 _359_.B.t9 VGND 0.10089f
C37758 _359_.B.n0 VGND 0.12594f
C37759 _359_.B.n1 VGND 0.23882f
C37760 _359_.B.t5 VGND 0.07679f
C37761 _359_.B.t11 VGND 0.09197f
C37762 _359_.B.n2 VGND 0.11718f
C37763 _359_.B.n3 VGND 0.19591f
C37764 _359_.B.n4 VGND 0.96547f
C37765 _359_.B.t10 VGND 0.07088f
C37766 _359_.B.t3 VGND 0.09456f
C37767 _359_.B.n5 VGND 0.11735f
C37768 _359_.B.n6 VGND 0.82294f
C37769 _359_.B.t6 VGND 0.09197f
C37770 _359_.B.t4 VGND 0.09011f
C37771 _359_.B.n7 VGND 0.12443f
C37772 _359_.B.n8 VGND 0.66846f
C37773 _359_.B.n9 VGND 1.14201f
C37774 _359_.B.t8 VGND 0.10644f
C37775 _359_.B.t7 VGND 0.06315f
C37776 _359_.B.n10 VGND 0.11123f
C37777 _359_.B.n11 VGND 2.34669f
C37778 _324_.C.t5 VGND 0.01002f
C37779 _324_.C.t6 VGND 0.01002f
C37780 _324_.C.n0 VGND 0.02041f
C37781 _324_.C.t4 VGND 0.01002f
C37782 _324_.C.t7 VGND 0.01002f
C37783 _324_.C.n1 VGND 0.02886f
C37784 _324_.C.n2 VGND 0.1737f
C37785 _324_.C.t2 VGND 0.0372f
C37786 _324_.C.t3 VGND 0.02687f
C37787 _324_.C.n3 VGND 0.06473f
C37788 _324_.C.n4 VGND 0.09569f
C37789 _324_.C.t1 VGND 0.02687f
C37790 _324_.C.t0 VGND 0.0372f
C37791 _324_.C.n5 VGND 0.06537f
C37792 _324_.C.t19 VGND 0.0808f
C37793 _324_.C.t26 VGND 0.0704f
C37794 _324_.C.n6 VGND 0.11215f
C37795 _324_.C.t8 VGND 0.05574f
C37796 _324_.C.t23 VGND 0.09528f
C37797 _324_.C.n7 VGND 0.10009f
C37798 _324_.C.t30 VGND 0.05574f
C37799 _324_.C.t14 VGND 0.09528f
C37800 _324_.C.n8 VGND 0.10006f
C37801 _324_.C.n9 VGND 0.04954f
C37802 _324_.C.n10 VGND 0.89677f
C37803 _324_.C.t13 VGND 0.04955f
C37804 _324_.C.t31 VGND 0.07936f
C37805 _324_.C.n11 VGND 0.11238f
C37806 _324_.C.t9 VGND 0.04955f
C37807 _324_.C.t27 VGND 0.07936f
C37808 _324_.C.n12 VGND 0.1008f
C37809 _324_.C.n13 VGND 0.01556f
C37810 _324_.C.t29 VGND 0.08427f
C37811 _324_.C.t22 VGND 0.06555f
C37812 _324_.C.n14 VGND 0.09501f
C37813 _324_.C.n15 VGND 0.89737f
C37814 _324_.C.t18 VGND 0.08427f
C37815 _324_.C.t32 VGND 0.06555f
C37816 _324_.C.n16 VGND 0.09501f
C37817 _324_.C.t15 VGND 0.09528f
C37818 _324_.C.t21 VGND 0.05574f
C37819 _324_.C.n17 VGND 0.10103f
C37820 _324_.C.t28 VGND 0.09528f
C37821 _324_.C.t16 VGND 0.05574f
C37822 _324_.C.n18 VGND 0.10006f
C37823 _324_.C.t24 VGND 0.07061f
C37824 _324_.C.t11 VGND 0.0808f
C37825 _324_.C.n19 VGND 0.11227f
C37826 _324_.C.n20 VGND 0.81617f
C37827 _324_.C.t12 VGND 0.06886f
C37828 _324_.C.t20 VGND 0.08268f
C37829 _324_.C.n21 VGND 0.11017f
C37830 _324_.C.n22 VGND 0.11257f
C37831 _324_.C.n23 VGND 1.04391f
C37832 _324_.C.n24 VGND 0.50465f
C37833 _324_.C.n25 VGND 0.94464f
C37834 _324_.C.n26 VGND 1.04313f
C37835 _324_.C.t17 VGND 0.06555f
C37836 _324_.C.t33 VGND 0.08427f
C37837 _324_.C.n27 VGND 0.09502f
C37838 _324_.C.n28 VGND 1.81992f
C37839 _324_.C.t25 VGND 0.04797f
C37840 _324_.C.t10 VGND 0.06119f
C37841 _324_.C.n29 VGND 0.10057f
C37842 _324_.C.n30 VGND 2.06113f
C37843 _324_.C.n31 VGND 0.47221f
C37844 _304_.ZN.t9 VGND 0.00686f
C37845 _304_.ZN.t0 VGND 0.02292f
C37846 _304_.ZN.n0 VGND 0.04772f
C37847 _304_.ZN.t6 VGND 0.0126f
C37848 _304_.ZN.t5 VGND 0.0126f
C37849 _304_.ZN.n1 VGND 0.0252f
C37850 _304_.ZN.n2 VGND 0.09191f
C37851 _304_.ZN.t1 VGND 0.02292f
C37852 _304_.ZN.t8 VGND 0.00686f
C37853 _304_.ZN.n3 VGND 0.0434f
C37854 _304_.ZN.n4 VGND 0.05147f
C37855 _304_.ZN.t15 VGND 0.04939f
C37856 _304_.ZN.n5 VGND 0.03767f
C37857 _304_.ZN.t11 VGND 0.04939f
C37858 _304_.ZN.n6 VGND 0.03872f
C37859 _304_.ZN.t17 VGND 0.05301f
C37860 _304_.ZN.n7 VGND 0.0513f
C37861 _304_.ZN.t13 VGND 0.05301f
C37862 _304_.ZN.n8 VGND 0.0513f
C37863 _304_.ZN.t16 VGND 0.04939f
C37864 _304_.ZN.n9 VGND 0.03759f
C37865 _304_.ZN.n10 VGND 0.08378f
C37866 _304_.ZN.t10 VGND 0.05301f
C37867 _304_.ZN.n11 VGND 0.0513f
C37868 _304_.ZN.t12 VGND 0.05301f
C37869 _304_.ZN.n12 VGND 0.0513f
C37870 _304_.ZN.t14 VGND 0.04939f
C37871 _304_.ZN.n13 VGND 0.03759f
C37872 _304_.ZN.n14 VGND 0.04236f
C37873 _304_.ZN.n15 VGND 0.18752f
C37874 _304_.ZN.n16 VGND 0.19308f
C37875 _304_.ZN.t4 VGND 0.01682f
C37876 _304_.ZN.t7 VGND 0.01682f
C37877 _304_.ZN.n17 VGND 0.04694f
C37878 _304_.ZN.t2 VGND 0.01659f
C37879 _304_.ZN.t3 VGND 0.01659f
C37880 _304_.ZN.n18 VGND 0.03718f
C37881 _304_.ZN.n19 VGND 0.15007f
C37882 clkbuf_1_0__f_clk.I.t13 VGND 0.06811f
C37883 clkbuf_1_0__f_clk.I.t0 VGND 0.04919f
C37884 clkbuf_1_0__f_clk.I.n0 VGND 0.1383f
C37885 clkbuf_1_0__f_clk.I.t14 VGND 0.04919f
C37886 clkbuf_1_0__f_clk.I.t1 VGND 0.06811f
C37887 clkbuf_1_0__f_clk.I.n1 VGND 0.11731f
C37888 clkbuf_1_0__f_clk.I.n2 VGND 0.41539f
C37889 clkbuf_1_0__f_clk.I.t56 VGND 0.18777f
C37890 clkbuf_1_0__f_clk.I.t53 VGND 0.07258f
C37891 clkbuf_1_0__f_clk.I.t59 VGND 0.12971f
C37892 clkbuf_1_0__f_clk.I.n3 VGND 0.3546f
C37893 clkbuf_1_0__f_clk.I.t38 VGND 0.07258f
C37894 clkbuf_1_0__f_clk.I.t48 VGND 0.12971f
C37895 clkbuf_1_0__f_clk.I.n4 VGND 0.25202f
C37896 clkbuf_1_0__f_clk.I.t43 VGND 0.07258f
C37897 clkbuf_1_0__f_clk.I.t51 VGND 0.12971f
C37898 clkbuf_1_0__f_clk.I.n5 VGND 0.25202f
C37899 clkbuf_1_0__f_clk.I.t33 VGND 0.19653f
C37900 clkbuf_1_0__f_clk.I.t58 VGND 0.07258f
C37901 clkbuf_1_0__f_clk.I.t40 VGND 0.12971f
C37902 clkbuf_1_0__f_clk.I.n6 VGND 0.35701f
C37903 clkbuf_1_0__f_clk.I.t37 VGND 0.07258f
C37904 clkbuf_1_0__f_clk.I.t46 VGND 0.12971f
C37905 clkbuf_1_0__f_clk.I.n7 VGND 0.25202f
C37906 clkbuf_1_0__f_clk.I.t42 VGND 0.07258f
C37907 clkbuf_1_0__f_clk.I.t50 VGND 0.12971f
C37908 clkbuf_1_0__f_clk.I.n8 VGND 0.2995f
C37909 clkbuf_1_0__f_clk.I.t47 VGND 0.19653f
C37910 clkbuf_1_0__f_clk.I.t41 VGND 0.12971f
C37911 clkbuf_1_0__f_clk.I.t49 VGND 0.07211f
C37912 clkbuf_1_0__f_clk.I.n9 VGND 0.35748f
C37913 clkbuf_1_0__f_clk.I.t34 VGND 0.12971f
C37914 clkbuf_1_0__f_clk.I.t45 VGND 0.07211f
C37915 clkbuf_1_0__f_clk.I.n10 VGND 0.25249f
C37916 clkbuf_1_0__f_clk.I.t54 VGND 0.18777f
C37917 clkbuf_1_0__f_clk.I.t57 VGND 0.12971f
C37918 clkbuf_1_0__f_clk.I.t35 VGND 0.07211f
C37919 clkbuf_1_0__f_clk.I.n11 VGND 0.35507f
C37920 clkbuf_1_0__f_clk.I.t55 VGND 0.12971f
C37921 clkbuf_1_0__f_clk.I.t32 VGND 0.07211f
C37922 clkbuf_1_0__f_clk.I.n12 VGND 0.25249f
C37923 clkbuf_1_0__f_clk.I.t39 VGND 0.12971f
C37924 clkbuf_1_0__f_clk.I.t36 VGND 0.07211f
C37925 clkbuf_1_0__f_clk.I.n13 VGND 0.25249f
C37926 clkbuf_1_0__f_clk.I.t44 VGND 0.12971f
C37927 clkbuf_1_0__f_clk.I.t52 VGND 0.07211f
C37928 clkbuf_1_0__f_clk.I.n14 VGND 0.29997f
C37929 clkbuf_1_0__f_clk.I.n15 VGND 1.25521f
C37930 clkbuf_1_0__f_clk.I.n16 VGND 0.19795f
C37931 clkbuf_1_0__f_clk.I.t7 VGND 0.04919f
C37932 clkbuf_1_0__f_clk.I.t5 VGND 0.06811f
C37933 clkbuf_1_0__f_clk.I.n17 VGND 0.11731f
C37934 clkbuf_1_0__f_clk.I.n18 VGND 0.2888f
C37935 clkbuf_1_0__f_clk.I.t8 VGND 0.04919f
C37936 clkbuf_1_0__f_clk.I.t6 VGND 0.06811f
C37937 clkbuf_1_0__f_clk.I.n19 VGND 0.11731f
C37938 clkbuf_1_0__f_clk.I.n20 VGND 0.24068f
C37939 clkbuf_1_0__f_clk.I.t4 VGND 0.04919f
C37940 clkbuf_1_0__f_clk.I.t3 VGND 0.06811f
C37941 clkbuf_1_0__f_clk.I.n21 VGND 0.14023f
C37942 clkbuf_1_0__f_clk.I.t15 VGND 0.04919f
C37943 clkbuf_1_0__f_clk.I.t2 VGND 0.06811f
C37944 clkbuf_1_0__f_clk.I.n22 VGND 0.11731f
C37945 clkbuf_1_0__f_clk.I.n23 VGND 0.54659f
C37946 clkbuf_1_0__f_clk.I.t10 VGND 0.04919f
C37947 clkbuf_1_0__f_clk.I.t12 VGND 0.06811f
C37948 clkbuf_1_0__f_clk.I.n24 VGND 0.11731f
C37949 clkbuf_1_0__f_clk.I.n25 VGND 0.37515f
C37950 clkbuf_1_0__f_clk.I.t9 VGND 0.04919f
C37951 clkbuf_1_0__f_clk.I.t11 VGND 0.06811f
C37952 clkbuf_1_0__f_clk.I.n26 VGND 0.11731f
C37953 clkbuf_1_0__f_clk.I.n27 VGND 0.22719f
C37954 clkbuf_1_0__f_clk.I.n28 VGND 0.30617f
C37955 clkbuf_1_0__f_clk.I.t29 VGND 0.01956f
C37956 clkbuf_1_0__f_clk.I.t31 VGND 0.01956f
C37957 clkbuf_1_0__f_clk.I.n29 VGND 0.03964f
C37958 clkbuf_1_0__f_clk.I.t30 VGND 0.01956f
C37959 clkbuf_1_0__f_clk.I.t21 VGND 0.01956f
C37960 clkbuf_1_0__f_clk.I.n30 VGND 0.03964f
C37961 clkbuf_1_0__f_clk.I.t18 VGND 0.01956f
C37962 clkbuf_1_0__f_clk.I.t20 VGND 0.01956f
C37963 clkbuf_1_0__f_clk.I.n31 VGND 0.03964f
C37964 clkbuf_1_0__f_clk.I.t22 VGND 0.01956f
C37965 clkbuf_1_0__f_clk.I.t27 VGND 0.01956f
C37966 clkbuf_1_0__f_clk.I.n32 VGND 0.05386f
C37967 clkbuf_1_0__f_clk.I.n33 VGND 0.40454f
C37968 clkbuf_1_0__f_clk.I.n34 VGND 0.25926f
C37969 clkbuf_1_0__f_clk.I.n35 VGND 0.18258f
C37970 clkbuf_1_0__f_clk.I.t26 VGND 0.01956f
C37971 clkbuf_1_0__f_clk.I.t28 VGND 0.01956f
C37972 clkbuf_1_0__f_clk.I.n36 VGND 0.03964f
C37973 clkbuf_1_0__f_clk.I.t25 VGND 0.01956f
C37974 clkbuf_1_0__f_clk.I.t24 VGND 0.01956f
C37975 clkbuf_1_0__f_clk.I.n37 VGND 0.03964f
C37976 clkbuf_1_0__f_clk.I.t17 VGND 0.01956f
C37977 clkbuf_1_0__f_clk.I.t23 VGND 0.01956f
C37978 clkbuf_1_0__f_clk.I.n38 VGND 0.03964f
C37979 clkbuf_1_0__f_clk.I.t16 VGND 0.01956f
C37980 clkbuf_1_0__f_clk.I.t19 VGND 0.01956f
C37981 clkbuf_1_0__f_clk.I.n39 VGND 0.05386f
C37982 clkbuf_1_0__f_clk.I.n40 VGND 0.40454f
C37983 clkbuf_1_0__f_clk.I.n41 VGND 0.25926f
C37984 clkbuf_1_0__f_clk.I.n42 VGND 0.1801f
C37985 clkbuf_1_0__f_clk.I.n43 VGND 0.19282f
C37986 a_44296_24393.t12 VGND 0.04219f
C37987 a_44296_24393.t7 VGND 0.04219f
C37988 a_44296_24393.t13 VGND 0.05842f
C37989 a_44296_24393.n0 VGND 0.10181f
C37990 a_44296_24393.t5 VGND 0.04219f
C37991 a_44296_24393.t4 VGND 0.05842f
C37992 a_44296_24393.n1 VGND 0.10181f
C37993 a_44296_24393.t11 VGND 0.04219f
C37994 a_44296_24393.t2 VGND 0.05842f
C37995 a_44296_24393.n2 VGND 0.12544f
C37996 a_44296_24393.n3 VGND 0.40497f
C37997 a_44296_24393.n4 VGND 0.26004f
C37998 a_44296_24393.t1 VGND 0.05178f
C37999 a_44296_24393.t6 VGND 0.02084f
C38000 a_44296_24393.t3 VGND 0.02084f
C38001 a_44296_24393.n5 VGND 0.04236f
C38002 a_44296_24393.t10 VGND 0.02084f
C38003 a_44296_24393.t9 VGND 0.02084f
C38004 a_44296_24393.n6 VGND 0.04236f
C38005 a_44296_24393.t8 VGND 0.06562f
C38006 a_44296_24393.n7 VGND 0.41703f
C38007 a_44296_24393.n8 VGND 0.25146f
C38008 a_44296_24393.n9 VGND 0.20883f
C38009 a_44296_24393.t16 VGND 0.18298f
C38010 a_44296_24393.t45 VGND 0.12051f
C38011 a_44296_24393.n10 VGND 0.26983f
C38012 a_44296_24393.t42 VGND 0.18298f
C38013 a_44296_24393.t39 VGND 0.12051f
C38014 a_44296_24393.n11 VGND 0.30687f
C38015 a_44296_24393.t15 VGND 0.18298f
C38016 a_44296_24393.t44 VGND 0.12051f
C38017 a_44296_24393.n12 VGND 0.30687f
C38018 a_44296_24393.t29 VGND 0.18298f
C38019 a_44296_24393.t38 VGND 0.18298f
C38020 a_44296_24393.t25 VGND 0.12051f
C38021 a_44296_24393.n13 VGND 0.26983f
C38022 a_44296_24393.t36 VGND 0.18298f
C38023 a_44296_24393.t34 VGND 0.12051f
C38024 a_44296_24393.n14 VGND 0.30687f
C38025 a_44296_24393.t40 VGND 0.18298f
C38026 a_44296_24393.t37 VGND 0.12051f
C38027 a_44296_24393.n15 VGND 0.30687f
C38028 a_44296_24393.t14 VGND 0.18298f
C38029 a_44296_24393.t43 VGND 0.12051f
C38030 a_44296_24393.n16 VGND -0.57412f
C38031 a_44296_24393.t18 VGND 0.18298f
C38032 a_44296_24393.t35 VGND 0.12051f
C38033 a_44296_24393.n17 VGND 0.30687f
C38034 a_44296_24393.t23 VGND 0.18298f
C38035 a_44296_24393.t20 VGND 0.12051f
C38036 a_44296_24393.n18 VGND 0.30687f
C38037 a_44296_24393.t19 VGND 0.18298f
C38038 a_44296_24393.t17 VGND 0.12051f
C38039 a_44296_24393.n19 VGND 0.30687f
C38040 a_44296_24393.t24 VGND 0.18298f
C38041 a_44296_24393.t21 VGND 0.12051f
C38042 a_44296_24393.n20 VGND 0.30687f
C38043 a_44296_24393.t32 VGND 0.18298f
C38044 a_44296_24393.t22 VGND 0.12051f
C38045 a_44296_24393.n21 VGND 0.30687f
C38046 a_44296_24393.t28 VGND 0.18298f
C38047 a_44296_24393.t26 VGND 0.12051f
C38048 a_44296_24393.n22 VGND 0.30687f
C38049 a_44296_24393.t33 VGND 0.18298f
C38050 a_44296_24393.n23 VGND 0.15465f
C38051 a_44296_24393.t30 VGND 0.11992f
C38052 a_44296_24393.n24 VGND 0.15384f
C38053 a_44296_24393.t27 VGND 0.11992f
C38054 a_44296_24393.n25 VGND 0.15384f
C38055 a_44296_24393.n26 VGND 0.15465f
C38056 a_44296_24393.t41 VGND 0.18298f
C38057 a_44296_24393.t31 VGND 0.12051f
C38058 a_44296_24393.n27 VGND 0.83892f
C38059 a_44296_24393.n28 VGND 0.58145f
C38060 a_44296_24393.n29 VGND 0.21258f
C38061 a_44296_24393.n30 VGND 0.10181f
C38062 a_44296_24393.t0 VGND 0.05842f
C38063 VPWR.t759 VGND 0.00433f
C38064 VPWR.n0 VGND 0.01144f
C38065 VPWR.n1 VGND 0.05372f
C38066 VPWR.t4295 VGND 0.00433f
C38067 VPWR.t2315 VGND 0.00433f
C38068 VPWR.n2 VGND 0.01724f
C38069 VPWR.n3 VGND 0.58789f
C38070 VPWR.n4 VGND 0.00941f
C38071 VPWR.t4811 VGND 0.00433f
C38072 VPWR.t2817 VGND 0.00433f
C38073 VPWR.t3812 VGND 0.00433f
C38074 VPWR.t749 VGND 0.00433f
C38075 VPWR.t2006 VGND 0.00433f
C38076 VPWR.t380 VGND 0.00433f
C38077 VPWR.t3487 VGND 0.00433f
C38078 VPWR.t4536 VGND 0.00433f
C38079 VPWR.n5 VGND 0.03832f
C38080 VPWR.t2334 VGND 0.00433f
C38081 VPWR.t3328 VGND 0.00433f
C38082 VPWR.t2266 VGND 0.00433f
C38083 VPWR.t3276 VGND 0.00433f
C38084 VPWR.t597 VGND 0.00433f
C38085 VPWR.t4345 VGND 0.00433f
C38086 VPWR.t5793 VGND 0.00433f
C38087 VPWR.t2155 VGND 0.00433f
C38088 VPWR.t2333 VGND 0.05247f
C38089 VPWR.t3327 VGND 0.05996f
C38090 VPWR.t2265 VGND 0.05996f
C38091 VPWR.t3275 VGND 0.05996f
C38092 VPWR.t596 VGND 0.05996f
C38093 VPWR.t4344 VGND 0.05996f
C38094 VPWR.t5792 VGND 0.05996f
C38095 VPWR.t2154 VGND 0.04035f
C38096 VPWR.n6 VGND 0.03832f
C38097 VPWR.t4947 VGND 0.00433f
C38098 VPWR.n7 VGND 0.01089f
C38099 VPWR.n8 VGND 0.78236f
C38100 VPWR.n9 VGND 0.01186f
C38101 VPWR.t2038 VGND 0.00433f
C38102 VPWR.t6091 VGND 0.00433f
C38103 VPWR.t6432 VGND 0.00433f
C38104 VPWR.t5746 VGND 0.00433f
C38105 VPWR.t7139 VGND 0.00433f
C38106 VPWR.t5472 VGND 0.00433f
C38107 VPWR.t4027 VGND 0.00433f
C38108 VPWR.t6257 VGND 0.00433f
C38109 VPWR.t5697 VGND 0.00433f
C38110 VPWR.t1303 VGND 0.00433f
C38111 VPWR.t1662 VGND 0.00433f
C38112 VPWR.t1805 VGND 0.00433f
C38113 VPWR.t6295 VGND 0.00433f
C38114 VPWR.t2093 VGND 0.0202f
C38115 VPWR.t2094 VGND 0.00433f
C38116 VPWR.t3259 VGND 0.00433f
C38117 VPWR.t1174 VGND 0.00433f
C38118 VPWR.t2314 VGND 0.08751f
C38119 VPWR.t912 VGND 0.10001f
C38120 VPWR.t673 VGND 0.10001f
C38121 VPWR.t4300 VGND 0.10001f
C38122 VPWR.t1702 VGND 0.10001f
C38123 VPWR.t574 VGND 0.06731f
C38124 VPWR.t3258 VGND 0.025f
C38125 VPWR.t1173 VGND 0.04231f
C38126 VPWR.t3936 VGND 0.03751f
C38127 VPWR.n10 VGND 0.03642f
C38128 VPWR.t3937 VGND 0.00433f
C38129 VPWR.t575 VGND 0.00433f
C38130 VPWR.t4855 VGND 0.00433f
C38131 VPWR.t1703 VGND 0.00433f
C38132 VPWR.t1714 VGND 0.00433f
C38133 VPWR.t4301 VGND 0.00433f
C38134 VPWR.t5683 VGND 0.00433f
C38135 VPWR.t674 VGND 0.00433f
C38136 VPWR.t1810 VGND 0.00433f
C38137 VPWR.t913 VGND 0.00433f
C38138 VPWR.t3426 VGND 0.00433f
C38139 VPWR.n11 VGND 0.02171f
C38140 VPWR.n12 VGND 0.02171f
C38141 VPWR.n13 VGND 0.0207f
C38142 VPWR.n14 VGND 0.01577f
C38143 VPWR.n15 VGND 0.02171f
C38144 VPWR.n16 VGND 0.01144f
C38145 VPWR.n17 VGND 0.01189f
C38146 VPWR.n18 VGND 0.00912f
C38147 VPWR.n19 VGND 0.0085f
C38148 VPWR.n20 VGND 0.01144f
C38149 VPWR.t3441 VGND 0.00433f
C38150 VPWR.t1115 VGND 0.00433f
C38151 VPWR.t3857 VGND 0.00433f
C38152 VPWR.t1701 VGND 0.00433f
C38153 VPWR.t3563 VGND 0.00433f
C38154 VPWR.t1824 VGND 0.00433f
C38155 VPWR.t3832 VGND 0.00433f
C38156 VPWR.t2691 VGND 0.00433f
C38157 VPWR.t4756 VGND 0.00433f
C38158 VPWR.t4263 VGND 0.00433f
C38159 VPWR.t3692 VGND 0.00433f
C38160 VPWR.t5736 VGND 0.00433f
C38161 VPWR.t4099 VGND 0.00433f
C38162 VPWR.t3137 VGND 0.00433f
C38163 VPWR.t6009 VGND 0.00433f
C38164 VPWR.t5973 VGND 0.00433f
C38165 VPWR.t1878 VGND 0.00433f
C38166 VPWR.n21 VGND 0.01144f
C38167 VPWR.n22 VGND 0.01568f
C38168 VPWR.n23 VGND 0.02079f
C38169 VPWR.n24 VGND 0.02171f
C38170 VPWR.n25 VGND 0.01577f
C38171 VPWR.n26 VGND 0.0207f
C38172 VPWR.n27 VGND 0.02171f
C38173 VPWR.n28 VGND 0.02171f
C38174 VPWR.n29 VGND 0.01762f
C38175 VPWR.n30 VGND 0.01189f
C38176 VPWR.n31 VGND 0.05372f
C38177 VPWR.t1114 VGND 0.08751f
C38178 VPWR.t1700 VGND 0.10001f
C38179 VPWR.t1823 VGND 0.10001f
C38180 VPWR.t2690 VGND 0.10001f
C38181 VPWR.t4262 VGND 0.10001f
C38182 VPWR.t3691 VGND 0.10001f
C38183 VPWR.t3136 VGND 0.10001f
C38184 VPWR.t5972 VGND 0.06731f
C38185 VPWR.n32 VGND 0.03642f
C38186 VPWR.t1877 VGND 0.03751f
C38187 VPWR.t2037 VGND 0.05001f
C38188 VPWR.t6090 VGND 0.05001f
C38189 VPWR.t6431 VGND 0.05001f
C38190 VPWR.t5745 VGND 0.05001f
C38191 VPWR.t7138 VGND 0.05001f
C38192 VPWR.t5471 VGND 0.05001f
C38193 VPWR.t4026 VGND 0.05001f
C38194 VPWR.t6256 VGND 0.05001f
C38195 VPWR.t5696 VGND 0.05001f
C38196 VPWR.t1302 VGND 0.05001f
C38197 VPWR.t1661 VGND 0.05001f
C38198 VPWR.t1804 VGND 0.04231f
C38199 VPWR.t6294 VGND 0.0202f
C38200 VPWR.n33 VGND 0.05372f
C38201 VPWR.t4290 VGND 0.00433f
C38202 VPWR.t2973 VGND 0.00433f
C38203 VPWR.t6023 VGND 0.00433f
C38204 VPWR.t2972 VGND 0.05481f
C38205 VPWR.n34 VGND 0.03642f
C38206 VPWR.t957 VGND 0.00433f
C38207 VPWR.t3959 VGND 0.00433f
C38208 VPWR.t368 VGND 0.00433f
C38209 VPWR.t5458 VGND 0.00433f
C38210 VPWR.t3553 VGND 0.00433f
C38211 VPWR.t1870 VGND 0.00433f
C38212 VPWR.t5686 VGND 0.00433f
C38213 VPWR.t5103 VGND 0.00433f
C38214 VPWR.t5478 VGND 0.00433f
C38215 VPWR.t4216 VGND 0.00433f
C38216 VPWR.t6225 VGND 0.00433f
C38217 VPWR.t6267 VGND 0.00433f
C38218 VPWR.t1043 VGND 0.00433f
C38219 VPWR.t467 VGND 0.00433f
C38220 VPWR.t5364 VGND 0.00433f
C38221 VPWR.t519 VGND 0.00433f
C38222 VPWR.t6022 VGND 0.03751f
C38223 VPWR.t956 VGND 0.05001f
C38224 VPWR.t3958 VGND 0.05001f
C38225 VPWR.t367 VGND 0.05001f
C38226 VPWR.t5457 VGND 0.05001f
C38227 VPWR.t3552 VGND 0.05001f
C38228 VPWR.t1869 VGND 0.05001f
C38229 VPWR.t5685 VGND 0.05001f
C38230 VPWR.t5102 VGND 0.05001f
C38231 VPWR.t5477 VGND 0.05001f
C38232 VPWR.t4215 VGND 0.05001f
C38233 VPWR.t6224 VGND 0.05001f
C38234 VPWR.t6266 VGND 0.05001f
C38235 VPWR.t1042 VGND 0.05001f
C38236 VPWR.t466 VGND 0.05001f
C38237 VPWR.t5363 VGND 0.04231f
C38238 VPWR.t518 VGND 0.0202f
C38239 VPWR.n35 VGND 0.05372f
C38240 VPWR.t2043 VGND 0.00433f
C38241 VPWR.t4928 VGND 0.00433f
C38242 VPWR.t5982 VGND 0.00433f
C38243 VPWR.t4613 VGND 0.00433f
C38244 VPWR.n36 VGND 0.01929f
C38245 VPWR.n37 VGND 0.78236f
C38246 VPWR.t6119 VGND 0.00433f
C38247 VPWR.n38 VGND 0.00918f
C38248 VPWR.t3606 VGND 0.00433f
C38249 VPWR.t5267 VGND 0.00433f
C38250 VPWR.t5389 VGND 0.00433f
C38251 VPWR.t3779 VGND 0.00433f
C38252 VPWR.t1199 VGND 0.00433f
C38253 VPWR.t75 VGND 0.00433f
C38254 VPWR.t5651 VGND 0.00433f
C38255 VPWR.t3700 VGND 0.00433f
C38256 VPWR.t2971 VGND 0.00433f
C38257 VPWR.t7091 VGND 0.00433f
C38258 VPWR.t3867 VGND 0.00433f
C38259 VPWR.t4241 VGND 0.00433f
C38260 VPWR.t3504 VGND 0.00433f
C38261 VPWR.t785 VGND 0.00433f
C38262 VPWR.t3682 VGND 0.00433f
C38263 VPWR.t4946 VGND 0.05247f
C38264 VPWR.t6222 VGND 0.05996f
C38265 VPWR.t2688 VGND 0.05996f
C38266 VPWR.t3758 VGND 0.05996f
C38267 VPWR.t5734 VGND 0.05996f
C38268 VPWR.t2567 VGND 0.05996f
C38269 VPWR.t3438 VGND 0.05996f
C38270 VPWR.t3375 VGND 0.04035f
C38271 VPWR.t3699 VGND 0.04035f
C38272 VPWR.t2970 VGND 0.05996f
C38273 VPWR.t7090 VGND 0.05996f
C38274 VPWR.t3866 VGND 0.05996f
C38275 VPWR.t4240 VGND 0.05996f
C38276 VPWR.t3503 VGND 0.05996f
C38277 VPWR.t784 VGND 0.05996f
C38278 VPWR.t3681 VGND 0.05247f
C38279 VPWR.n39 VGND 0.03832f
C38280 VPWR.t3376 VGND 0.00433f
C38281 VPWR.t3439 VGND 0.00433f
C38282 VPWR.t2568 VGND 0.00433f
C38283 VPWR.t5735 VGND 0.00433f
C38284 VPWR.t3759 VGND 0.00433f
C38285 VPWR.t2689 VGND 0.00433f
C38286 VPWR.t6223 VGND 0.00433f
C38287 VPWR.n40 VGND 0.0178f
C38288 VPWR.n41 VGND 0.0178f
C38289 VPWR.n42 VGND 0.01679f
C38290 VPWR.n43 VGND 0.01186f
C38291 VPWR.n44 VGND 0.0178f
C38292 VPWR.n45 VGND 0.0178f
C38293 VPWR.n46 VGND 0.01839f
C38294 VPWR.n47 VGND 0.01189f
C38295 VPWR.n48 VGND 0.01371f
C38296 VPWR.n49 VGND 0.0178f
C38297 VPWR.n50 VGND 0.0178f
C38298 VPWR.n51 VGND 0.01679f
C38299 VPWR.n52 VGND 0.01186f
C38300 VPWR.n53 VGND 0.0178f
C38301 VPWR.n54 VGND 0.0178f
C38302 VPWR.n55 VGND 0.01839f
C38303 VPWR.n56 VGND 0.01189f
C38304 VPWR.n57 VGND 0.03832f
C38305 VPWR.t6118 VGND 0.05247f
C38306 VPWR.t3605 VGND 0.05996f
C38307 VPWR.t5266 VGND 0.05996f
C38308 VPWR.t5388 VGND 0.05996f
C38309 VPWR.t3778 VGND 0.05996f
C38310 VPWR.t1198 VGND 0.05996f
C38311 VPWR.t74 VGND 0.05996f
C38312 VPWR.t5650 VGND 0.04035f
C38313 VPWR.n58 VGND 0.03832f
C38314 VPWR.t5518 VGND 0.00433f
C38315 VPWR.t3135 VGND 0.00433f
C38316 VPWR.t7093 VGND 0.00433f
C38317 VPWR.t2977 VGND 0.00433f
C38318 VPWR.t561 VGND 0.00433f
C38319 VPWR.t6438 VGND 0.00433f
C38320 VPWR.t917 VGND 0.00433f
C38321 VPWR.t2424 VGND 0.00433f
C38322 VPWR.t5517 VGND 0.05247f
C38323 VPWR.t3134 VGND 0.05996f
C38324 VPWR.t7092 VGND 0.05996f
C38325 VPWR.t2976 VGND 0.05996f
C38326 VPWR.t560 VGND 0.05996f
C38327 VPWR.t6437 VGND 0.05996f
C38328 VPWR.t916 VGND 0.05996f
C38329 VPWR.t2423 VGND 0.04035f
C38330 VPWR.n59 VGND 0.03832f
C38331 VPWR.t955 VGND 0.00433f
C38332 VPWR.t1822 VGND 0.00433f
C38333 VPWR.n60 VGND 0.01293f
C38334 VPWR.n61 VGND 1.23893f
C38335 VPWR.t5226 VGND 0.00433f
C38336 VPWR.n62 VGND 0.00878f
C38337 VPWR.t6124 VGND 0.00433f
C38338 VPWR.t1542 VGND 0.00433f
C38339 VPWR.t4141 VGND 0.00433f
C38340 VPWR.t4292 VGND 0.00433f
C38341 VPWR.t4779 VGND 0.00433f
C38342 VPWR.t3518 VGND 0.00433f
C38343 VPWR.t4735 VGND 0.00433f
C38344 VPWR.t4923 VGND 0.00433f
C38345 VPWR.t455 VGND 0.00433f
C38346 VPWR.t4350 VGND 0.00433f
C38347 VPWR.t2683 VGND 0.00433f
C38348 VPWR.t1820 VGND 0.00433f
C38349 VPWR.t5536 VGND 0.00433f
C38350 VPWR.t4745 VGND 0.00433f
C38351 VPWR.t550 VGND 0.00433f
C38352 VPWR.t6226 VGND 0.00433f
C38353 VPWR.t1552 VGND 0.00433f
C38354 VPWR.t2882 VGND 0.00433f
C38355 VPWR.t513 VGND 0.00433f
C38356 VPWR.t5687 VGND 0.00433f
C38357 VPWR.t390 VGND 0.00433f
C38358 VPWR.t2989 VGND 0.00433f
C38359 VPWR.t1285 VGND 0.00433f
C38360 VPWR.t4582 VGND 0.00433f
C38361 VPWR.t1980 VGND 0.00433f
C38362 VPWR.t1485 VGND 0.00433f
C38363 VPWR.t2607 VGND 0.00433f
C38364 VPWR.t3842 VGND 0.00433f
C38365 VPWR.t1630 VGND 0.00433f
C38366 VPWR.t4939 VGND 0.00433f
C38367 VPWR.t549 VGND 0.06731f
C38368 VPWR.t1551 VGND 0.10001f
C38369 VPWR.t512 VGND 0.10001f
C38370 VPWR.t389 VGND 0.10001f
C38371 VPWR.t1284 VGND 0.10001f
C38372 VPWR.t1484 VGND 0.10001f
C38373 VPWR.t2606 VGND 0.10001f
C38374 VPWR.t1629 VGND 0.08271f
C38375 VPWR.n63 VGND 0.02102f
C38376 VPWR.t1100 VGND 0.00433f
C38377 VPWR.t2042 VGND 0.08751f
C38378 VPWR.t4612 VGND 0.10001f
C38379 VPWR.t1190 VGND 0.10001f
C38380 VPWR.t1186 VGND 0.10001f
C38381 VPWR.t2624 VGND 0.10001f
C38382 VPWR.t952 VGND 0.10001f
C38383 VPWR.t1145 VGND 0.06731f
C38384 VPWR.t1099 VGND 0.0202f
C38385 VPWR.t5726 VGND 0.0298f
C38386 VPWR.n64 VGND 0.03642f
C38387 VPWR.t5727 VGND 0.00433f
C38388 VPWR.t1146 VGND 0.00433f
C38389 VPWR.t3619 VGND 0.00433f
C38390 VPWR.t5576 VGND 0.00433f
C38391 VPWR.t953 VGND 0.00433f
C38392 VPWR.t2625 VGND 0.00433f
C38393 VPWR.t2978 VGND 0.00433f
C38394 VPWR.t1187 VGND 0.00433f
C38395 VPWR.t7079 VGND 0.00433f
C38396 VPWR.t1191 VGND 0.00433f
C38397 VPWR.t5664 VGND 0.00433f
C38398 VPWR.n65 VGND 0.02171f
C38399 VPWR.n66 VGND 0.0207f
C38400 VPWR.n67 VGND 0.01577f
C38401 VPWR.n68 VGND 0.02171f
C38402 VPWR.n69 VGND 0.02171f
C38403 VPWR.n70 VGND 0.01144f
C38404 VPWR.n71 VGND 0.01189f
C38405 VPWR.n72 VGND 0.00912f
C38406 VPWR.n73 VGND 0.01189f
C38407 VPWR.n74 VGND 0.01762f
C38408 VPWR.n75 VGND 0.02171f
C38409 VPWR.n76 VGND 0.02171f
C38410 VPWR.n77 VGND 0.0207f
C38411 VPWR.n78 VGND 0.01577f
C38412 VPWR.n79 VGND 0.02171f
C38413 VPWR.n80 VGND 0.02171f
C38414 VPWR.n81 VGND 0.02079f
C38415 VPWR.n82 VGND 0.00541f
C38416 VPWR.t4556 VGND 0.00433f
C38417 VPWR.n83 VGND 0.01023f
C38418 VPWR.n84 VGND 0.01189f
C38419 VPWR.n85 VGND 0.03642f
C38420 VPWR.t4744 VGND 0.03751f
C38421 VPWR.t4555 VGND 0.05001f
C38422 VPWR.t5225 VGND 0.05001f
C38423 VPWR.t6123 VGND 0.05001f
C38424 VPWR.t1541 VGND 0.05001f
C38425 VPWR.t4140 VGND 0.05001f
C38426 VPWR.t4291 VGND 0.05001f
C38427 VPWR.t4778 VGND 0.05001f
C38428 VPWR.t3517 VGND 0.05001f
C38429 VPWR.t4734 VGND 0.05001f
C38430 VPWR.t4922 VGND 0.05001f
C38431 VPWR.t454 VGND 0.05001f
C38432 VPWR.t4349 VGND 0.05001f
C38433 VPWR.t2682 VGND 0.05001f
C38434 VPWR.t1819 VGND 0.04231f
C38435 VPWR.t5535 VGND 0.0202f
C38436 VPWR.n86 VGND 0.02102f
C38437 VPWR.t663 VGND 0.00433f
C38438 VPWR.n87 VGND 0.03642f
C38439 VPWR.t6206 VGND 0.00433f
C38440 VPWR.t4503 VGND 0.00433f
C38441 VPWR.t5843 VGND 0.00433f
C38442 VPWR.t814 VGND 0.00433f
C38443 VPWR.t3526 VGND 0.00433f
C38444 VPWR.t432 VGND 0.00433f
C38445 VPWR.t345 VGND 0.00433f
C38446 VPWR.t4402 VGND 0.00433f
C38447 VPWR.t6197 VGND 0.00433f
C38448 VPWR.t2790 VGND 0.00433f
C38449 VPWR.t2211 VGND 0.00433f
C38450 VPWR.t3695 VGND 0.00433f
C38451 VPWR.t2372 VGND 0.00433f
C38452 VPWR.t5080 VGND 0.00433f
C38453 VPWR.t2311 VGND 0.00433f
C38454 VPWR.t6011 VGND 0.00433f
C38455 VPWR.t662 VGND 0.0298f
C38456 VPWR.t6205 VGND 0.03271f
C38457 VPWR.t4502 VGND 0.05001f
C38458 VPWR.t5842 VGND 0.05001f
C38459 VPWR.t813 VGND 0.05001f
C38460 VPWR.t3525 VGND 0.05001f
C38461 VPWR.t431 VGND 0.05001f
C38462 VPWR.t344 VGND 0.05001f
C38463 VPWR.t4401 VGND 0.05001f
C38464 VPWR.t6196 VGND 0.05001f
C38465 VPWR.t2789 VGND 0.05001f
C38466 VPWR.t2210 VGND 0.05001f
C38467 VPWR.t3694 VGND 0.05001f
C38468 VPWR.t2371 VGND 0.05001f
C38469 VPWR.t5079 VGND 0.05001f
C38470 VPWR.t2310 VGND 0.04231f
C38471 VPWR.t6010 VGND 0.0202f
C38472 VPWR.n88 VGND 0.05372f
C38473 VPWR.t5802 VGND 0.00433f
C38474 VPWR.t4250 VGND 0.00433f
C38475 VPWR.t650 VGND 0.00433f
C38476 VPWR.t1374 VGND 0.00433f
C38477 VPWR.t4885 VGND 0.00433f
C38478 VPWR.t2280 VGND 0.00433f
C38479 VPWR.t3707 VGND 0.00433f
C38480 VPWR.t77 VGND 0.00433f
C38481 VPWR.t357 VGND 0.00433f
C38482 VPWR.t637 VGND 0.00433f
C38483 VPWR.t1301 VGND 0.00433f
C38484 VPWR.t4730 VGND 0.00433f
C38485 VPWR.t1365 VGND 0.00433f
C38486 VPWR.t1470 VGND 0.00433f
C38487 VPWR.t3126 VGND 0.00433f
C38488 VPWR.t1508 VGND 0.00433f
C38489 VPWR.t4249 VGND 0.08751f
C38490 VPWR.t649 VGND 0.10001f
C38491 VPWR.t2279 VGND 0.10001f
C38492 VPWR.t76 VGND 0.10001f
C38493 VPWR.t356 VGND 0.10001f
C38494 VPWR.t1300 VGND 0.10001f
C38495 VPWR.t1364 VGND 0.10001f
C38496 VPWR.t1507 VGND 0.06731f
C38497 VPWR.n89 VGND 0.02233f
C38498 VPWR.n90 VGND 0.02171f
C38499 VPWR.n91 VGND 0.02171f
C38500 VPWR.n92 VGND 0.01577f
C38501 VPWR.n93 VGND 0.0207f
C38502 VPWR.n94 VGND 0.02134f
C38503 VPWR.n95 VGND 0.0184f
C38504 VPWR.t4968 VGND 0.00433f
C38505 VPWR.t4286 VGND 0.00433f
C38506 VPWR.n96 VGND 0.01513f
C38507 VPWR.t5101 VGND 0.00433f
C38508 VPWR.t3743 VGND 0.00433f
C38509 VPWR.t6439 VGND 0.00433f
C38510 VPWR.t1608 VGND 0.00433f
C38511 VPWR.t5418 VGND 0.00433f
C38512 VPWR.t2664 VGND 0.00433f
C38513 VPWR.t4620 VGND 0.00433f
C38514 VPWR.t2000 VGND 0.00433f
C38515 VPWR.t2016 VGND 0.00433f
C38516 VPWR.t3957 VGND 0.00433f
C38517 VPWR.t87 VGND 0.00433f
C38518 VPWR.t5513 VGND 0.00433f
C38519 VPWR.t754 VGND 0.0202f
C38520 VPWR.t755 VGND 0.00433f
C38521 VPWR.t3209 VGND 0.00433f
C38522 VPWR.t4507 VGND 0.00433f
C38523 VPWR.t6171 VGND 0.00433f
C38524 VPWR.t7078 VGND 0.00433f
C38525 VPWR.t5263 VGND 0.00433f
C38526 VPWR.t2775 VGND 0.00433f
C38527 VPWR.t3702 VGND 0.00433f
C38528 VPWR.t1197 VGND 0.00433f
C38529 VPWR.t5432 VGND 0.00433f
C38530 VPWR.t5795 VGND 0.00433f
C38531 VPWR.t5240 VGND 0.00433f
C38532 VPWR.t2548 VGND 0.00433f
C38533 VPWR.t5180 VGND 0.00433f
C38534 VPWR.t376 VGND 0.00433f
C38535 VPWR.t4471 VGND 0.00433f
C38536 VPWR.t3208 VGND 0.04231f
C38537 VPWR.t4506 VGND 0.05001f
C38538 VPWR.t6170 VGND 0.05001f
C38539 VPWR.t7077 VGND 0.05001f
C38540 VPWR.t5262 VGND 0.05001f
C38541 VPWR.t2774 VGND 0.05001f
C38542 VPWR.t3701 VGND 0.05001f
C38543 VPWR.t1196 VGND 0.05001f
C38544 VPWR.t5431 VGND 0.05001f
C38545 VPWR.t5794 VGND 0.05001f
C38546 VPWR.t5239 VGND 0.05001f
C38547 VPWR.t2547 VGND 0.05001f
C38548 VPWR.t5179 VGND 0.05001f
C38549 VPWR.t375 VGND 0.05001f
C38550 VPWR.t4470 VGND 0.03271f
C38551 VPWR.t6442 VGND 0.0298f
C38552 VPWR.n97 VGND 0.03642f
C38553 VPWR.t6443 VGND 0.00433f
C38554 VPWR.n98 VGND 0.02102f
C38555 VPWR.t2800 VGND 0.00433f
C38556 VPWR.t1462 VGND 0.00433f
C38557 VPWR.t6072 VGND 0.00433f
C38558 VPWR.t443 VGND 0.00433f
C38559 VPWR.t3367 VGND 0.00433f
C38560 VPWR.t696 VGND 0.00433f
C38561 VPWR.t6285 VGND 0.00433f
C38562 VPWR.t5137 VGND 0.00433f
C38563 VPWR.t1154 VGND 0.00433f
C38564 VPWR.t1231 VGND 0.00433f
C38565 VPWR.t3999 VGND 0.00433f
C38566 VPWR.t3314 VGND 0.00433f
C38567 VPWR.t1458 VGND 0.00433f
C38568 VPWR.t1246 VGND 0.00433f
C38569 VPWR.t3920 VGND 0.00433f
C38570 VPWR.t2799 VGND 0.0202f
C38571 VPWR.t1461 VGND 0.04231f
C38572 VPWR.t6071 VGND 0.05001f
C38573 VPWR.t442 VGND 0.05001f
C38574 VPWR.t3366 VGND 0.05001f
C38575 VPWR.t695 VGND 0.05001f
C38576 VPWR.t6284 VGND 0.05001f
C38577 VPWR.t5136 VGND 0.05001f
C38578 VPWR.t1153 VGND 0.05001f
C38579 VPWR.t1230 VGND 0.05001f
C38580 VPWR.t3998 VGND 0.05001f
C38581 VPWR.t3313 VGND 0.05001f
C38582 VPWR.t1457 VGND 0.05001f
C38583 VPWR.t1245 VGND 0.05001f
C38584 VPWR.t3919 VGND 0.05001f
C38585 VPWR.t707 VGND 0.03751f
C38586 VPWR.n99 VGND 0.03642f
C38587 VPWR.t708 VGND 0.00433f
C38588 VPWR.t6451 VGND 0.00433f
C38589 VPWR.t1917 VGND 0.00433f
C38590 VPWR.t7071 VGND 0.00433f
C38591 VPWR.t1219 VGND 0.00433f
C38592 VPWR.t5573 VGND 0.00433f
C38593 VPWR.t6233 VGND 0.00433f
C38594 VPWR.t3786 VGND 0.00433f
C38595 VPWR.t4729 VGND 0.00433f
C38596 VPWR.t1548 VGND 0.00433f
C38597 VPWR.t5749 VGND 0.00433f
C38598 VPWR.t656 VGND 0.00433f
C38599 VPWR.t4426 VGND 0.00433f
C38600 VPWR.t7081 VGND 0.00433f
C38601 VPWR.t3502 VGND 0.00433f
C38602 VPWR.t79 VGND 0.00433f
C38603 VPWR.t3843 VGND 0.00433f
C38604 VPWR.t1916 VGND 0.06731f
C38605 VPWR.t1218 VGND 0.10001f
C38606 VPWR.t5572 VGND 0.10001f
C38607 VPWR.t3785 VGND 0.10001f
C38608 VPWR.t1547 VGND 0.10001f
C38609 VPWR.t655 VGND 0.10001f
C38610 VPWR.t3501 VGND 0.10001f
C38611 VPWR.t78 VGND 0.08271f
C38612 VPWR.n100 VGND 0.02102f
C38613 VPWR.t4259 VGND 0.00433f
C38614 VPWR.t4258 VGND 0.0202f
C38615 VPWR.t5416 VGND 0.0298f
C38616 VPWR.n101 VGND 0.03642f
C38617 VPWR.t5417 VGND 0.00433f
C38618 VPWR.t2404 VGND 0.00433f
C38619 VPWR.t2871 VGND 0.00433f
C38620 VPWR.t7133 VGND 0.00433f
C38621 VPWR.t3075 VGND 0.00433f
C38622 VPWR.t6362 VGND 0.00433f
C38623 VPWR.t2587 VGND 0.00431f
C38624 VPWR.t4118 VGND 0.00433f
C38625 VPWR.t139 VGND 0.00116f
C38626 VPWR.t6491 VGND 0.00116f
C38627 VPWR.n102 VGND 0.00236f
C38628 VPWR.t6895 VGND 0.00185f
C38629 VPWR.t4390 VGND 0.00219f
C38630 VPWR.n103 VGND 0.00433f
C38631 VPWR.t6098 VGND 0.00255f
C38632 VPWR.n104 VGND 0.01415f
C38633 VPWR.n105 VGND 0.13412f
C38634 VPWR.t3670 VGND 0.00127f
C38635 VPWR.n106 VGND 0.00342f
C38636 VPWR.n107 VGND 0.00619f
C38637 VPWR.t3222 VGND 0.00433f
C38638 VPWR.n108 VGND 0.00115f
C38639 VPWR.t3411 VGND 0.0202f
C38640 VPWR.t2751 VGND 0.00433f
C38641 VPWR.n109 VGND 0.00115f
C38642 VPWR.t6321 VGND 0.00433f
C38643 VPWR.t1255 VGND 0.00431f
C38644 VPWR.t2520 VGND 0.00107f
C38645 VPWR.n110 VGND 0.00292f
C38646 VPWR.t613 VGND 0.00427f
C38647 VPWR.t1257 VGND 0.00183f
C38648 VPWR.t2228 VGND 0.00157f
C38649 VPWR.n111 VGND 0.00508f
C38650 VPWR.t4090 VGND 0.00203f
C38651 VPWR.t4092 VGND 0.0031f
C38652 VPWR.t2563 VGND 0.00114f
C38653 VPWR.t2556 VGND 0.00114f
C38654 VPWR.n112 VGND 0.00231f
C38655 VPWR.t6403 VGND 0.00425f
C38656 VPWR.t4088 VGND 0.00114f
C38657 VPWR.t4083 VGND 0.00114f
C38658 VPWR.n113 VGND 0.00231f
C38659 VPWR.t4388 VGND 0.00433f
C38660 VPWR.t2750 VGND 0.02147f
C38661 VPWR.t6215 VGND 0.01772f
C38662 VPWR.n114 VGND 0.02438f
C38663 VPWR.t104 VGND 0.02478f
C38664 VPWR.t1676 VGND 0.03014f
C38665 VPWR.t6320 VGND 0.02411f
C38666 VPWR.t4251 VGND 0.03271f
C38667 VPWR.t105 VGND 0.03427f
C38668 VPWR.t4084 VGND 0.03181f
C38669 VPWR.t3413 VGND 0.02612f
C38670 VPWR.t614 VGND 0.02913f
C38671 VPWR.t2519 VGND 0.03561f
C38672 VPWR.t2227 VGND 0.03885f
C38673 VPWR.t612 VGND 0.02992f
C38674 VPWR.t1256 VGND 0.03349f
C38675 VPWR.t4089 VGND 0.02489f
C38676 VPWR.t3635 VGND 0.0154f
C38677 VPWR.t6854 VGND 0.01172f
C38678 VPWR.t4091 VGND 0.025f
C38679 VPWR.t2555 VGND 0.02545f
C38680 VPWR.t6402 VGND 0.02277f
C38681 VPWR.t2562 VGND 0.03784f
C38682 VPWR.t4082 VGND 0.0173f
C38683 VPWR.t4387 VGND 0.02277f
C38684 VPWR.t4087 VGND 0.03326f
C38685 VPWR.t2557 VGND 0.02701f
C38686 VPWR.n115 VGND 0.02649f
C38687 VPWR.t2561 VGND 0.00114f
C38688 VPWR.t2558 VGND 0.00114f
C38689 VPWR.n116 VGND 0.00231f
C38690 VPWR.t6849 VGND 0.00114f
C38691 VPWR.t4086 VGND 0.00114f
C38692 VPWR.n117 VGND 0.00231f
C38693 VPWR.t882 VGND 0.00433f
C38694 VPWR.t5753 VGND 0.00433f
C38695 VPWR.t6413 VGND 0.00114f
C38696 VPWR.t6411 VGND 0.00306f
C38697 VPWR.n118 VGND 0.00423f
C38698 VPWR.n119 VGND 0.00426f
C38699 VPWR.n120 VGND 0.20174f
C38700 VPWR.n121 VGND 0.13412f
C38701 VPWR.t5779 VGND 0.00433f
C38702 VPWR.t4995 VGND 0.00433f
C38703 VPWR.n122 VGND 0.01238f
C38704 VPWR.t2955 VGND 0.00431f
C38705 VPWR.t949 VGND 0.00427f
C38706 VPWR.t3659 VGND 0.00107f
C38707 VPWR.n123 VGND 0.00292f
C38708 VPWR.t6966 VGND 0.0202f
C38709 VPWR.t6967 VGND 0.00425f
C38710 VPWR.t4562 VGND 0.00334f
C38711 VPWR.n124 VGND 0.00145f
C38712 VPWR.t7110 VGND 0.00132f
C38713 VPWR.t6971 VGND 0.00132f
C38714 VPWR.n125 VGND 0.00267f
C38715 VPWR.t6987 VGND 0.00196f
C38716 VPWR.t1084 VGND 0.00157f
C38717 VPWR.n126 VGND 0.00539f
C38718 VPWR.t3647 VGND 0.00433f
C38719 VPWR.t113 VGND 0.00431f
C38720 VPWR.t3493 VGND 0.00433f
C38721 VPWR.t6259 VGND 0.00433f
C38722 VPWR.t6214 VGND 0.00433f
C38723 VPWR.t478 VGND 0.00516f
C38724 VPWR.t6528 VGND 0.00425f
C38725 VPWR.t3472 VGND 0.00375f
C38726 VPWR.t3993 VGND 0.00434f
C38727 VPWR.t2351 VGND 0.00132f
C38728 VPWR.t6530 VGND 0.00132f
C38729 VPWR.n127 VGND 0.00266f
C38730 VPWR.t4561 VGND 0.01172f
C38731 VPWR.t6968 VGND 0.02277f
C38732 VPWR.t6970 VGND 0.02277f
C38733 VPWR.t4558 VGND 0.02277f
C38734 VPWR.t7109 VGND 0.02277f
C38735 VPWR.t6986 VGND 0.02724f
C38736 VPWR.t1083 VGND 0.0173f
C38737 VPWR.t3646 VGND 0.03516f
C38738 VPWR.t3492 VGND 0.01172f
C38739 VPWR.t112 VGND 0.03304f
C38740 VPWR.t7111 VGND 0.04309f
C38741 VPWR.t6258 VGND 0.03717f
C38742 VPWR.t474 VGND 0.0125f
C38743 VPWR.t6213 VGND 0.02199f
C38744 VPWR.t3473 VGND 0.03795f
C38745 VPWR.t6527 VGND 0.02802f
C38746 VPWR.t477 VGND 0.03672f
C38747 VPWR.t3470 VGND 0.02355f
C38748 VPWR.t3471 VGND 0.02645f
C38749 VPWR.t3992 VGND 0.02277f
C38750 VPWR.t6529 VGND 0.03125f
C38751 VPWR.t2350 VGND 0.03237f
C38752 VPWR.n128 VGND 0.02649f
C38753 VPWR.t6541 VGND 0.00132f
C38754 VPWR.t2358 VGND 0.00132f
C38755 VPWR.n129 VGND 0.00266f
C38756 VPWR.t3483 VGND 0.0033f
C38757 VPWR.t6770 VGND 0.00425f
C38758 VPWR.t481 VGND 0.00196f
C38759 VPWR.t3183 VGND 0.00157f
C38760 VPWR.n130 VGND 0.00539f
C38761 VPWR.n131 VGND 0.00981f
C38762 VPWR.n132 VGND 0.13412f
C38763 VPWR.n133 VGND 0.13412f
C38764 VPWR.t3869 VGND 0.00427f
C38765 VPWR.n134 VGND 0.00461f
C38766 VPWR.t5915 VGND 0.00107f
C38767 VPWR.n135 VGND 0.00292f
C38768 VPWR.t4709 VGND 0.00433f
C38769 VPWR.n136 VGND 0.03006f
C38770 VPWR.t4748 VGND 0.00433f
C38771 VPWR.n137 VGND 0.00115f
C38772 VPWR.t4041 VGND 0.00433f
C38773 VPWR.t5912 VGND 0.00255f
C38774 VPWR.t2784 VGND 0.00427f
C38775 VPWR.t38 VGND 0.00116f
C38776 VPWR.t6489 VGND 0.00116f
C38777 VPWR.n138 VGND 0.00236f
C38778 VPWR.t3163 VGND 0.00107f
C38779 VPWR.n139 VGND 0.00292f
C38780 VPWR.t1636 VGND 0.00433f
C38781 VPWR.t476 VGND 0.00431f
C38782 VPWR.n140 VGND 0.00115f
C38783 VPWR.t355 VGND 0.00433f
C38784 VPWR.t6318 VGND 0.00255f
C38785 VPWR.t3129 VGND 0.01772f
C38786 VPWR.t6073 VGND 0.01775f
C38787 VPWR.t4040 VGND 0.02143f
C38788 VPWR.t40 VGND 0.0173f
C38789 VPWR.t6153 VGND 0.03271f
C38790 VPWR.t4747 VGND 0.02411f
C38791 VPWR.t435 VGND 0.03014f
C38792 VPWR.t39 VGND 0.02478f
C38793 VPWR.n141 VGND 0.02438f
C38794 VPWR.t5911 VGND 0.03561f
C38795 VPWR.t2783 VGND 0.04822f
C38796 VPWR.t37 VGND 0.03885f
C38797 VPWR.t3162 VGND 0.02277f
C38798 VPWR.t6488 VGND 0.02556f
C38799 VPWR.t2781 VGND 0.01953f
C38800 VPWR.t6319 VGND 0.03058f
C38801 VPWR.t1635 VGND 0.03047f
C38802 VPWR.t6387 VGND 0.0154f
C38803 VPWR.t475 VGND 0.01931f
C38804 VPWR.t3130 VGND 0.02277f
C38805 VPWR.t4837 VGND 0.02411f
C38806 VPWR.t2323 VGND 0.02322f
C38807 VPWR.t6386 VGND 0.01831f
C38808 VPWR.t6676 VGND 0.00826f
C38809 VPWR.n142 VGND 0.05913f
C38810 VPWR.t6317 VGND 0.0211f
C38811 VPWR.t354 VGND 0.02244f
C38812 VPWR.n143 VGND 0.0295f
C38813 VPWR.t6389 VGND 0.00116f
C38814 VPWR.t6471 VGND 0.00116f
C38815 VPWR.n144 VGND 0.00236f
C38816 VPWR.t4204 VGND 0.00427f
C38817 VPWR.t463 VGND 0.00107f
C38818 VPWR.n145 VGND 0.00292f
C38819 VPWR.t6679 VGND 0.00429f
C38820 VPWR.n146 VGND 0.00115f
C38821 VPWR.t372 VGND 0.00433f
C38822 VPWR.t6994 VGND 0.0019f
C38823 VPWR.t6293 VGND 0.00255f
C38824 VPWR.t170 VGND 0.00156f
C38825 VPWR.n147 VGND 0.00505f
C38826 VPWR.t6740 VGND 0.00116f
C38827 VPWR.t6475 VGND 0.00116f
C38828 VPWR.n148 VGND 0.00236f
C38829 VPWR.t6989 VGND 0.00374f
C38830 VPWR.t5856 VGND 0.00427f
C38831 VPWR.t2574 VGND 0.01733f
C38832 VPWR.t6388 VGND 0.02835f
C38833 VPWR.t6470 VGND 0.03483f
C38834 VPWR.t4203 VGND 0.01395f
C38835 VPWR.t462 VGND 0.025f
C38836 VPWR.t4201 VGND 0.01183f
C38837 VPWR.t6990 VGND 0.01741f
C38838 VPWR.t6291 VGND 0.02277f
C38839 VPWR.t4560 VGND 0.03047f
C38840 VPWR.t2990 VGND 0.02634f
C38841 VPWR.t6741 VGND 0.025f
C38842 VPWR.t6678 VGND 0.03338f
C38843 VPWR.t2966 VGND 0.03382f
C38844 VPWR.t932 VGND 0.04063f
C38845 VPWR.t6776 VGND 0.02389f
C38846 VPWR.t371 VGND 0.02969f
C38847 VPWR.n150 VGND 0.01275f
C38848 VPWR.t6292 VGND 0.01485f
C38849 VPWR.t6993 VGND 0.02545f
C38850 VPWR.t169 VGND 0.04554f
C38851 VPWR.t6739 VGND 0.02902f
C38852 VPWR.t5707 VGND 0.02277f
C38853 VPWR.t6474 VGND 0.02389f
C38854 VPWR.t171 VGND 0.01172f
C38855 VPWR.t6988 VGND 0.03656f
C38856 VPWR.t5855 VGND 0.04309f
C38857 VPWR.n151 VGND 0.04256f
C38858 VPWR.t4072 VGND 0.00107f
C38859 VPWR.n152 VGND 0.00292f
C38860 VPWR.t1994 VGND 0.00433f
C38861 VPWR.t1384 VGND 0.00433f
C38862 VPWR.t4331 VGND 0.00433f
C38863 VPWR.n153 VGND 0.00115f
C38864 VPWR.t2802 VGND 0.00433f
C38865 VPWR.t6364 VGND 0.00433f
C38866 VPWR.t4423 VGND 0.00255f
C38867 VPWR.t7028 VGND 0.00116f
C38868 VPWR.t6465 VGND 0.00116f
C38869 VPWR.n154 VGND 0.00236f
C38870 VPWR.t1996 VGND 0.00433f
C38871 VPWR.t4715 VGND 0.00433f
C38872 VPWR.t4053 VGND 0.00433f
C38873 VPWR.t2416 VGND 0.00433f
C38874 VPWR.t2246 VGND 0.00433f
C38875 VPWR.t3203 VGND 0.00433f
C38876 VPWR.t2956 VGND 0.02356f
C38877 VPWR.t2801 VGND 0.01563f
C38878 VPWR.t4071 VGND 0.03192f
C38879 VPWR.t5857 VGND 0.03326f
C38880 VPWR.t1993 VGND 0.01741f
C38881 VPWR.t4421 VGND 0.0173f
C38882 VPWR.t7030 VGND 0.03271f
C38883 VPWR.t1383 VGND 0.03338f
C38884 VPWR.t4742 VGND 0.05001f
C38885 VPWR.t4330 VGND 0.02411f
C38886 VPWR.t5089 VGND 0.01764f
C38887 VPWR.t7029 VGND 0.02478f
C38888 VPWR.n156 VGND 0.03945f
C38889 VPWR.t4422 VGND 0.0461f
C38890 VPWR.t6363 VGND 0.04822f
C38891 VPWR.t7027 VGND 0.04085f
C38892 VPWR.t6464 VGND 0.03192f
C38893 VPWR.t1995 VGND 0.01395f
C38894 VPWR.t4714 VGND 0.03271f
C38895 VPWR.t4052 VGND 0.05001f
C38896 VPWR.t2415 VGND 0.05001f
C38897 VPWR.t2245 VGND 0.0298f
C38898 VPWR.t3202 VGND 0.06143f
C38899 VPWR.t5499 VGND 0.00433f
C38900 VPWR.t2615 VGND 0.00433f
C38901 VPWR.t5434 VGND 0.00433f
C38902 VPWR.t3946 VGND 0.00433f
C38903 VPWR.t1414 VGND 0.00433f
C38904 VPWR.t1594 VGND 0.00433f
C38905 VPWR.t5776 VGND 0.00433f
C38906 VPWR.t6459 VGND 0.00433f
C38907 VPWR.t601 VGND 0.00433f
C38908 VPWR.t2432 VGND 0.00433f
C38909 VPWR.t5282 VGND 0.00433f
C38910 VPWR.t5532 VGND 0.00433f
C38911 VPWR.t4128 VGND 0.00433f
C38912 VPWR.t4593 VGND 0.00433f
C38913 VPWR.t6211 VGND 0.00433f
C38914 VPWR.t665 VGND 0.00433f
C38915 VPWR.t2794 VGND 0.00433f
C38916 VPWR.t5498 VGND 0.05001f
C38917 VPWR.t2614 VGND 0.0173f
C38918 VPWR.t5433 VGND 0.04521f
C38919 VPWR.t3945 VGND 0.05001f
C38920 VPWR.t1413 VGND 0.05001f
C38921 VPWR.t1593 VGND 0.05001f
C38922 VPWR.t5775 VGND 0.05001f
C38923 VPWR.t6458 VGND 0.05001f
C38924 VPWR.t600 VGND 0.05001f
C38925 VPWR.t2431 VGND 0.05001f
C38926 VPWR.t5281 VGND 0.05001f
C38927 VPWR.t5531 VGND 0.05001f
C38928 VPWR.t4127 VGND 0.05001f
C38929 VPWR.t4592 VGND 0.05001f
C38930 VPWR.t6210 VGND 0.05001f
C38931 VPWR.t664 VGND 0.0298f
C38932 VPWR.t2793 VGND 0.04122f
C38933 VPWR.t2128 VGND 0.00433f
C38934 VPWR.t5988 VGND 0.00433f
C38935 VPWR.t1477 VGND 0.00433f
C38936 VPWR.t6440 VGND 0.00433f
C38937 VPWR.t5902 VGND 0.00433f
C38938 VPWR.t6354 VGND 0.00433f
C38939 VPWR.t2687 VGND 0.00433f
C38940 VPWR.t1238 VGND 0.00433f
C38941 VPWR.t3616 VGND 0.00433f
C38942 VPWR.t3370 VGND 0.00433f
C38943 VPWR.t4974 VGND 0.00433f
C38944 VPWR.t2992 VGND 0.00433f
C38945 VPWR.t667 VGND 0.00433f
C38946 VPWR.t5124 VGND 0.00433f
C38947 VPWR.t3601 VGND 0.00433f
C38948 VPWR.t7089 VGND 0.00433f
C38949 VPWR.t2127 VGND 0.08271f
C38950 VPWR.t1476 VGND 0.10001f
C38951 VPWR.t5901 VGND 0.10001f
C38952 VPWR.t1237 VGND 0.10001f
C38953 VPWR.t3369 VGND 0.10001f
C38954 VPWR.t2991 VGND 0.10001f
C38955 VPWR.t666 VGND 0.10001f
C38956 VPWR.t3600 VGND 0.06731f
C38957 VPWR.n157 VGND 0.02233f
C38958 VPWR.n158 VGND 0.02171f
C38959 VPWR.n159 VGND 0.02171f
C38960 VPWR.n160 VGND 0.01577f
C38961 VPWR.n161 VGND 0.0207f
C38962 VPWR.n162 VGND 0.02171f
C38963 VPWR.n163 VGND 0.02171f
C38964 VPWR.n164 VGND 0.01568f
C38965 VPWR.n165 VGND 0.01165f
C38966 VPWR.n166 VGND 0.01144f
C38967 VPWR.n167 VGND 0.01085f
C38968 VPWR.n168 VGND 0.01085f
C38969 VPWR.n169 VGND 0.01017f
C38970 VPWR.n170 VGND 0.13412f
C38971 VPWR.t4944 VGND 0.00433f
C38972 VPWR.n171 VGND 0.0098f
C38973 VPWR.t1606 VGND 0.00433f
C38974 VPWR.t2098 VGND 0.00433f
C38975 VPWR.t5265 VGND 0.00433f
C38976 VPWR.t5834 VGND 0.00433f
C38977 VPWR.t5100 VGND 0.00433f
C38978 VPWR.t5332 VGND 0.00433f
C38979 VPWR.t4059 VGND 0.00433f
C38980 VPWR.t5781 VGND 0.00433f
C38981 VPWR.t3500 VGND 0.00433f
C38982 VPWR.t331 VGND 0.00433f
C38983 VPWR.t2386 VGND 0.00433f
C38984 VPWR.t4486 VGND 0.00433f
C38985 VPWR.t1852 VGND 0.00433f
C38986 VPWR.t5637 VGND 0.00433f
C38987 VPWR.t4392 VGND 0.00433f
C38988 VPWR.t3645 VGND 0.00433f
C38989 VPWR.t6350 VGND 0.00433f
C38990 VPWR.t5300 VGND 0.00433f
C38991 VPWR.t6242 VGND 0.00433f
C38992 VPWR.t449 VGND 0.00433f
C38993 VPWR.t5575 VGND 0.00433f
C38994 VPWR.t5331 VGND 0.0298f
C38995 VPWR.t4058 VGND 0.05001f
C38996 VPWR.t5780 VGND 0.05001f
C38997 VPWR.t3499 VGND 0.05001f
C38998 VPWR.t330 VGND 0.05001f
C38999 VPWR.t2385 VGND 0.05001f
C39000 VPWR.t4485 VGND 0.05001f
C39001 VPWR.t1851 VGND 0.05001f
C39002 VPWR.t5636 VGND 0.05001f
C39003 VPWR.t4391 VGND 0.05001f
C39004 VPWR.t3644 VGND 0.05001f
C39005 VPWR.t6349 VGND 0.05001f
C39006 VPWR.t5299 VGND 0.05001f
C39007 VPWR.t6241 VGND 0.04521f
C39008 VPWR.t448 VGND 0.0173f
C39009 VPWR.t5574 VGND 0.03271f
C39010 VPWR.t3271 VGND 0.04122f
C39011 VPWR.t3272 VGND 0.00433f
C39012 VPWR.t5381 VGND 0.00433f
C39013 VPWR.t2679 VGND 0.00433f
C39014 VPWR.t1386 VGND 0.00433f
C39015 VPWR.t4098 VGND 0.00433f
C39016 VPWR.n172 VGND 0.01082f
C39017 VPWR.t5645 VGND 0.00433f
C39018 VPWR.n173 VGND 0.01082f
C39019 VPWR.t4951 VGND 0.00433f
C39020 VPWR.t5954 VGND 0.00433f
C39021 VPWR.t3123 VGND 0.00433f
C39022 VPWR.t2026 VGND 0.00433f
C39023 VPWR.t2137 VGND 0.00433f
C39024 VPWR.t1179 VGND 0.00433f
C39025 VPWR.t3847 VGND 0.00433f
C39026 VPWR.t2909 VGND 0.00433f
C39027 VPWR.t1002 VGND 0.00433f
C39028 VPWR.t2080 VGND 0.00433f
C39029 VPWR.t4074 VGND 0.00433f
C39030 VPWR.t4895 VGND 0.00433f
C39031 VPWR.t6302 VGND 0.00433f
C39032 VPWR.t3781 VGND 0.00433f
C39033 VPWR.t3728 VGND 0.00433f
C39034 VPWR.t99 VGND 0.00116f
C39035 VPWR.t6666 VGND 0.00116f
C39036 VPWR.n174 VGND 0.00236f
C39037 VPWR.t5764 VGND 0.00433f
C39038 VPWR.t1468 VGND 0.00255f
C39039 VPWR.t5222 VGND 0.00433f
C39040 VPWR.t4542 VGND 0.00433f
C39041 VPWR.t1178 VGND 0.0298f
C39042 VPWR.t3846 VGND 0.05001f
C39043 VPWR.t2908 VGND 0.05001f
C39044 VPWR.t1001 VGND 0.05001f
C39045 VPWR.t2079 VGND 0.05001f
C39046 VPWR.t4073 VGND 0.05001f
C39047 VPWR.t4894 VGND 0.05001f
C39048 VPWR.t6301 VGND 0.03271f
C39049 VPWR.t3780 VGND 0.0298f
C39050 VPWR.t3727 VGND 0.03271f
C39051 VPWR.t6665 VGND 0.0173f
C39052 VPWR.t5763 VGND 0.02277f
C39053 VPWR.t98 VGND 0.05001f
C39054 VPWR.t5221 VGND 0.04822f
C39055 VPWR.t1467 VGND 0.03271f
C39056 VPWR.t5470 VGND 0.01775f
C39057 VPWR.t4541 VGND 0.02143f
C39058 VPWR.n175 VGND 0.02438f
C39059 VPWR.t101 VGND 0.02478f
C39060 VPWR.t2058 VGND 0.01764f
C39061 VPWR.n176 VGND 0.02504f
C39062 VPWR.n177 VGND 0.00115f
C39063 VPWR.t4718 VGND 0.00433f
C39064 VPWR.n178 VGND 0.13412f
C39065 VPWR.t83 VGND 0.00433f
C39066 VPWR.t2708 VGND 0.01775f
C39067 VPWR.t82 VGND 0.02143f
C39068 VPWR.t2001 VGND 0.0202f
C39069 VPWR.t2705 VGND 0.0018f
C39070 VPWR.t2002 VGND 0.00181f
C39071 VPWR.n179 VGND 0.00494f
C39072 VPWR.t2576 VGND 0.00431f
C39073 VPWR.t6882 VGND 0.00203f
C39074 VPWR.t2707 VGND 0.00431f
C39075 VPWR.t6169 VGND 0.00433f
C39076 VPWR.t3199 VGND 0.00433f
C39077 VPWR.t886 VGND 0.00433f
C39078 VPWR.t959 VGND 0.00394f
C39079 VPWR.t6581 VGND 0.00394f
C39080 VPWR.t6347 VGND 0.00433f
C39081 VPWR.t5877 VGND 0.00433f
C39082 VPWR.t6434 VGND 0.00433f
C39083 VPWR.t487 VGND 0.00433f
C39084 VPWR.t5328 VGND 0.00433f
C39085 VPWR.t1832 VGND 0.00433f
C39086 VPWR.t2818 VGND 0.00433f
C39087 VPWR.t2575 VGND 0.01261f
C39088 VPWR.t2704 VGND 0.02366f
C39089 VPWR.t6881 VGND 0.02523f
C39090 VPWR.t6582 VGND 0.01172f
C39091 VPWR.t2706 VGND 0.0125f
C39092 VPWR.t6168 VGND 0.02534f
C39093 VPWR.t6885 VGND 0.04521f
C39094 VPWR.t3198 VGND 0.0173f
C39095 VPWR.t885 VGND 0.03271f
C39096 VPWR.t958 VGND 0.0298f
C39097 VPWR.t6346 VGND 0.02277f
C39098 VPWR.t6580 VGND 0.03271f
C39099 VPWR.t5876 VGND 0.06731f
C39100 VPWR.t486 VGND 0.08271f
C39101 VPWR.t1831 VGND 0.05001f
C39102 VPWR.n180 VGND 0.02872f
C39103 VPWR.t5568 VGND 0.00431f
C39104 VPWR.t6822 VGND 0.00433f
C39105 VPWR.t2950 VGND 0.00375f
C39106 VPWR.t5567 VGND 0.025f
C39107 VPWR.t5665 VGND 0.03538f
C39108 VPWR.t6821 VGND 0.025f
C39109 VPWR.t214 VGND 0.01172f
C39110 VPWR.n181 VGND 0.04468f
C39111 VPWR.t6820 VGND 0.00394f
C39112 VPWR.n182 VGND 0.13412f
C39113 VPWR.n183 VGND 0.13412f
C39114 VPWR.t5976 VGND 0.00255f
C39115 VPWR.n184 VGND 0.00849f
C39116 VPWR.t585 VGND 0.00427f
C39117 VPWR.t7045 VGND 0.00116f
C39118 VPWR.t6662 VGND 0.00116f
C39119 VPWR.n185 VGND 0.00236f
C39120 VPWR.t589 VGND 0.00603f
C39121 VPWR.t1310 VGND 0.0202f
C39122 VPWR.t1311 VGND 0.00433f
C39123 VPWR.t978 VGND 0.00433f
C39124 VPWR.t5184 VGND 0.00433f
C39125 VPWR.t4467 VGND 0.00431f
C39126 VPWR.t4957 VGND 0.00433f
C39127 VPWR.t4740 VGND 0.00433f
C39128 VPWR.t2854 VGND 0.00433f
C39129 VPWR.t5559 VGND 0.00433f
C39130 VPWR.t6454 VGND 0.00433f
C39131 VPWR.t2893 VGND 0.00603f
C39132 VPWR.t364 VGND 0.00433f
C39133 VPWR.t2895 VGND 0.00427f
C39134 VPWR.t5426 VGND 0.00107f
C39135 VPWR.n186 VGND 0.00292f
C39136 VPWR.t3543 VGND 0.00433f
C39137 VPWR.t977 VGND 0.03538f
C39138 VPWR.t204 VGND 0.04309f
C39139 VPWR.t6290 VGND 0.03192f
C39140 VPWR.t5183 VGND 0.02277f
C39141 VPWR.t4466 VGND 0.0298f
C39142 VPWR.t4956 VGND 0.0173f
C39143 VPWR.t4739 VGND 0.05001f
C39144 VPWR.t2853 VGND 0.05001f
C39145 VPWR.t5558 VGND 0.04521f
C39146 VPWR.t6453 VGND 0.04744f
C39147 VPWR.t2892 VGND 0.05001f
C39148 VPWR.t363 VGND 0.02277f
C39149 VPWR.t2894 VGND 0.03271f
C39150 VPWR.t3542 VGND 0.02154f
C39151 VPWR.t5425 VGND 0.03192f
C39152 VPWR.t2890 VGND 0.02846f
C39153 VPWR.t5422 VGND 0.025f
C39154 VPWR.n187 VGND 0.02716f
C39155 VPWR.n188 VGND 0.00115f
C39156 VPWR.n189 VGND 0.00446f
C39157 VPWR.n190 VGND 0.13412f
C39158 VPWR.n191 VGND 0.13412f
C39159 VPWR.t4574 VGND 0.00433f
C39160 VPWR.n192 VGND 0.00695f
C39161 VPWR.t4337 VGND 0.00433f
C39162 VPWR.t7132 VGND 0.00433f
C39163 VPWR.t5950 VGND 0.00473f
C39164 VPWR.t5247 VGND 0.00433f
C39165 VPWR.t5952 VGND 0.00427f
C39166 VPWR.t5312 VGND 0.00433f
C39167 VPWR.t1121 VGND 0.00473f
C39168 VPWR.t5990 VGND 0.00473f
C39169 VPWR.t1119 VGND 0.00427f
C39170 VPWR.t5992 VGND 0.00427f
C39171 VPWR.t609 VGND 0.00427f
C39172 VPWR.t1127 VGND 0.00473f
C39173 VPWR.t607 VGND 0.00473f
C39174 VPWR.t1125 VGND 0.00427f
C39175 VPWR.t5322 VGND 0.00427f
C39176 VPWR.t2141 VGND 0.00433f
C39177 VPWR.t5320 VGND 0.00473f
C39178 VPWR.t3796 VGND 0.00433f
C39179 VPWR.t3763 VGND 0.00433f
C39180 VPWR.t3390 VGND 0.00433f
C39181 VPWR.t5246 VGND 0.03248f
C39182 VPWR.t5949 VGND 0.03271f
C39183 VPWR.t5311 VGND 0.02288f
C39184 VPWR.t5951 VGND 0.0173f
C39185 VPWR.t1120 VGND 0.03248f
C39186 VPWR.t5989 VGND 0.02791f
C39187 VPWR.t1118 VGND 0.02712f
C39188 VPWR.t5991 VGND 0.0125f
C39189 VPWR.t608 VGND 0.03248f
C39190 VPWR.t1126 VGND 0.02791f
C39191 VPWR.t606 VGND 0.02791f
C39192 VPWR.t1124 VGND 0.03248f
C39193 VPWR.t2140 VGND 0.01172f
C39194 VPWR.t5321 VGND 0.03483f
C39195 VPWR.t5319 VGND 0.04309f
C39196 VPWR.t3795 VGND 0.03538f
C39197 VPWR.t3762 VGND 0.0298f
C39198 VPWR.t3389 VGND 0.03271f
C39199 VPWR.n193 VGND 0.03352f
C39200 VPWR.t6312 VGND 0.00433f
C39201 VPWR.t4769 VGND 0.00433f
C39202 VPWR.n194 VGND 0.00735f
C39203 VPWR.n195 VGND 0.13412f
C39204 VPWR.n196 VGND 0.13412f
C39205 VPWR.t3574 VGND 0.00473f
C39206 VPWR.n197 VGND 0.00652f
C39207 VPWR.t4061 VGND 0.00473f
C39208 VPWR.t3572 VGND 0.00427f
C39209 VPWR.t2364 VGND 0.00427f
C39210 VPWR.t1514 VGND 0.00427f
C39211 VPWR.t2366 VGND 0.00473f
C39212 VPWR.t1512 VGND 0.00473f
C39213 VPWR.n198 VGND 0.0391f
C39214 VPWR.t1518 VGND 0.00427f
C39215 VPWR.t4666 VGND 0.00433f
C39216 VPWR.t1516 VGND 0.00473f
C39217 VPWR.t5484 VGND 0.00433f
C39218 VPWR.t2917 VGND 0.00427f
C39219 VPWR.t6156 VGND 0.00433f
C39220 VPWR.t2915 VGND 0.00473f
C39221 VPWR.t2264 VGND 0.00433f
C39222 VPWR.t5407 VGND 0.00433f
C39223 VPWR.t5224 VGND 0.00433f
C39224 VPWR.t2763 VGND 0.00433f
C39225 VPWR.t992 VGND 0.00433f
C39226 VPWR.t4705 VGND 0.00433f
C39227 VPWR.t1452 VGND 0.00433f
C39228 VPWR.t1517 VGND 0.0298f
C39229 VPWR.t4665 VGND 0.02791f
C39230 VPWR.t1515 VGND 0.04521f
C39231 VPWR.t5483 VGND 0.01172f
C39232 VPWR.t2916 VGND 0.03483f
C39233 VPWR.t2914 VGND 0.04309f
C39234 VPWR.t6155 VGND 0.03248f
C39235 VPWR.t2263 VGND 0.03271f
C39236 VPWR.t5406 VGND 0.04231f
C39237 VPWR.t5223 VGND 0.03271f
C39238 VPWR.t2762 VGND 0.05001f
C39239 VPWR.t991 VGND 0.05001f
C39240 VPWR.t4704 VGND 0.04231f
C39241 VPWR.t1451 VGND 0.0202f
C39242 VPWR.n199 VGND 0.05372f
C39243 VPWR.t4736 VGND 0.00433f
C39244 VPWR.t388 VGND 0.00433f
C39245 VPWR.t4839 VGND 0.00433f
C39246 VPWR.t387 VGND 0.05481f
C39247 VPWR.n200 VGND 0.03642f
C39248 VPWR.t5230 VGND 0.00433f
C39249 VPWR.t5892 VGND 0.00433f
C39250 VPWR.t7122 VGND 0.00433f
C39251 VPWR.t1481 VGND 0.00433f
C39252 VPWR.t3332 VGND 0.00433f
C39253 VPWR.t5729 VGND 0.00433f
C39254 VPWR.t4457 VGND 0.00433f
C39255 VPWR.t812 VGND 0.00433f
C39256 VPWR.t4635 VGND 0.00433f
C39257 VPWR.t4917 VGND 0.00433f
C39258 VPWR.t3027 VGND 0.00433f
C39259 VPWR.t5150 VGND 0.00433f
C39260 VPWR.t386 VGND 0.00433f
C39261 VPWR.t3415 VGND 0.00433f
C39262 VPWR.t2476 VGND 0.00433f
C39263 VPWR.t2996 VGND 0.00433f
C39264 VPWR.t4838 VGND 0.03751f
C39265 VPWR.t5229 VGND 0.05001f
C39266 VPWR.t5891 VGND 0.05001f
C39267 VPWR.t7121 VGND 0.05001f
C39268 VPWR.t1480 VGND 0.05001f
C39269 VPWR.t3331 VGND 0.05001f
C39270 VPWR.t5728 VGND 0.05001f
C39271 VPWR.t4456 VGND 0.05001f
C39272 VPWR.t811 VGND 0.05001f
C39273 VPWR.t4634 VGND 0.05001f
C39274 VPWR.t4916 VGND 0.05001f
C39275 VPWR.t3026 VGND 0.05001f
C39276 VPWR.t5149 VGND 0.05001f
C39277 VPWR.t385 VGND 0.05001f
C39278 VPWR.t3414 VGND 0.05001f
C39279 VPWR.t2475 VGND 0.04231f
C39280 VPWR.t2995 VGND 0.0202f
C39281 VPWR.n201 VGND 0.05372f
C39282 VPWR.t1807 VGND 0.00433f
C39283 VPWR.t3080 VGND 0.00433f
C39284 VPWR.t5554 VGND 0.00433f
C39285 VPWR.t4853 VGND 0.00433f
C39286 VPWR.t1632 VGND 0.00433f
C39287 VPWR.t4731 VGND 0.00433f
C39288 VPWR.t1510 VGND 0.00433f
C39289 VPWR.t2421 VGND 0.00433f
C39290 VPWR.t1560 VGND 0.00433f
C39291 VPWR.t5543 VGND 0.00433f
C39292 VPWR.t4942 VGND 0.00433f
C39293 VPWR.t4306 VGND 0.00433f
C39294 VPWR.t4139 VGND 0.00433f
C39295 VPWR.t67 VGND 0.00433f
C39296 VPWR.t521 VGND 0.00433f
C39297 VPWR.t1806 VGND 0.08751f
C39298 VPWR.t4852 VGND 0.10001f
C39299 VPWR.t1631 VGND 0.10001f
C39300 VPWR.t1509 VGND 0.10001f
C39301 VPWR.t1559 VGND 0.10001f
C39302 VPWR.t4305 VGND 0.10001f
C39303 VPWR.t66 VGND 0.06731f
C39304 VPWR.n202 VGND 0.03642f
C39305 VPWR.t3657 VGND 0.00433f
C39306 VPWR.t520 VGND 0.0298f
C39307 VPWR.t3656 VGND 0.0202f
C39308 VPWR.n203 VGND 0.02102f
C39309 VPWR.t1148 VGND 0.00433f
C39310 VPWR.t4002 VGND 0.00433f
C39311 VPWR.t3641 VGND 0.00433f
C39312 VPWR.t5310 VGND 0.00433f
C39313 VPWR.t6135 VGND 0.00433f
C39314 VPWR.t1895 VGND 0.00433f
C39315 VPWR.t4356 VGND 0.00433f
C39316 VPWR.t3704 VGND 0.00433f
C39317 VPWR.t2722 VGND 0.00433f
C39318 VPWR.t700 VGND 0.00433f
C39319 VPWR.t2220 VGND 0.00433f
C39320 VPWR.t451 VGND 0.00433f
C39321 VPWR.t5031 VGND 0.00433f
C39322 VPWR.t5064 VGND 0.00433f
C39323 VPWR.t424 VGND 0.00433f
C39324 VPWR.t3648 VGND 0.00433f
C39325 VPWR.t2926 VGND 0.00433f
C39326 VPWR.t1147 VGND 0.08271f
C39327 VPWR.t3640 VGND 0.10001f
C39328 VPWR.t1894 VGND 0.10001f
C39329 VPWR.t3703 VGND 0.10001f
C39330 VPWR.t699 VGND 0.10001f
C39331 VPWR.t450 VGND 0.10001f
C39332 VPWR.t5030 VGND 0.10001f
C39333 VPWR.t423 VGND 0.06731f
C39334 VPWR.n204 VGND 0.03642f
C39335 VPWR.t2645 VGND 0.00433f
C39336 VPWR.t4319 VGND 0.00433f
C39337 VPWR.t1416 VGND 0.00433f
C39338 VPWR.t2434 VGND 0.00433f
C39339 VPWR.t5042 VGND 0.00433f
C39340 VPWR.t3719 VGND 0.00433f
C39341 VPWR.t2845 VGND 0.00433f
C39342 VPWR.t2053 VGND 0.00433f
C39343 VPWR.t828 VGND 0.00433f
C39344 VPWR.t2712 VGND 0.00433f
C39345 VPWR.t1305 VGND 0.00433f
C39346 VPWR.t2374 VGND 0.00433f
C39347 VPWR.t5383 VGND 0.00433f
C39348 VPWR.t2633 VGND 0.00433f
C39349 VPWR.t5167 VGND 0.00433f
C39350 VPWR.t2925 VGND 0.03751f
C39351 VPWR.t2644 VGND 0.05001f
C39352 VPWR.t4318 VGND 0.05001f
C39353 VPWR.t1415 VGND 0.05001f
C39354 VPWR.t2433 VGND 0.05001f
C39355 VPWR.t5041 VGND 0.05001f
C39356 VPWR.t3718 VGND 0.05001f
C39357 VPWR.t2844 VGND 0.05001f
C39358 VPWR.t2052 VGND 0.05001f
C39359 VPWR.t827 VGND 0.05001f
C39360 VPWR.t2711 VGND 0.05001f
C39361 VPWR.t1304 VGND 0.05001f
C39362 VPWR.t2373 VGND 0.05001f
C39363 VPWR.t5382 VGND 0.05001f
C39364 VPWR.t2632 VGND 0.04231f
C39365 VPWR.t5166 VGND 0.0202f
C39366 VPWR.n205 VGND 0.02102f
C39367 VPWR.t3768 VGND 0.00433f
C39368 VPWR.n206 VGND 0.03642f
C39369 VPWR.t3653 VGND 0.00433f
C39370 VPWR.t1650 VGND 0.00433f
C39371 VPWR.t611 VGND 0.00433f
C39372 VPWR.t3885 VGND 0.00433f
C39373 VPWR.t4394 VGND 0.00433f
C39374 VPWR.t5773 VGND 0.00433f
C39375 VPWR.t4925 VGND 0.00433f
C39376 VPWR.t1566 VGND 0.00433f
C39377 VPWR.t2847 VGND 0.00433f
C39378 VPWR.t5069 VGND 0.00433f
C39379 VPWR.t1534 VGND 0.00433f
C39380 VPWR.t5377 VGND 0.00433f
C39381 VPWR.t3706 VGND 0.00433f
C39382 VPWR.t1967 VGND 0.00433f
C39383 VPWR.t5105 VGND 0.00433f
C39384 VPWR.t5964 VGND 0.00433f
C39385 VPWR.t3767 VGND 0.0298f
C39386 VPWR.t3652 VGND 0.03271f
C39387 VPWR.t1649 VGND 0.05001f
C39388 VPWR.t610 VGND 0.05001f
C39389 VPWR.t3884 VGND 0.05001f
C39390 VPWR.t4393 VGND 0.05001f
C39391 VPWR.t5772 VGND 0.05001f
C39392 VPWR.t4924 VGND 0.05001f
C39393 VPWR.t1565 VGND 0.05001f
C39394 VPWR.t2846 VGND 0.05001f
C39395 VPWR.t5068 VGND 0.05001f
C39396 VPWR.t1533 VGND 0.05001f
C39397 VPWR.t5376 VGND 0.05001f
C39398 VPWR.t3705 VGND 0.05001f
C39399 VPWR.t1966 VGND 0.05001f
C39400 VPWR.t5104 VGND 0.04231f
C39401 VPWR.t5963 VGND 0.0202f
C39402 VPWR.n207 VGND 0.05372f
C39403 VPWR.t2012 VGND 0.00433f
C39404 VPWR.t3602 VGND 0.00433f
C39405 VPWR.t1347 VGND 0.00433f
C39406 VPWR.t3427 VGND 0.00433f
C39407 VPWR.t3197 VGND 0.00433f
C39408 VPWR.t1969 VGND 0.00433f
C39409 VPWR.t4257 VGND 0.00433f
C39410 VPWR.t3952 VGND 0.00433f
C39411 VPWR.t2981 VGND 0.00433f
C39412 VPWR.t1975 VGND 0.00433f
C39413 VPWR.t1496 VGND 0.00433f
C39414 VPWR.t7142 VGND 0.00433f
C39415 VPWR.t4271 VGND 0.00433f
C39416 VPWR.t1570 VGND 0.00433f
C39417 VPWR.t1544 VGND 0.00433f
C39418 VPWR.t2131 VGND 0.00433f
C39419 VPWR.t2011 VGND 0.08751f
C39420 VPWR.t1346 VGND 0.10001f
C39421 VPWR.t1968 VGND 0.10001f
C39422 VPWR.t3951 VGND 0.10001f
C39423 VPWR.t1974 VGND 0.10001f
C39424 VPWR.t1495 VGND 0.10001f
C39425 VPWR.t1569 VGND 0.10001f
C39426 VPWR.t1543 VGND 0.06731f
C39427 VPWR.n208 VGND 0.02233f
C39428 VPWR.n209 VGND 0.02171f
C39429 VPWR.n210 VGND 0.02171f
C39430 VPWR.n211 VGND 0.01577f
C39431 VPWR.n212 VGND 0.0207f
C39432 VPWR.n213 VGND 0.02171f
C39433 VPWR.n214 VGND 0.02171f
C39434 VPWR.n215 VGND 0.01568f
C39435 VPWR.n216 VGND 0.01097f
C39436 VPWR.n217 VGND 0.01144f
C39437 VPWR.n218 VGND 0.00986f
C39438 VPWR.n219 VGND 0.0083f
C39439 VPWR.n220 VGND 0.00837f
C39440 VPWR.n221 VGND 0.01085f
C39441 VPWR.n222 VGND 0.01085f
C39442 VPWR.n223 VGND 0.01085f
C39443 VPWR.n224 VGND 0.01085f
C39444 VPWR.n225 VGND 0.00839f
C39445 VPWR.n226 VGND 0.00985f
C39446 VPWR.n227 VGND 0.01085f
C39447 VPWR.n228 VGND 0.01085f
C39448 VPWR.n229 VGND 0.01085f
C39449 VPWR.n230 VGND 0.01085f
C39450 VPWR.n231 VGND 0.01085f
C39451 VPWR.n232 VGND 0.01085f
C39452 VPWR.n233 VGND 0.0085f
C39453 VPWR.n234 VGND 0.01077f
C39454 VPWR.n235 VGND 0.00735f
C39455 VPWR.n236 VGND 0.01189f
C39456 VPWR.n237 VGND 0.01144f
C39457 VPWR.n238 VGND 0.01085f
C39458 VPWR.n239 VGND 0.01085f
C39459 VPWR.n240 VGND 0.01085f
C39460 VPWR.n241 VGND 0.01085f
C39461 VPWR.n242 VGND 0.01085f
C39462 VPWR.n243 VGND 0.00839f
C39463 VPWR.n244 VGND 0.00985f
C39464 VPWR.n245 VGND 0.01085f
C39465 VPWR.n246 VGND 0.01085f
C39466 VPWR.n247 VGND 0.01085f
C39467 VPWR.n248 VGND 0.01085f
C39468 VPWR.n249 VGND 0.01085f
C39469 VPWR.n250 VGND 0.01085f
C39470 VPWR.n251 VGND 0.01023f
C39471 VPWR.n252 VGND 0.01189f
C39472 VPWR.n253 VGND 0.00541f
C39473 VPWR.n254 VGND 0.01878f
C39474 VPWR.n255 VGND 0.10419f
C39475 VPWR.t4789 VGND 0.00433f
C39476 VPWR.n256 VGND 0.01634f
C39477 VPWR.t5130 VGND 0.00433f
C39478 VPWR.t5854 VGND 0.00433f
C39479 VPWR.t5691 VGND 0.00433f
C39480 VPWR.t3320 VGND 0.00433f
C39481 VPWR.t4289 VGND 0.00433f
C39482 VPWR.t1572 VGND 0.00433f
C39483 VPWR.t1963 VGND 0.00433f
C39484 VPWR.t6014 VGND 0.00433f
C39485 VPWR.t5129 VGND 0.04035f
C39486 VPWR.t5853 VGND 0.05996f
C39487 VPWR.t5690 VGND 0.05996f
C39488 VPWR.t3319 VGND 0.05996f
C39489 VPWR.t4288 VGND 0.05996f
C39490 VPWR.t1571 VGND 0.05996f
C39491 VPWR.t1962 VGND 0.05996f
C39492 VPWR.t6013 VGND 0.05247f
C39493 VPWR.n257 VGND 0.03832f
C39494 VPWR.t6323 VGND 0.00433f
C39495 VPWR.n258 VGND 0.01389f
C39496 VPWR.n259 VGND 0.32859f
C39497 VPWR.t4416 VGND 0.00433f
C39498 VPWR.n260 VGND 0.01042f
C39499 VPWR.t1724 VGND 0.00433f
C39500 VPWR.t1780 VGND 0.00433f
C39501 VPWR.t3613 VGND 0.00433f
C39502 VPWR.t2946 VGND 0.00433f
C39503 VPWR.t5474 VGND 0.00433f
C39504 VPWR.t2937 VGND 0.00433f
C39505 VPWR.t2887 VGND 0.00433f
C39506 VPWR.t2686 VGND 0.00433f
C39507 VPWR.t2945 VGND 0.06731f
C39508 VPWR.t2936 VGND 0.08271f
C39509 VPWR.t2685 VGND 0.05481f
C39510 VPWR.n261 VGND 0.05372f
C39511 VPWR.t2139 VGND 0.00433f
C39512 VPWR.t532 VGND 0.00433f
C39513 VPWR.t4104 VGND 0.00433f
C39514 VPWR.t4949 VGND 0.00433f
C39515 VPWR.t4166 VGND 0.00433f
C39516 VPWR.t3905 VGND 0.00433f
C39517 VPWR.t5330 VGND 0.00433f
C39518 VPWR.t4440 VGND 0.00433f
C39519 VPWR.t1376 VGND 0.00433f
C39520 VPWR.t2138 VGND 0.0202f
C39521 VPWR.t531 VGND 0.04231f
C39522 VPWR.t4103 VGND 0.05001f
C39523 VPWR.t4948 VGND 0.05001f
C39524 VPWR.t4165 VGND 0.05001f
C39525 VPWR.t3904 VGND 0.05001f
C39526 VPWR.t5329 VGND 0.05001f
C39527 VPWR.t4439 VGND 0.05001f
C39528 VPWR.t1375 VGND 0.05001f
C39529 VPWR.t4618 VGND 0.03751f
C39530 VPWR.n262 VGND 0.03642f
C39531 VPWR.t4619 VGND 0.00433f
C39532 VPWR.t915 VGND 0.00433f
C39533 VPWR.t1236 VGND 0.00433f
C39534 VPWR.n263 VGND 0.01535f
C39535 VPWR.n264 VGND 0.32859f
C39536 VPWR.t868 VGND 0.00433f
C39537 VPWR.n265 VGND 0.01144f
C39538 VPWR.t3384 VGND 0.00433f
C39539 VPWR.t65 VGND 0.00433f
C39540 VPWR.t2668 VGND 0.00433f
C39541 VPWR.t4198 VGND 0.00433f
C39542 VPWR.t2975 VGND 0.00433f
C39543 VPWR.t3383 VGND 0.04035f
C39544 VPWR.t64 VGND 0.05996f
C39545 VPWR.t2667 VGND 0.05996f
C39546 VPWR.t4197 VGND 0.05996f
C39547 VPWR.t2974 VGND 0.05334f
C39548 VPWR.n266 VGND 0.05473f
C39549 VPWR.t846 VGND 0.00433f
C39550 VPWR.t6148 VGND 0.00433f
C39551 VPWR.t5033 VGND 0.00433f
C39552 VPWR.t307 VGND 0.00433f
C39553 VPWR.t773 VGND 0.00433f
C39554 VPWR.t845 VGND 0.02065f
C39555 VPWR.t6147 VGND 0.04231f
C39556 VPWR.t5032 VGND 0.05001f
C39557 VPWR.t306 VGND 0.05001f
C39558 VPWR.t772 VGND 0.05001f
C39559 VPWR.t3894 VGND 0.03751f
C39560 VPWR.n267 VGND 0.03642f
C39561 VPWR.t3895 VGND 0.00433f
C39562 VPWR.t4191 VGND 0.00433f
C39563 VPWR.t863 VGND 0.00433f
C39564 VPWR.t5983 VGND 0.00433f
C39565 VPWR.t5245 VGND 0.00433f
C39566 VPWR.t2510 VGND 0.00433f
C39567 VPWR.t3013 VGND 0.00433f
C39568 VPWR.t5882 VGND 0.00433f
C39569 VPWR.t690 VGND 0.00433f
C39570 VPWR.t1176 VGND 0.00433f
C39571 VPWR.t6360 VGND 0.00433f
C39572 VPWR.t4230 VGND 0.00433f
C39573 VPWR.t1433 VGND 0.00433f
C39574 VPWR.t862 VGND 0.06731f
C39575 VPWR.t5244 VGND 0.10001f
C39576 VPWR.t2509 VGND 0.10001f
C39577 VPWR.t689 VGND 0.08271f
C39578 VPWR.t1175 VGND 0.05001f
C39579 VPWR.t1432 VGND 0.05001f
C39580 VPWR.n268 VGND 0.01214f
C39581 VPWR.n269 VGND 0.01588f
C39582 VPWR.n270 VGND 0.02171f
C39583 VPWR.n271 VGND 0.02059f
C39584 VPWR.n272 VGND 0.01402f
C39585 VPWR.n273 VGND 0.13412f
C39586 VPWR.t3452 VGND 0.00433f
C39587 VPWR.n274 VGND 0.01073f
C39588 VPWR.t830 VGND 0.00433f
C39589 VPWR.t3948 VGND 0.00433f
C39590 VPWR.t4641 VGND 0.00433f
C39591 VPWR.t2061 VGND 0.00433f
C39592 VPWR.t3050 VGND 0.00433f
C39593 VPWR.t2450 VGND 0.00433f
C39594 VPWR.t3551 VGND 0.00433f
C39595 VPWR.t3032 VGND 0.00433f
C39596 VPWR.t1671 VGND 0.00433f
C39597 VPWR.t6084 VGND 0.00433f
C39598 VPWR.t2924 VGND 0.00433f
C39599 VPWR.t1250 VGND 0.00433f
C39600 VPWR.t5669 VGND 0.00433f
C39601 VPWR.t473 VGND 0.00433f
C39602 VPWR.t3380 VGND 0.00433f
C39603 VPWR.n275 VGND 0.01013f
C39604 VPWR.n276 VGND 0.00985f
C39605 VPWR.n277 VGND 0.01085f
C39606 VPWR.n278 VGND 0.01085f
C39607 VPWR.n279 VGND 0.01085f
C39608 VPWR.n280 VGND 0.01085f
C39609 VPWR.n281 VGND 0.01085f
C39610 VPWR.n282 VGND 0.00834f
C39611 VPWR.n283 VGND 0.00665f
C39612 VPWR.t3550 VGND 0.025f
C39613 VPWR.t3031 VGND 0.04521f
C39614 VPWR.t1670 VGND 0.05001f
C39615 VPWR.t6083 VGND 0.05001f
C39616 VPWR.t2923 VGND 0.05001f
C39617 VPWR.t1249 VGND 0.05001f
C39618 VPWR.t5668 VGND 0.05001f
C39619 VPWR.t472 VGND 0.05001f
C39620 VPWR.t3379 VGND 0.05001f
C39621 VPWR.t3451 VGND 0.05001f
C39622 VPWR.t829 VGND 0.05001f
C39623 VPWR.t3947 VGND 0.05001f
C39624 VPWR.t4640 VGND 0.05001f
C39625 VPWR.t2060 VGND 0.05001f
C39626 VPWR.t3049 VGND 0.0298f
C39627 VPWR.t2449 VGND 0.06143f
C39628 VPWR.t499 VGND 0.00433f
C39629 VPWR.t4857 VGND 0.00433f
C39630 VPWR.t7141 VGND 0.00433f
C39631 VPWR.t493 VGND 0.00433f
C39632 VPWR.t7086 VGND 0.00433f
C39633 VPWR.t3856 VGND 0.00433f
C39634 VPWR.t392 VGND 0.00433f
C39635 VPWR.t1195 VGND 0.00433f
C39636 VPWR.t4930 VGND 0.00433f
C39637 VPWR.t1926 VGND 0.00433f
C39638 VPWR.t5956 VGND 0.00433f
C39639 VPWR.t2193 VGND 0.00433f
C39640 VPWR.t2230 VGND 0.00433f
C39641 VPWR.t4544 VGND 0.00433f
C39642 VPWR.t2408 VGND 0.00433f
C39643 VPWR.t6056 VGND 0.00433f
C39644 VPWR.t5108 VGND 0.00433f
C39645 VPWR.t498 VGND 0.05001f
C39646 VPWR.t4856 VGND 0.0173f
C39647 VPWR.t7140 VGND 0.04521f
C39648 VPWR.t492 VGND 0.05001f
C39649 VPWR.t7085 VGND 0.05001f
C39650 VPWR.t3855 VGND 0.05001f
C39651 VPWR.t391 VGND 0.05001f
C39652 VPWR.t1194 VGND 0.05001f
C39653 VPWR.t4929 VGND 0.05001f
C39654 VPWR.t1925 VGND 0.05001f
C39655 VPWR.t5955 VGND 0.05001f
C39656 VPWR.t2192 VGND 0.05001f
C39657 VPWR.t2229 VGND 0.05001f
C39658 VPWR.t4543 VGND 0.05001f
C39659 VPWR.t2407 VGND 0.05001f
C39660 VPWR.t6055 VGND 0.0298f
C39661 VPWR.t5107 VGND 0.06143f
C39662 VPWR.t1418 VGND 0.00433f
C39663 VPWR.t2798 VGND 0.00433f
C39664 VPWR.t3177 VGND 0.00433f
C39665 VPWR.t7124 VGND 0.00433f
C39666 VPWR.t3467 VGND 0.00433f
C39667 VPWR.t3334 VGND 0.00433f
C39668 VPWR.t4807 VGND 0.00433f
C39669 VPWR.t4459 VGND 0.00433f
C39670 VPWR.t5360 VGND 0.00433f
C39671 VPWR.t4637 VGND 0.00433f
C39672 VPWR.t4595 VGND 0.00433f
C39673 VPWR.t2250 VGND 0.00433f
C39674 VPWR.n284 VGND 0.01027f
C39675 VPWR.t745 VGND 0.00433f
C39676 VPWR.n285 VGND 0.00971f
C39677 VPWR.t3589 VGND 0.00433f
C39678 VPWR.t6110 VGND 0.00433f
C39679 VPWR.t3214 VGND 0.00433f
C39680 VPWR.t5061 VGND 0.00433f
C39681 VPWR.t3545 VGND 0.00433f
C39682 VPWR.t3627 VGND 0.00433f
C39683 VPWR.t5542 VGND 0.00433f
C39684 VPWR.t4654 VGND 0.00433f
C39685 VPWR.t4254 VGND 0.00433f
C39686 VPWR.t4815 VGND 0.00433f
C39687 VPWR.t945 VGND 0.00433f
C39688 VPWR.t3887 VGND 0.00433f
C39689 VPWR.t4941 VGND 0.00433f
C39690 VPWR.t5453 VGND 0.00433f
C39691 VPWR.t3365 VGND 0.00433f
C39692 VPWR.t2494 VGND 0.00433f
C39693 VPWR.t3775 VGND 0.00433f
C39694 VPWR.t2472 VGND 0.00433f
C39695 VPWR.t783 VGND 0.00433f
C39696 VPWR.t3816 VGND 0.00433f
C39697 VPWR.t3854 VGND 0.00433f
C39698 VPWR.t4447 VGND 0.00433f
C39699 VPWR.t3094 VGND 0.00433f
C39700 VPWR.t4653 VGND 0.0298f
C39701 VPWR.t4253 VGND 0.05001f
C39702 VPWR.t4814 VGND 0.05001f
C39703 VPWR.t944 VGND 0.05001f
C39704 VPWR.t3886 VGND 0.05001f
C39705 VPWR.t4940 VGND 0.05001f
C39706 VPWR.t5452 VGND 0.05001f
C39707 VPWR.t3364 VGND 0.05001f
C39708 VPWR.t2493 VGND 0.05001f
C39709 VPWR.t3774 VGND 0.05001f
C39710 VPWR.t2471 VGND 0.05001f
C39711 VPWR.t782 VGND 0.05001f
C39712 VPWR.t3815 VGND 0.05001f
C39713 VPWR.t3853 VGND 0.04521f
C39714 VPWR.t4446 VGND 0.0173f
C39715 VPWR.t3093 VGND 0.05001f
C39716 VPWR.t3190 VGND 0.06143f
C39717 VPWR.t3191 VGND 0.00433f
C39718 VPWR.t5852 VGND 0.00433f
C39719 VPWR.t4767 VGND 0.00433f
C39720 VPWR.t1090 VGND 0.00433f
C39721 VPWR.t2201 VGND 0.00433f
C39722 VPWR.t2889 VGND 0.00433f
C39723 VPWR.t4759 VGND 0.00433f
C39724 VPWR.t5841 VGND 0.00433f
C39725 VPWR.t5037 VGND 0.00433f
C39726 VPWR.t1008 VGND 0.00433f
C39727 VPWR.t1229 VGND 0.00433f
C39728 VPWR.t2133 VGND 0.00433f
C39729 VPWR.t1707 VGND 0.00433f
C39730 VPWR.t4190 VGND 0.00433f
C39731 VPWR.t1646 VGND 0.00433f
C39732 VPWR.t3318 VGND 0.00433f
C39733 VPWR.t5851 VGND 0.0298f
C39734 VPWR.t4766 VGND 0.05001f
C39735 VPWR.t1089 VGND 0.05001f
C39736 VPWR.t2200 VGND 0.05001f
C39737 VPWR.t2888 VGND 0.05001f
C39738 VPWR.t4758 VGND 0.05001f
C39739 VPWR.t5840 VGND 0.05001f
C39740 VPWR.t5036 VGND 0.05001f
C39741 VPWR.t1007 VGND 0.05001f
C39742 VPWR.t1228 VGND 0.05001f
C39743 VPWR.t2132 VGND 0.05001f
C39744 VPWR.t1706 VGND 0.05001f
C39745 VPWR.t4189 VGND 0.05001f
C39746 VPWR.t1645 VGND 0.04521f
C39747 VPWR.t3317 VGND 0.025f
C39748 VPWR.n286 VGND 0.00665f
C39749 VPWR.n287 VGND 0.00834f
C39750 VPWR.n288 VGND 0.01085f
C39751 VPWR.n289 VGND 0.01085f
C39752 VPWR.n290 VGND 0.01085f
C39753 VPWR.n291 VGND 0.01085f
C39754 VPWR.n292 VGND 0.01085f
C39755 VPWR.n293 VGND 0.00985f
C39756 VPWR.n294 VGND 0.01013f
C39757 VPWR.n295 VGND 0.01073f
C39758 VPWR.n296 VGND 0.00656f
C39759 VPWR.n297 VGND 0.00924f
C39760 VPWR.n298 VGND 0.01085f
C39761 VPWR.n299 VGND 0.01085f
C39762 VPWR.n300 VGND 0.01085f
C39763 VPWR.n301 VGND 0.01085f
C39764 VPWR.n302 VGND 0.01144f
C39765 VPWR.n303 VGND 0.01189f
C39766 VPWR.n304 VGND 0.00758f
C39767 VPWR.n305 VGND 0.00544f
C39768 VPWR.n306 VGND 0.01023f
C39769 VPWR.n307 VGND 0.01085f
C39770 VPWR.n308 VGND 0.01085f
C39771 VPWR.n309 VGND 0.01085f
C39772 VPWR.n310 VGND 0.01085f
C39773 VPWR.n311 VGND 0.01085f
C39774 VPWR.n312 VGND 0.01085f
C39775 VPWR.n313 VGND 0.01085f
C39776 VPWR.n314 VGND 0.01085f
C39777 VPWR.n315 VGND 0.01085f
C39778 VPWR.n316 VGND 0.01085f
C39779 VPWR.n317 VGND 0.01085f
C39780 VPWR.n318 VGND 0.01085f
C39781 VPWR.n319 VGND 0.01085f
C39782 VPWR.n320 VGND 0.01144f
C39783 VPWR.t1766 VGND 0.00433f
C39784 VPWR.t5173 VGND 0.00433f
C39785 VPWR.t4298 VGND 0.00433f
C39786 VPWR.t6151 VGND 0.00433f
C39787 VPWR.t4862 VGND 0.00433f
C39788 VPWR.t5482 VGND 0.00433f
C39789 VPWR.t4707 VGND 0.00433f
C39790 VPWR.t2057 VGND 0.00433f
C39791 VPWR.t2213 VGND 0.00433f
C39792 VPWR.t1422 VGND 0.00433f
C39793 VPWR.n321 VGND 0.01085f
C39794 VPWR.n322 VGND 0.01085f
C39795 VPWR.n323 VGND 0.01085f
C39796 VPWR.n324 VGND 0.01085f
C39797 VPWR.n325 VGND 0.01085f
C39798 VPWR.n326 VGND 0.01085f
C39799 VPWR.n327 VGND 0.01085f
C39800 VPWR.n328 VGND 0.01023f
C39801 VPWR.n329 VGND 0.00544f
C39802 VPWR.n330 VGND 0.00758f
C39803 VPWR.n331 VGND 0.01189f
C39804 VPWR.t5541 VGND 0.06143f
C39805 VPWR.t1765 VGND 0.05001f
C39806 VPWR.t5172 VGND 0.0173f
C39807 VPWR.t4297 VGND 0.04521f
C39808 VPWR.t6150 VGND 0.05001f
C39809 VPWR.t4861 VGND 0.05001f
C39810 VPWR.t5481 VGND 0.05001f
C39811 VPWR.t4706 VGND 0.05001f
C39812 VPWR.t2056 VGND 0.05001f
C39813 VPWR.t2212 VGND 0.05001f
C39814 VPWR.t1421 VGND 0.05001f
C39815 VPWR.t744 VGND 0.05001f
C39816 VPWR.t3588 VGND 0.05001f
C39817 VPWR.t6109 VGND 0.05001f
C39818 VPWR.t3213 VGND 0.05001f
C39819 VPWR.t5060 VGND 0.05001f
C39820 VPWR.t3544 VGND 0.0298f
C39821 VPWR.t3626 VGND 0.06143f
C39822 VPWR.t4009 VGND 0.00433f
C39823 VPWR.t4513 VGND 0.00433f
C39824 VPWR.t6089 VGND 0.00433f
C39825 VPWR.t3597 VGND 0.00433f
C39826 VPWR.t5631 VGND 0.00433f
C39827 VPWR.t4590 VGND 0.00433f
C39828 VPWR.t4352 VGND 0.00433f
C39829 VPWR.t4455 VGND 0.00433f
C39830 VPWR.t6219 VGND 0.00433f
C39831 VPWR.t6209 VGND 0.00433f
C39832 VPWR.t61 VGND 0.00433f
C39833 VPWR.t3808 VGND 0.00433f
C39834 VPWR.t3726 VGND 0.00433f
C39835 VPWR.t4025 VGND 0.00433f
C39836 VPWR.t1655 VGND 0.00433f
C39837 VPWR.t1466 VGND 0.00433f
C39838 VPWR.t4526 VGND 0.00433f
C39839 VPWR.t4008 VGND 0.05001f
C39840 VPWR.t4512 VGND 0.0173f
C39841 VPWR.t6088 VGND 0.04521f
C39842 VPWR.t3596 VGND 0.05001f
C39843 VPWR.t5630 VGND 0.05001f
C39844 VPWR.t4589 VGND 0.05001f
C39845 VPWR.t4351 VGND 0.05001f
C39846 VPWR.t4454 VGND 0.05001f
C39847 VPWR.t6218 VGND 0.05001f
C39848 VPWR.t6208 VGND 0.05001f
C39849 VPWR.t60 VGND 0.05001f
C39850 VPWR.t3807 VGND 0.05001f
C39851 VPWR.t3725 VGND 0.05001f
C39852 VPWR.t4024 VGND 0.05001f
C39853 VPWR.t1654 VGND 0.05001f
C39854 VPWR.t1465 VGND 0.0298f
C39855 VPWR.t4525 VGND 0.06143f
C39856 VPWR.t3818 VGND 0.00433f
C39857 VPWR.t4915 VGND 0.00433f
C39858 VPWR.t489 VGND 0.00433f
C39859 VPWR.t676 VGND 0.00433f
C39860 VPWR.t2627 VGND 0.00433f
C39861 VPWR.t4875 VGND 0.00433f
C39862 VPWR.t6192 VGND 0.00433f
C39863 VPWR.t3354 VGND 0.00433f
C39864 VPWR.t4491 VGND 0.00433f
C39865 VPWR.t6054 VGND 0.00433f
C39866 VPWR.t4615 VGND 0.00433f
C39867 VPWR.t3169 VGND 0.00433f
C39868 VPWR.t4152 VGND 0.00433f
C39869 VPWR.t5273 VGND 0.00433f
C39870 VPWR.t1854 VGND 0.00433f
C39871 VPWR.t2842 VGND 0.00433f
C39872 VPWR.t1562 VGND 0.00433f
C39873 VPWR.t3817 VGND 0.05001f
C39874 VPWR.t4914 VGND 0.0173f
C39875 VPWR.t488 VGND 0.04521f
C39876 VPWR.t675 VGND 0.05001f
C39877 VPWR.t2626 VGND 0.05001f
C39878 VPWR.t4874 VGND 0.05001f
C39879 VPWR.t6191 VGND 0.05001f
C39880 VPWR.t3353 VGND 0.05001f
C39881 VPWR.t4490 VGND 0.05001f
C39882 VPWR.t6053 VGND 0.05001f
C39883 VPWR.t4614 VGND 0.05001f
C39884 VPWR.t3168 VGND 0.05001f
C39885 VPWR.t4151 VGND 0.05001f
C39886 VPWR.t5272 VGND 0.05001f
C39887 VPWR.t1853 VGND 0.05001f
C39888 VPWR.t2841 VGND 0.0298f
C39889 VPWR.t1561 VGND 0.04122f
C39890 VPWR.t581 VGND 0.00433f
C39891 VPWR.t1914 VGND 0.00433f
C39892 VPWR.t4101 VGND 0.00433f
C39893 VPWR.t5451 VGND 0.00433f
C39894 VPWR.t3109 VGND 0.00433f
C39895 VPWR.t1392 VGND 0.00433f
C39896 VPWR.t1336 VGND 0.00433f
C39897 VPWR.t3079 VGND 0.00433f
C39898 VPWR.t2528 VGND 0.00433f
C39899 VPWR.t6326 VGND 0.00433f
C39900 VPWR.t4575 VGND 0.00433f
C39901 VPWR.t3386 VGND 0.00433f
C39902 VPWR.t3981 VGND 0.00433f
C39903 VPWR.t5742 VGND 0.00433f
C39904 VPWR.t5647 VGND 0.00433f
C39905 VPWR.t3903 VGND 0.00433f
C39906 VPWR.t580 VGND 0.08271f
C39907 VPWR.t4100 VGND 0.10001f
C39908 VPWR.t1391 VGND 0.10001f
C39909 VPWR.t1335 VGND 0.10001f
C39910 VPWR.t2527 VGND 0.10001f
C39911 VPWR.t3385 VGND 0.10001f
C39912 VPWR.t3980 VGND 0.10001f
C39913 VPWR.t3902 VGND 0.06731f
C39914 VPWR.n332 VGND 0.02233f
C39915 VPWR.n333 VGND 0.02171f
C39916 VPWR.n334 VGND 0.02171f
C39917 VPWR.n335 VGND 0.01577f
C39918 VPWR.n336 VGND 0.0207f
C39919 VPWR.n337 VGND 0.02171f
C39920 VPWR.n338 VGND 0.02171f
C39921 VPWR.n339 VGND 0.01568f
C39922 VPWR.n340 VGND 0.01165f
C39923 VPWR.n341 VGND 0.01144f
C39924 VPWR.n342 VGND 0.01085f
C39925 VPWR.n343 VGND 0.01085f
C39926 VPWR.n344 VGND 0.01085f
C39927 VPWR.n345 VGND 0.01085f
C39928 VPWR.n346 VGND 0.01085f
C39929 VPWR.n347 VGND 0.00608f
C39930 VPWR.t4354 VGND 0.00433f
C39931 VPWR.n348 VGND 0.01042f
C39932 VPWR.t4546 VGND 0.00433f
C39933 VPWR.t682 VGND 0.00433f
C39934 VPWR.t5725 VGND 0.00433f
C39935 VPWR.t1475 VGND 0.00433f
C39936 VPWR.t6160 VGND 0.00433f
C39937 VPWR.t4396 VGND 0.00433f
C39938 VPWR.t3618 VGND 0.00433f
C39939 VPWR.t428 VGND 0.00433f
C39940 VPWR.t3929 VGND 0.00433f
C39941 VPWR.t3263 VGND 0.00433f
C39942 VPWR.t1845 VGND 0.00433f
C39943 VPWR.t4032 VGND 0.00433f
C39944 VPWR.t4163 VGND 0.00433f
C39945 VPWR.t3247 VGND 0.00433f
C39946 VPWR.t5771 VGND 0.00433f
C39947 VPWR.t4362 VGND 0.00433f
C39948 VPWR.t459 VGND 0.00433f
C39949 VPWR.t1279 VGND 0.00433f
C39950 VPWR.t4919 VGND 0.00433f
C39951 VPWR.t1450 VGND 0.00433f
C39952 VPWR.t3226 VGND 0.00433f
C39953 VPWR.t2270 VGND 0.00433f
C39954 VPWR.t5979 VGND 0.00433f
C39955 VPWR.t2715 VGND 0.00433f
C39956 VPWR.t3928 VGND 0.0298f
C39957 VPWR.t3262 VGND 0.05001f
C39958 VPWR.t1844 VGND 0.05001f
C39959 VPWR.t4031 VGND 0.05001f
C39960 VPWR.t4162 VGND 0.05001f
C39961 VPWR.t3246 VGND 0.05001f
C39962 VPWR.t5770 VGND 0.05001f
C39963 VPWR.t4361 VGND 0.05001f
C39964 VPWR.t458 VGND 0.05001f
C39965 VPWR.t1278 VGND 0.05001f
C39966 VPWR.t4918 VGND 0.05001f
C39967 VPWR.t1449 VGND 0.05001f
C39968 VPWR.t3225 VGND 0.05001f
C39969 VPWR.t2269 VGND 0.04521f
C39970 VPWR.t5978 VGND 0.0173f
C39971 VPWR.t2714 VGND 0.03271f
C39972 VPWR.t496 VGND 0.04122f
C39973 VPWR.t497 VGND 0.00433f
C39974 VPWR.t3232 VGND 0.00433f
C39975 VPWR.t2145 VGND 0.00433f
C39976 VPWR.t5822 VGND 0.00433f
C39977 VPWR.t4019 VGND 0.00433f
C39978 VPWR.t5604 VGND 0.00473f
C39979 VPWR.t1072 VGND 0.00433f
C39980 VPWR.t5602 VGND 0.00427f
C39981 VPWR.t6039 VGND 0.00433f
C39982 VPWR.t5241 VGND 0.00433f
C39983 VPWR.t1782 VGND 0.00433f
C39984 VPWR.t5045 VGND 0.00433f
C39985 VPWR.t4308 VGND 0.00433f
C39986 VPWR.t3788 VGND 0.00433f
C39987 VPWR.t4770 VGND 0.00433f
C39988 VPWR.t3609 VGND 0.00433f
C39989 VPWR.t591 VGND 0.00433f
C39990 VPWR.t3231 VGND 0.0298f
C39991 VPWR.t2144 VGND 0.04521f
C39992 VPWR.t5821 VGND 0.0173f
C39993 VPWR.t4018 VGND 0.04521f
C39994 VPWR.t1071 VGND 0.03248f
C39995 VPWR.t5603 VGND 0.05001f
C39996 VPWR.t6038 VGND 0.02791f
C39997 VPWR.t5601 VGND 0.0173f
C39998 VPWR.t1781 VGND 0.06731f
C39999 VPWR.t4307 VGND 0.10001f
C40000 VPWR.t3787 VGND 0.10001f
C40001 VPWR.t590 VGND 0.08271f
C40002 VPWR.t6179 VGND 0.04122f
C40003 VPWR.t6180 VGND 0.00433f
C40004 VPWR.t2219 VGND 0.00433f
C40005 VPWR.t4970 VGND 0.00433f
C40006 VPWR.t4540 VGND 0.00433f
C40007 VPWR.t1134 VGND 0.00433f
C40008 VPWR.t2010 VGND 0.00433f
C40009 VPWR.t757 VGND 0.00433f
C40010 VPWR.t6001 VGND 0.00433f
C40011 VPWR.t6194 VGND 0.00433f
C40012 VPWR.t5700 VGND 0.00433f
C40013 VPWR.t2430 VGND 0.00433f
C40014 VPWR.t2320 VGND 0.00433f
C40015 VPWR.t4368 VGND 0.00433f
C40016 VPWR.t2518 VGND 0.00433f
C40017 VPWR.t4848 VGND 0.00433f
C40018 VPWR.t4311 VGND 0.00433f
C40019 VPWR.t724 VGND 0.00433f
C40020 VPWR.t2218 VGND 0.0298f
C40021 VPWR.t4969 VGND 0.05001f
C40022 VPWR.t4539 VGND 0.05001f
C40023 VPWR.t1133 VGND 0.05001f
C40024 VPWR.t2009 VGND 0.05001f
C40025 VPWR.t756 VGND 0.05001f
C40026 VPWR.t6000 VGND 0.05001f
C40027 VPWR.t6193 VGND 0.05001f
C40028 VPWR.t5699 VGND 0.05001f
C40029 VPWR.t2429 VGND 0.05001f
C40030 VPWR.t2319 VGND 0.05001f
C40031 VPWR.t4367 VGND 0.05001f
C40032 VPWR.t2517 VGND 0.05001f
C40033 VPWR.t4847 VGND 0.04521f
C40034 VPWR.t4310 VGND 0.0173f
C40035 VPWR.t723 VGND 0.05001f
C40036 VPWR.t5768 VGND 0.06143f
C40037 VPWR.t5769 VGND 0.00433f
C40038 VPWR.t3185 VGND 0.00433f
C40039 VPWR.t5679 VGND 0.00433f
C40040 VPWR.t2757 VGND 0.00433f
C40041 VPWR.t3516 VGND 0.00433f
C40042 VPWR.t4358 VGND 0.00433f
C40043 VPWR.t1774 VGND 0.00433f
C40044 VPWR.t1277 VGND 0.00433f
C40045 VPWR.t1172 VGND 0.00433f
C40046 VPWR.t1448 VGND 0.00433f
C40047 VPWR.t605 VGND 0.00433f
C40048 VPWR.t4907 VGND 0.00433f
C40049 VPWR.t2143 VGND 0.00433f
C40050 VPWR.t1880 VGND 0.00433f
C40051 VPWR.t4196 VGND 0.00433f
C40052 VPWR.t5163 VGND 0.00433f
C40053 VPWR.t3184 VGND 0.0298f
C40054 VPWR.t5678 VGND 0.05001f
C40055 VPWR.t2756 VGND 0.05001f
C40056 VPWR.t3515 VGND 0.05001f
C40057 VPWR.t4357 VGND 0.05001f
C40058 VPWR.t1773 VGND 0.05001f
C40059 VPWR.t1276 VGND 0.05001f
C40060 VPWR.t1171 VGND 0.05001f
C40061 VPWR.t1447 VGND 0.05001f
C40062 VPWR.t604 VGND 0.05001f
C40063 VPWR.t4906 VGND 0.05001f
C40064 VPWR.t2142 VGND 0.05001f
C40065 VPWR.t1879 VGND 0.05001f
C40066 VPWR.t4195 VGND 0.04521f
C40067 VPWR.t5162 VGND 0.025f
C40068 VPWR.n349 VGND 0.00665f
C40069 VPWR.n350 VGND 0.00834f
C40070 VPWR.n351 VGND 0.01085f
C40071 VPWR.n352 VGND 0.01085f
C40072 VPWR.n353 VGND 0.01085f
C40073 VPWR.n354 VGND 0.01085f
C40074 VPWR.n355 VGND 0.01085f
C40075 VPWR.n356 VGND 0.00985f
C40076 VPWR.n357 VGND 0.01013f
C40077 VPWR.n358 VGND 0.01073f
C40078 VPWR.n359 VGND 0.13412f
C40079 VPWR.t1058 VGND 0.00433f
C40080 VPWR.n360 VGND 0.01073f
C40081 VPWR.t3463 VGND 0.00427f
C40082 VPWR.t4403 VGND 0.0202f
C40083 VPWR.t4404 VGND 0.00433f
C40084 VPWR.t1182 VGND 0.00433f
C40085 VPWR.t1181 VGND 0.025f
C40086 VPWR.n361 VGND 0.00754f
C40087 VPWR.n362 VGND 0.00738f
C40088 VPWR.t4824 VGND 0.00433f
C40089 VPWR.t3802 VGND 0.00433f
C40090 VPWR.t1373 VGND 0.00433f
C40091 VPWR.t4809 VGND 0.00433f
C40092 VPWR.t5008 VGND 0.00433f
C40093 VPWR.t4579 VGND 0.00433f
C40094 VPWR.n363 VGND 0.0085f
C40095 VPWR.n364 VGND 0.00738f
C40096 VPWR.n365 VGND 0.00974f
C40097 VPWR.n366 VGND 0.0085f
C40098 VPWR.n367 VGND 0.00896f
C40099 VPWR.n368 VGND 0.00754f
C40100 VPWR.n369 VGND 0.01189f
C40101 VPWR.n370 VGND 0.02102f
C40102 VPWR.t4823 VGND 0.03271f
C40103 VPWR.t3801 VGND 0.04231f
C40104 VPWR.t1372 VGND 0.03271f
C40105 VPWR.t4808 VGND 0.05001f
C40106 VPWR.t5007 VGND 0.05001f
C40107 VPWR.t4578 VGND 0.04231f
C40108 VPWR.t1057 VGND 0.0154f
C40109 VPWR.t3462 VGND 0.0202f
C40110 VPWR.n371 VGND 0.03162f
C40111 VPWR.t3461 VGND 0.00473f
C40112 VPWR.t7126 VGND 0.00433f
C40113 VPWR.t309 VGND 0.00427f
C40114 VPWR.t3447 VGND 0.00433f
C40115 VPWR.t311 VGND 0.00473f
C40116 VPWR.t3121 VGND 0.00427f
C40117 VPWR.t2875 VGND 0.00433f
C40118 VPWR.t3119 VGND 0.00473f
C40119 VPWR.t471 VGND 0.00433f
C40120 VPWR.t3460 VGND 0.0173f
C40121 VPWR.t7125 VGND 0.01172f
C40122 VPWR.t308 VGND 0.03483f
C40123 VPWR.t310 VGND 0.04309f
C40124 VPWR.t3446 VGND 0.03248f
C40125 VPWR.t3120 VGND 0.0298f
C40126 VPWR.t2874 VGND 0.02791f
C40127 VPWR.t3118 VGND 0.05001f
C40128 VPWR.t470 VGND 0.0737f
C40129 VPWR.t1576 VGND 0.00433f
C40130 VPWR.t2322 VGND 0.00433f
C40131 VPWR.t1064 VGND 0.00433f
C40132 VPWR.t1768 VGND 0.00427f
C40133 VPWR.t4891 VGND 0.00433f
C40134 VPWR.t1770 VGND 0.00473f
C40135 VPWR.t5667 VGND 0.00433f
C40136 VPWR.t5316 VGND 0.00433f
C40137 VPWR.t1720 VGND 0.00433f
C40138 VPWR.t3621 VGND 0.00433f
C40139 VPWR.t7076 VGND 0.00433f
C40140 VPWR.t5349 VGND 0.00433f
C40141 VPWR.t5075 VGND 0.00473f
C40142 VPWR.t3155 VGND 0.00473f
C40143 VPWR.t5073 VGND 0.00427f
C40144 VPWR.t3153 VGND 0.00427f
C40145 VPWR.t5785 VGND 0.00427f
C40146 VPWR.t1575 VGND 0.03271f
C40147 VPWR.t2321 VGND 0.0298f
C40148 VPWR.t1063 VGND 0.01172f
C40149 VPWR.t1767 VGND 0.03483f
C40150 VPWR.t1769 VGND 0.04309f
C40151 VPWR.t4890 VGND 0.04498f
C40152 VPWR.t5666 VGND 0.03271f
C40153 VPWR.t5315 VGND 0.0298f
C40154 VPWR.t1719 VGND 0.03271f
C40155 VPWR.t3620 VGND 0.05001f
C40156 VPWR.t7075 VGND 0.05001f
C40157 VPWR.t5348 VGND 0.0173f
C40158 VPWR.t5074 VGND 0.03538f
C40159 VPWR.t3154 VGND 0.02791f
C40160 VPWR.t5072 VGND 0.02712f
C40161 VPWR.t3152 VGND 0.0125f
C40162 VPWR.t5784 VGND 0.0173f
C40163 VPWR.n372 VGND 0.03162f
C40164 VPWR.t5828 VGND 0.00473f
C40165 VPWR.t5783 VGND 0.00473f
C40166 VPWR.t4843 VGND 0.00473f
C40167 VPWR.t5826 VGND 0.00427f
C40168 VPWR.t2503 VGND 0.00427f
C40169 VPWR.t4841 VGND 0.00427f
C40170 VPWR.t1489 VGND 0.00427f
C40171 VPWR.t2501 VGND 0.00473f
C40172 VPWR.t1965 VGND 0.00433f
C40173 VPWR.t1487 VGND 0.00473f
C40174 VPWR.t2512 VGND 0.00433f
C40175 VPWR.t5782 VGND 0.04018f
C40176 VPWR.t5827 VGND 0.04577f
C40177 VPWR.t5825 VGND 0.03751f
C40178 VPWR.t4842 VGND 0.01172f
C40179 VPWR.t4840 VGND 0.01172f
C40180 VPWR.t2502 VGND 0.01172f
C40181 VPWR.t2500 VGND 0.01172f
C40182 VPWR.t1488 VGND 0.03751f
C40183 VPWR.t1486 VGND 0.04309f
C40184 VPWR.t1964 VGND 0.03248f
C40185 VPWR.t2511 VGND 0.0202f
C40186 VPWR.n373 VGND 0.02102f
C40187 VPWR.t2864 VGND 0.00473f
C40188 VPWR.t5115 VGND 0.00473f
C40189 VPWR.t2862 VGND 0.00427f
C40190 VPWR.t2860 VGND 0.00427f
C40191 VPWR.t5113 VGND 0.00427f
C40192 VPWR.t5493 VGND 0.00427f
C40193 VPWR.t2858 VGND 0.00473f
C40194 VPWR.t5491 VGND 0.00473f
C40195 VPWR.t2863 VGND 0.03538f
C40196 VPWR.t5114 VGND 0.02791f
C40197 VPWR.t2861 VGND 0.01462f
C40198 VPWR.t5112 VGND 0.0154f
C40199 VPWR.t2859 VGND 0.0154f
C40200 VPWR.t5492 VGND 0.01462f
C40201 VPWR.t2857 VGND 0.02791f
C40202 VPWR.t5490 VGND 0.04018f
C40203 VPWR.n374 VGND 0.0391f
C40204 VPWR.t3421 VGND 0.00427f
C40205 VPWR.t3069 VGND 0.00427f
C40206 VPWR.t3420 VGND 0.00473f
C40207 VPWR.t3067 VGND 0.00473f
C40208 VPWR.t5236 VGND 0.00433f
C40209 VPWR.t5583 VGND 0.00433f
C40210 VPWR.t2815 VGND 0.00433f
C40211 VPWR.t3777 VGND 0.00433f
C40212 VPWR.t3549 VGND 0.00433f
C40213 VPWR.t3404 VGND 0.00433f
C40214 VPWR.t2454 VGND 0.00433f
C40215 VPWR.t6763 VGND 0.00116f
C40216 VPWR.t6416 VGND 0.00116f
C40217 VPWR.n375 VGND 0.00236f
C40218 VPWR.t4323 VGND 0.00433f
C40219 VPWR.t438 VGND 0.00255f
C40220 VPWR.t4329 VGND 0.00394f
C40221 VPWR.t4461 VGND 0.00394f
C40222 VPWR.n376 VGND 0.00115f
C40223 VPWR.t4328 VGND 0.01727f
C40224 VPWR.t3068 VGND 0.03963f
C40225 VPWR.t3066 VGND 0.06039f
C40226 VPWR.t5235 VGND 0.03271f
C40227 VPWR.t5582 VGND 0.0173f
C40228 VPWR.t2814 VGND 0.04521f
C40229 VPWR.t3776 VGND 0.05001f
C40230 VPWR.t3548 VGND 0.05001f
C40231 VPWR.t3403 VGND 0.0173f
C40232 VPWR.t6762 VGND 0.0298f
C40233 VPWR.t2453 VGND 0.02277f
C40234 VPWR.t6415 VGND 0.0173f
C40235 VPWR.t4322 VGND 0.02244f
C40236 VPWR.t437 VGND 0.02668f
C40237 VPWR.t5977 VGND 0.01772f
C40238 VPWR.n377 VGND 0.04365f
C40239 VPWR.t6414 VGND 0.01886f
C40240 VPWR.t4460 VGND 0.01652f
C40241 VPWR.t2739 VGND 0.01183f
C40242 VPWR.t942 VGND 0.0202f
C40243 VPWR.n378 VGND 0.03709f
C40244 VPWR.t2738 VGND 0.00107f
C40245 VPWR.n379 VGND 0.00292f
C40246 VPWR.t469 VGND 0.00219f
C40247 VPWR.t301 VGND 0.00185f
C40248 VPWR.n380 VGND 0.00433f
C40249 VPWR.t4564 VGND 0.00427f
C40250 VPWR.t2254 VGND 0.00433f
C40251 VPWR.t4803 VGND 0.00433f
C40252 VPWR.t4662 VGND 0.00433f
C40253 VPWR.t6417 VGND 0.0413f
C40254 VPWR.t4463 VGND 0.03181f
C40255 VPWR.t439 VGND 0.02277f
C40256 VPWR.t302 VGND 0.01741f
C40257 VPWR.t4565 VGND 0.02277f
C40258 VPWR.t468 VGND 0.02768f
C40259 VPWR.t2737 VGND 0.03125f
C40260 VPWR.t300 VGND 0.03259f
C40261 VPWR.t4462 VGND 0.02902f
C40262 VPWR.t4563 VGND 0.01395f
C40263 VPWR.t2253 VGND 0.025f
C40264 VPWR.t4802 VGND 0.0298f
C40265 VPWR.t4661 VGND 0.03538f
C40266 VPWR.n381 VGND 0.01912f
C40267 VPWR.t5002 VGND 0.00203f
C40268 VPWR.n382 VGND 0.00162f
C40269 VPWR.t3611 VGND 0.00219f
C40270 VPWR.t4799 VGND 0.00185f
C40271 VPWR.n383 VGND 0.00433f
C40272 VPWR.t4133 VGND 0.00149f
C40273 VPWR.t7100 VGND 0.00281f
C40274 VPWR.n384 VGND 0.00388f
C40275 VPWR.t5001 VGND 0.0336f
C40276 VPWR.t131 VGND 0.02277f
C40277 VPWR.t4800 VGND 0.02277f
C40278 VPWR.t4795 VGND 0.02277f
C40279 VPWR.t5153 VGND 0.02277f
C40280 VPWR.t3610 VGND 0.02277f
C40281 VPWR.t4132 VGND 0.03125f
C40282 VPWR.t4798 VGND 0.05179f
C40283 VPWR.t136 VGND 0.03192f
C40284 VPWR.n385 VGND 0.01767f
C40285 VPWR.t1908 VGND 0.00427f
C40286 VPWR.t1922 VGND 0.00427f
C40287 VPWR.t3082 VGND 0.00107f
C40288 VPWR.n386 VGND 0.00292f
C40289 VPWR.t2463 VGND 0.00107f
C40290 VPWR.n387 VGND 0.00292f
C40291 VPWR.n388 VGND 0.00115f
C40292 VPWR.n389 VGND 0.00115f
C40293 VPWR.t2078 VGND 0.00255f
C40294 VPWR.t2599 VGND 0.00255f
C40295 VPWR.t200 VGND 0.00116f
C40296 VPWR.t6668 VGND 0.00116f
C40297 VPWR.n390 VGND 0.00236f
C40298 VPWR.t7033 VGND 0.00116f
C40299 VPWR.t6642 VGND 0.00116f
C40300 VPWR.n391 VGND 0.00236f
C40301 VPWR.t1113 VGND 0.01526f
C40302 VPWR.t2077 VGND 0.01925f
C40303 VPWR.t1907 VGND 0.03561f
C40304 VPWR.t1921 VGND 0.03885f
C40305 VPWR.t3081 VGND 0.03885f
C40306 VPWR.t2462 VGND 0.02768f
C40307 VPWR.t1905 VGND 0.02009f
C40308 VPWR.t2076 VGND 0.025f
C40309 VPWR.t1923 VGND 0.025f
C40310 VPWR.t2597 VGND 0.02422f
C40311 VPWR.t197 VGND 0.03181f
C40312 VPWR.t7034 VGND 0.03338f
C40313 VPWR.t1046 VGND 0.03248f
C40314 VPWR.t5552 VGND 0.025f
C40315 VPWR.t1918 VGND 0.01652f
C40316 VPWR.t198 VGND 0.02401f
C40317 VPWR.t464 VGND 0.02462f
C40318 VPWR.t7031 VGND 0.02406f
C40319 VPWR.n392 VGND 0.01946f
C40320 VPWR.n394 VGND 0.02426f
C40321 VPWR.t2598 VGND 0.03918f
C40322 VPWR.t199 VGND 0.04599f
C40323 VPWR.t6667 VGND 0.025f
C40324 VPWR.t7032 VGND 0.01395f
C40325 VPWR.t6641 VGND 0.0125f
C40326 VPWR.t2949 VGND 0.02063f
C40327 VPWR.t6949 VGND 0.02428f
C40328 VPWR.t6819 VGND 0.02428f
C40329 VPWR.t6611 VGND 0.02211f
C40330 VPWR.t3398 VGND 0.01615f
C40331 VPWR.t6606 VGND 0.03024f
C40332 VPWR.t6954 VGND 0.03122f
C40333 VPWR.t6804 VGND 0.02791f
C40334 VPWR.t2951 VGND 0.05066f
C40335 VPWR.t4699 VGND 0.05001f
C40336 VPWR.t4684 VGND 0.03672f
C40337 VPWR.t6390 VGND 0.0125f
C40338 VPWR.t3911 VGND 0.02277f
C40339 VPWR.t6829 VGND 0.02277f
C40340 VPWR.t6286 VGND 0.01261f
C40341 VPWR.t3401 VGND 0.0154f
C40342 VPWR.n395 VGND 0.04122f
C40343 VPWR.t3402 VGND 0.00425f
C40344 VPWR.t6287 VGND 0.00394f
C40345 VPWR.t3912 VGND 0.00394f
C40346 VPWR.t4685 VGND 0.00399f
C40347 VPWR.t6394 VGND 0.00516f
C40348 VPWR.t4700 VGND 0.00145f
C40349 VPWR.t2952 VGND 0.00224f
C40350 VPWR.n396 VGND 0.00444f
C40351 VPWR.t6708 VGND 0.00132f
C40352 VPWR.t6805 VGND 0.00132f
C40353 VPWR.n397 VGND 0.00266f
C40354 VPWR.t3399 VGND 0.00394f
C40355 VPWR.n398 VGND 0.00919f
C40356 VPWR.n399 VGND 0.0088f
C40357 VPWR.n400 VGND 0.00949f
C40358 VPWR.n401 VGND 0.01573f
C40359 VPWR.n402 VGND 0.00941f
C40360 VPWR.n403 VGND 0.00899f
C40361 VPWR.n404 VGND 0.00611f
C40362 VPWR.n405 VGND 0.0099f
C40363 VPWR.n406 VGND 0.00586f
C40364 VPWR.n407 VGND 0.00518f
C40365 VPWR.n408 VGND 0.0092f
C40366 VPWR.n409 VGND 0.01677f
C40367 VPWR.n410 VGND 0.01674f
C40368 VPWR.n411 VGND 0.01848f
C40369 VPWR.n412 VGND 0.01758f
C40370 VPWR.n413 VGND 0.00766f
C40371 VPWR.n414 VGND 0.00901f
C40372 VPWR.n415 VGND 0.01065f
C40373 VPWR.n416 VGND 0.01266f
C40374 VPWR.n417 VGND 0.00833f
C40375 VPWR.n418 VGND 0.0053f
C40376 VPWR.n419 VGND 0.00898f
C40377 VPWR.n420 VGND 0.00622f
C40378 VPWR.n421 VGND 0.01034f
C40379 VPWR.n422 VGND 0.00583f
C40380 VPWR.n423 VGND 0.00594f
C40381 VPWR.n424 VGND 0.00725f
C40382 VPWR.n425 VGND 0.00665f
C40383 VPWR.n426 VGND 0.01343f
C40384 VPWR.n427 VGND 0.00822f
C40385 VPWR.n428 VGND 0.00375f
C40386 VPWR.n429 VGND 0.02119f
C40387 VPWR.n430 VGND 0.006f
C40388 VPWR.n431 VGND 0.00801f
C40389 VPWR.n432 VGND 0.01074f
C40390 VPWR.n433 VGND 0.00641f
C40391 VPWR.n434 VGND 0.00994f
C40392 VPWR.n435 VGND 0.00784f
C40393 VPWR.n436 VGND 0.01234f
C40394 VPWR.n437 VGND 0.01197f
C40395 VPWR.n438 VGND 0.00564f
C40396 VPWR.n439 VGND 0.00974f
C40397 VPWR.n440 VGND 0.01023f
C40398 VPWR.n441 VGND 0.00627f
C40399 VPWR.n442 VGND 0.00588f
C40400 VPWR.n443 VGND 0.01101f
C40401 VPWR.n444 VGND 0.01415f
C40402 VPWR.n445 VGND 0.01189f
C40403 VPWR.n446 VGND 0.0059f
C40404 VPWR.n447 VGND 0.00593f
C40405 VPWR.n448 VGND 0.00646f
C40406 VPWR.n449 VGND 0.00708f
C40407 VPWR.n450 VGND 0.00708f
C40408 VPWR.n451 VGND 0.00646f
C40409 VPWR.n452 VGND 0.00593f
C40410 VPWR.n453 VGND 0.00577f
C40411 VPWR.n454 VGND 0.01266f
C40412 VPWR.n455 VGND 0.0058f
C40413 VPWR.n456 VGND 0.13412f
C40414 VPWR.t5608 VGND 0.00427f
C40415 VPWR.n457 VGND 0.00878f
C40416 VPWR.t2604 VGND 0.00473f
C40417 VPWR.t1711 VGND 0.00473f
C40418 VPWR.t2605 VGND 0.00427f
C40419 VPWR.t1709 VGND 0.00427f
C40420 VPWR.t2601 VGND 0.00427f
C40421 VPWR.t1727 VGND 0.0173f
C40422 VPWR.t1728 VGND 0.00427f
C40423 VPWR.t1732 VGND 0.00427f
C40424 VPWR.t2868 VGND 0.00473f
C40425 VPWR.t1730 VGND 0.00473f
C40426 VPWR.t2870 VGND 0.00427f
C40427 VPWR.t4497 VGND 0.00473f
C40428 VPWR.t5327 VGND 0.00433f
C40429 VPWR.t4499 VGND 0.00427f
C40430 VPWR.t505 VGND 0.00473f
C40431 VPWR.t5188 VGND 0.00427f
C40432 VPWR.t507 VGND 0.00427f
C40433 VPWR.t5190 VGND 0.00473f
C40434 VPWR.t6165 VGND 0.00473f
C40435 VPWR.t509 VGND 0.00427f
C40436 VPWR.t6163 VGND 0.00427f
C40437 VPWR.t511 VGND 0.00473f
C40438 VPWR.t4143 VGND 0.00473f
C40439 VPWR.t4607 VGND 0.00427f
C40440 VPWR.t4145 VGND 0.00427f
C40441 VPWR.t4609 VGND 0.00473f
C40442 VPWR.t3113 VGND 0.00473f
C40443 VPWR.t1731 VGND 0.03248f
C40444 VPWR.t2867 VGND 0.02791f
C40445 VPWR.t1729 VGND 0.02791f
C40446 VPWR.t2869 VGND 0.03248f
C40447 VPWR.t5326 VGND 0.03248f
C40448 VPWR.t4496 VGND 0.03271f
C40449 VPWR.t4498 VGND 0.0221f
C40450 VPWR.t504 VGND 0.01172f
C40451 VPWR.t5187 VGND 0.02791f
C40452 VPWR.t506 VGND 0.02791f
C40453 VPWR.t5189 VGND 0.01172f
C40454 VPWR.t6164 VGND 0.01172f
C40455 VPWR.t508 VGND 0.02791f
C40456 VPWR.t6162 VGND 0.02791f
C40457 VPWR.t510 VGND 0.01172f
C40458 VPWR.t4142 VGND 0.01172f
C40459 VPWR.t4606 VGND 0.02791f
C40460 VPWR.t4144 VGND 0.02791f
C40461 VPWR.t4608 VGND 0.01172f
C40462 VPWR.t3112 VGND 0.0298f
C40463 VPWR.n458 VGND 0.03162f
C40464 VPWR.t3115 VGND 0.00427f
C40465 VPWR.t751 VGND 0.00427f
C40466 VPWR.t1638 VGND 0.00473f
C40467 VPWR.t753 VGND 0.00473f
C40468 VPWR.t1492 VGND 0.00427f
C40469 VPWR.t1640 VGND 0.00427f
C40470 VPWR.t2831 VGND 0.00473f
C40471 VPWR.t1494 VGND 0.00473f
C40472 VPWR.t6314 VGND 0.00473f
C40473 VPWR.t2829 VGND 0.00427f
C40474 VPWR.t2827 VGND 0.00427f
C40475 VPWR.t6316 VGND 0.00427f
C40476 VPWR.t2825 VGND 0.00473f
C40477 VPWR.t5403 VGND 0.00433f
C40478 VPWR.t5445 VGND 0.00433f
C40479 VPWR.t3114 VGND 0.0173f
C40480 VPWR.t750 VGND 0.0125f
C40481 VPWR.t752 VGND 0.03248f
C40482 VPWR.t1637 VGND 0.03326f
C40483 VPWR.t1639 VGND 0.03003f
C40484 VPWR.t1491 VGND 0.03003f
C40485 VPWR.t1493 VGND 0.03326f
C40486 VPWR.t2830 VGND 0.03326f
C40487 VPWR.t2828 VGND 0.03963f
C40488 VPWR.t6313 VGND 0.0154f
C40489 VPWR.t2826 VGND 0.02288f
C40490 VPWR.t6315 VGND 0.02288f
C40491 VPWR.t2824 VGND 0.0154f
C40492 VPWR.t5402 VGND 0.025f
C40493 VPWR.t5444 VGND 0.025f
C40494 VPWR.n459 VGND 0.00665f
C40495 VPWR.n460 VGND 0.00738f
C40496 VPWR.n461 VGND 0.00705f
C40497 VPWR.n462 VGND 0.00655f
C40498 VPWR.n463 VGND 0.00646f
C40499 VPWR.n464 VGND 0.00593f
C40500 VPWR.n465 VGND 0.00655f
C40501 VPWR.n466 VGND 0.0054f
C40502 VPWR.n467 VGND 0.0054f
C40503 VPWR.n468 VGND 0.0077f
C40504 VPWR.n469 VGND 0.0077f
C40505 VPWR.n470 VGND 0.00345f
C40506 VPWR.n471 VGND 0.00724f
C40507 VPWR.n472 VGND 0.00494f
C40508 VPWR.n473 VGND 0.00557f
C40509 VPWR.n474 VGND 0.00642f
C40510 VPWR.n475 VGND 0.01077f
C40511 VPWR.n476 VGND 0.0063f
C40512 VPWR.n477 VGND 0.00584f
C40513 VPWR.n478 VGND 0.00655f
C40514 VPWR.n479 VGND 0.00655f
C40515 VPWR.n480 VGND 0.00584f
C40516 VPWR.n481 VGND 0.00584f
C40517 VPWR.n482 VGND 0.00655f
C40518 VPWR.n483 VGND 0.00655f
C40519 VPWR.n484 VGND 0.00584f
C40520 VPWR.n485 VGND 0.00584f
C40521 VPWR.n486 VGND 0.00655f
C40522 VPWR.n487 VGND 0.00655f
C40523 VPWR.n488 VGND 0.00469f
C40524 VPWR.n489 VGND 0.00776f
C40525 VPWR.n490 VGND 0.00685f
C40526 VPWR.n491 VGND 0.00481f
C40527 VPWR.n492 VGND 0.00934f
C40528 VPWR.n493 VGND 0.00655f
C40529 VPWR.n494 VGND 0.00655f
C40530 VPWR.n495 VGND 0.00698f
C40531 VPWR.n496 VGND 0.00642f
C40532 VPWR.t1726 VGND 0.00473f
C40533 VPWR.t4724 VGND 0.00473f
C40534 VPWR.t736 VGND 0.00473f
C40535 VPWR.t4722 VGND 0.00427f
C40536 VPWR.t5340 VGND 0.00427f
C40537 VPWR.t734 VGND 0.00427f
C40538 VPWR.t3989 VGND 0.00427f
C40539 VPWR.t5338 VGND 0.00473f
C40540 VPWR.t3991 VGND 0.00473f
C40541 VPWR.t5088 VGND 0.00433f
C40542 VPWR.t3337 VGND 0.00427f
C40543 VPWR.t3339 VGND 0.00473f
C40544 VPWR.t5610 VGND 0.00473f
C40545 VPWR.t4096 VGND 0.00433f
C40546 VPWR.n497 VGND 0.00685f
C40547 VPWR.n498 VGND 0.00584f
C40548 VPWR.n499 VGND 0.00646f
C40549 VPWR.n500 VGND 0.01257f
C40550 VPWR.n501 VGND 0.00608f
C40551 VPWR.n502 VGND 0.00593f
C40552 VPWR.n503 VGND 0.00646f
C40553 VPWR.n504 VGND 0.00708f
C40554 VPWR.n505 VGND 0.00708f
C40555 VPWR.n506 VGND 0.00646f
C40556 VPWR.n507 VGND 0.00593f
C40557 VPWR.n508 VGND 0.00577f
C40558 VPWR.n509 VGND 0.0052f
C40559 VPWR.n510 VGND 0.01077f
C40560 VPWR.n511 VGND 0.0266f
C40561 VPWR.t1725 VGND 0.025f
C40562 VPWR.t4723 VGND 0.03538f
C40563 VPWR.t735 VGND 0.02791f
C40564 VPWR.t4721 VGND 0.01462f
C40565 VPWR.t733 VGND 0.0154f
C40566 VPWR.t5339 VGND 0.0154f
C40567 VPWR.t3988 VGND 0.01462f
C40568 VPWR.t5337 VGND 0.02791f
C40569 VPWR.t3990 VGND 0.04498f
C40570 VPWR.t3336 VGND 0.0173f
C40571 VPWR.t5087 VGND 0.02288f
C40572 VPWR.t3338 VGND 0.03538f
C40573 VPWR.t5609 VGND 0.05269f
C40574 VPWR.t4095 VGND 0.02791f
C40575 VPWR.t5607 VGND 0.0173f
C40576 VPWR.t1710 VGND 0.06329f
C40577 VPWR.t1708 VGND 0.03963f
C40578 VPWR.n512 VGND 0.01544f
C40579 VPWR.t2603 VGND 0.00473f
C40580 VPWR.t3425 VGND 0.00473f
C40581 VPWR.t6745 VGND 0.00116f
C40582 VPWR.t6597 VGND 0.00116f
C40583 VPWR.n513 VGND 0.00236f
C40584 VPWR.t3423 VGND 0.00427f
C40585 VPWR.t5177 VGND 0.00427f
C40586 VPWR.t3943 VGND 0.00255f
C40587 VPWR.t5175 VGND 0.00473f
C40588 VPWR.t6249 VGND 0.00433f
C40589 VPWR.n514 VGND 0.00115f
C40590 VPWR.t5165 VGND 0.00433f
C40591 VPWR.t1945 VGND 0.00433f
C40592 VPWR.t878 VGND 0.00107f
C40593 VPWR.n515 VGND 0.00292f
C40594 VPWR.t1850 VGND 0.00433f
C40595 VPWR.t3252 VGND 0.00427f
C40596 VPWR.t1748 VGND 0.00433f
C40597 VPWR.t3784 VGND 0.01653f
C40598 VPWR.t5174 VGND 0.02333f
C40599 VPWR.t2600 VGND 0.0173f
C40600 VPWR.t2602 VGND 0.025f
C40601 VPWR.t3424 VGND 0.01395f
C40602 VPWR.t6744 VGND 0.02791f
C40603 VPWR.t3422 VGND 0.02277f
C40604 VPWR.t6596 VGND 0.01172f
C40605 VPWR.t5176 VGND 0.02244f
C40606 VPWR.t3942 VGND 0.02668f
C40607 VPWR.n517 VGND 0.03621f
C40608 VPWR.t6598 VGND 0.01909f
C40609 VPWR.t6157 VGND 0.03014f
C40610 VPWR.t6248 VGND 0.02411f
C40611 VPWR.t1019 VGND 0.0173f
C40612 VPWR.t6595 VGND 0.03271f
C40613 VPWR.t5164 VGND 0.03181f
C40614 VPWR.t3944 VGND 0.04309f
C40615 VPWR.t3253 VGND 0.02433f
C40616 VPWR.t1944 VGND 0.02768f
C40617 VPWR.t877 VGND 0.05001f
C40618 VPWR.t1849 VGND 0.03885f
C40619 VPWR.t3251 VGND 0.05001f
C40620 VPWR.t1747 VGND 0.06143f
C40621 VPWR.t730 VGND 0.00473f
C40622 VPWR.t304 VGND 0.00394f
C40623 VPWR.t3931 VGND 0.00394f
C40624 VPWR.t3933 VGND 0.00498f
C40625 VPWR.t4793 VGND 0.00114f
C40626 VPWR.t5006 VGND 0.00114f
C40627 VPWR.n518 VGND 0.00228f
C40628 VPWR.t4696 VGND 0.00334f
C40629 VPWR.t4325 VGND 0.00114f
C40630 VPWR.t3300 VGND 0.00114f
C40631 VPWR.n519 VGND 0.00228f
C40632 VPWR.t4321 VGND 0.00132f
C40633 VPWR.t3298 VGND 0.00132f
C40634 VPWR.n520 VGND 0.00267f
C40635 VPWR.t3296 VGND 0.00114f
C40636 VPWR.t4327 VGND 0.00114f
C40637 VPWR.n521 VGND 0.00228f
C40638 VPWR.t3055 VGND 0.00433f
C40639 VPWR.t5000 VGND 0.00114f
C40640 VPWR.t4805 VGND 0.00114f
C40641 VPWR.n522 VGND 0.0023f
C40642 VPWR.t196 VGND 0.00473f
C40643 VPWR.t3302 VGND 0.00433f
C40644 VPWR.t185 VGND 0.00431f
C40645 VPWR.t5392 VGND 0.00498f
C40646 VPWR.t729 VGND 0.0154f
C40647 VPWR.t303 VGND 0.02065f
C40648 VPWR.t2004 VGND 0.02277f
C40649 VPWR.t3930 VGND 0.025f
C40650 VPWR.t3960 VGND 0.02791f
C40651 VPWR.t3932 VGND 0.01172f
C40652 VPWR.t4792 VGND 0.01395f
C40653 VPWR.t5005 VGND 0.0154f
C40654 VPWR.t4695 VGND 0.01976f
C40655 VPWR.t4324 VGND 0.02277f
C40656 VPWR.t4320 VGND 0.02277f
C40657 VPWR.t3299 VGND 0.02277f
C40658 VPWR.t3297 VGND 0.02277f
C40659 VPWR.t3295 VGND 0.02433f
C40660 VPWR.t4326 VGND 0.02623f
C40661 VPWR.t4999 VGND 0.02925f
C40662 VPWR.t3054 VGND 0.02277f
C40663 VPWR.t4804 VGND 0.0173f
C40664 VPWR.t195 VGND 0.05079f
C40665 VPWR.t3301 VGND 0.02277f
C40666 VPWR.t3771 VGND 0.01172f
C40667 VPWR.t6620 VGND 0.025f
C40668 VPWR.t5391 VGND 0.0154f
C40669 VPWR.t184 VGND 0.0202f
C40670 VPWR.n523 VGND 0.02649f
C40671 VPWR.t133 VGND 0.00431f
C40672 VPWR.t5158 VGND 0.00187f
C40673 VPWR.t1168 VGND 0.00139f
C40674 VPWR.n524 VGND 0.00471f
C40675 VPWR.t5161 VGND 0.00425f
C40676 VPWR.t5004 VGND 0.00425f
C40677 VPWR.t6707 VGND 0.00433f
C40678 VPWR.t202 VGND 0.00429f
C40679 VPWR.t5156 VGND 0.00394f
C40680 VPWR.t4136 VGND 0.00394f
C40681 VPWR.t3274 VGND 0.00425f
C40682 VPWR.t5159 VGND 0.0173f
C40683 VPWR.t939 VGND 0.025f
C40684 VPWR.t132 VGND 0.0125f
C40685 VPWR.t4998 VGND 0.02534f
C40686 VPWR.t6715 VGND 0.02277f
C40687 VPWR.t5157 VGND 0.04298f
C40688 VPWR.t1167 VGND 0.04699f
C40689 VPWR.t5160 VGND 0.04431f
C40690 VPWR.t5996 VGND 0.03751f
C40691 VPWR.t5003 VGND 0.02277f
C40692 VPWR.t4134 VGND 0.02467f
C40693 VPWR.t4797 VGND 0.0154f
C40694 VPWR.t4465 VGND 0.01183f
C40695 VPWR.t4464 VGND 0.01172f
C40696 VPWR.t3200 VGND 0.03829f
C40697 VPWR.t6706 VGND 0.025f
C40698 VPWR.t5997 VGND 0.03449f
C40699 VPWR.t6731 VGND 0.02579f
C40700 VPWR.t5155 VGND 0.02579f
C40701 VPWR.t4135 VGND 0.02467f
C40702 VPWR.t3273 VGND 0.01183f
C40703 VPWR.n525 VGND 0.03162f
C40704 VPWR.t6717 VGND 0.00425f
C40705 VPWR.t3019 VGND 0.00379f
C40706 VPWR.t6798 VGND 0.00152f
C40707 VPWR.t6811 VGND 0.00152f
C40708 VPWR.n526 VGND 0.00306f
C40709 VPWR.t6710 VGND 0.0039f
C40710 VPWR.t3017 VGND 0.00147f
C40711 VPWR.t3023 VGND 0.00147f
C40712 VPWR.n527 VGND 0.00295f
C40713 VPWR.t6240 VGND 0.00529f
C40714 VPWR.n528 VGND 0.00208f
C40715 VPWR.t3021 VGND 0.00166f
C40716 VPWR.t4993 VGND 0.00183f
C40717 VPWR.n529 VGND 0.0043f
C40718 VPWR.t5439 VGND 0.00123f
C40719 VPWR.n530 VGND 0.00172f
C40720 VPWR.t232 VGND 0.00132f
C40721 VPWR.t230 VGND 0.00132f
C40722 VPWR.n531 VGND 0.00266f
C40723 VPWR.t4989 VGND 0.00132f
C40724 VPWR.t4991 VGND 0.00132f
C40725 VPWR.n532 VGND 0.00266f
C40726 VPWR.t234 VGND 0.00132f
C40727 VPWR.t228 VGND 0.00132f
C40728 VPWR.n533 VGND 0.00266f
C40729 VPWR.n534 VGND 0.00116f
C40730 VPWR.t4987 VGND 0.00332f
C40731 VPWR.t6716 VGND 0.01395f
C40732 VPWR.t3018 VGND 0.02355f
C40733 VPWR.t6797 VGND 0.0281f
C40734 VPWR.t4686 VGND 0.02211f
C40735 VPWR.t6810 VGND 0.02211f
C40736 VPWR.t4701 VGND 0.02211f
C40737 VPWR.t6709 VGND 0.01745f
C40738 VPWR.t3016 VGND 0.02851f
C40739 VPWR.t6239 VGND 0.02211f
C40740 VPWR.t3022 VGND 0.02905f
C40741 VPWR.t4688 VGND 0.03317f
C40742 VPWR.t3830 VGND 0.02211f
C40743 VPWR.t4680 VGND 0.01821f
C40744 VPWR.t3829 VGND 0.02769f
C40745 VPWR.t3020 VGND 0.04944f
C40746 VPWR.t5437 VGND 0.02724f
C40747 VPWR.t4992 VGND 0.01875f
C40748 VPWR.t5438 VGND 0.02277f
C40749 VPWR.t231 VGND 0.0317f
C40750 VPWR.t5047 VGND 0.02277f
C40751 VPWR.t229 VGND 0.01875f
C40752 VPWR.t5046 VGND 0.02277f
C40753 VPWR.t4988 VGND 0.02746f
C40754 VPWR.t4990 VGND 0.04398f
C40755 VPWR.t2504 VGND 0.02277f
C40756 VPWR.t233 VGND 0.01875f
C40757 VPWR.t2505 VGND 0.02277f
C40758 VPWR.t227 VGND 0.025f
C40759 VPWR.t6958 VGND 0.02277f
C40760 VPWR.t4986 VGND 0.0173f
C40761 VPWR.n535 VGND 0.042f
C40762 VPWR.t3400 VGND 0.00433f
C40763 VPWR.t6953 VGND 0.00431f
C40764 VPWR.t4270 VGND 0.00433f
C40765 VPWR.t4850 VGND 0.00433f
C40766 VPWR.t6824 VGND 0.00132f
C40767 VPWR.t6893 VGND 0.00132f
C40768 VPWR.n536 VGND 0.00266f
C40769 VPWR.t4683 VGND 0.00307f
C40770 VPWR.t6586 VGND 0.00516f
C40771 VPWR.t5121 VGND 0.00114f
C40772 VPWR.t6891 VGND 0.00114f
C40773 VPWR.n537 VGND 0.00229f
C40774 VPWR.t5824 VGND 0.00281f
C40775 VPWR.t5814 VGND 0.00149f
C40776 VPWR.n538 VGND 0.00388f
C40777 VPWR.t6419 VGND 0.00307f
C40778 VPWR.n539 VGND 0.00162f
C40779 VPWR.t5147 VGND 0.00181f
C40780 VPWR.t6423 VGND 0.0018f
C40781 VPWR.n540 VGND 0.00494f
C40782 VPWR.t6584 VGND 0.00203f
C40783 VPWR.t3352 VGND 0.00203f
C40784 VPWR.t2377 VGND 0.04309f
C40785 VPWR.t3397 VGND 0.03672f
C40786 VPWR.t6952 VGND 0.0125f
C40787 VPWR.t4269 VGND 0.03829f
C40788 VPWR.t6823 VGND 0.05001f
C40789 VPWR.t4849 VGND 0.02277f
C40790 VPWR.t6892 VGND 0.0173f
C40791 VPWR.t3349 VGND 0.02902f
C40792 VPWR.t4682 VGND 0.02277f
C40793 VPWR.t6585 VGND 0.02099f
C40794 VPWR.t5120 VGND 0.02456f
C40795 VPWR.t6890 VGND 0.02534f
C40796 VPWR.t5823 VGND 0.02277f
C40797 VPWR.t6418 VGND 0.02902f
C40798 VPWR.t5813 VGND 0.01518f
C40799 VPWR.t6377 VGND 0.03561f
C40800 VPWR.t5146 VGND 0.02277f
C40801 VPWR.t960 VGND 0.02634f
C40802 VPWR.t6583 VGND 0.02634f
C40803 VPWR.t6422 VGND 0.01306f
C40804 VPWR.t3351 VGND 0.0125f
C40805 VPWR.t3716 VGND 0.0173f
C40806 VPWR.t4717 VGND 0.03338f
C40807 VPWR.t100 VGND 0.05068f
C40808 VPWR.t1469 VGND 0.03672f
C40809 VPWR.t213 VGND 0.01741f
C40810 VPWR.t6033 VGND 0.025f
C40811 VPWR.t2577 VGND 0.02768f
C40812 VPWR.t2240 VGND 0.02277f
C40813 VPWR.t2331 VGND 0.02154f
C40814 VPWR.t6035 VGND 0.03561f
C40815 VPWR.t3934 VGND 0.04822f
C40816 VPWR.t2578 VGND 0.03706f
C40817 VPWR.t2392 VGND 0.02277f
C40818 VPWR.t6591 VGND 0.02735f
C40819 VPWR.t6379 VGND 0.0154f
C40820 VPWR.t6609 VGND 0.0173f
C40821 VPWR.t2196 VGND 0.02277f
C40822 VPWR.t3346 VGND 0.0298f
C40823 VPWR.t5618 VGND 0.01172f
C40824 VPWR.t4473 VGND 0.03271f
C40825 VPWR.t3348 VGND 0.0173f
C40826 VPWR.t5796 VGND 0.03717f
C40827 VPWR.t6886 VGND 0.0173f
C40828 VPWR.n541 VGND 0.0295f
C40829 VPWR.t6887 VGND 0.00433f
C40830 VPWR.t5797 VGND 0.00433f
C40831 VPWR.t5619 VGND 0.00433f
C40832 VPWR.t4474 VGND 0.00431f
C40833 VPWR.t2197 VGND 0.00433f
C40834 VPWR.n542 VGND 0.00145f
C40835 VPWR.t6592 VGND 0.00203f
C40836 VPWR.t6380 VGND 0.00196f
C40837 VPWR.t2393 VGND 0.00157f
C40838 VPWR.n543 VGND 0.00539f
C40839 VPWR.t2579 VGND 0.0018f
C40840 VPWR.t3935 VGND 0.00181f
C40841 VPWR.n544 VGND 0.00494f
C40842 VPWR.t6036 VGND 0.00427f
C40843 VPWR.t2332 VGND 0.00431f
C40844 VPWR.t2241 VGND 0.00107f
C40845 VPWR.n545 VGND 0.00292f
C40846 VPWR.n546 VGND 0.00778f
C40847 VPWR.n547 VGND 0.00922f
C40848 VPWR.n548 VGND 0.0105f
C40849 VPWR.n549 VGND 0.00962f
C40850 VPWR.n550 VGND 0.00832f
C40851 VPWR.n551 VGND 0.00492f
C40852 VPWR.n552 VGND 0.007f
C40853 VPWR.n553 VGND 0.00645f
C40854 VPWR.n554 VGND 0.00966f
C40855 VPWR.n555 VGND 0.008f
C40856 VPWR.n556 VGND 0.00723f
C40857 VPWR.n557 VGND 0.00756f
C40858 VPWR.n558 VGND 0.01139f
C40859 VPWR.n559 VGND 0.00438f
C40860 VPWR.n560 VGND 0.00623f
C40861 VPWR.n561 VGND 0.00572f
C40862 VPWR.n562 VGND 0.00822f
C40863 VPWR.n563 VGND 0.00882f
C40864 VPWR.n564 VGND 0.00739f
C40865 VPWR.n565 VGND 0.00317f
C40866 VPWR.n566 VGND 0.00901f
C40867 VPWR.n567 VGND 0.00923f
C40868 VPWR.n568 VGND 0.00526f
C40869 VPWR.n569 VGND 0.00627f
C40870 VPWR.n570 VGND 0.00665f
C40871 VPWR.n571 VGND 0.00657f
C40872 VPWR.n572 VGND 0.00829f
C40873 VPWR.n573 VGND 0.01337f
C40874 VPWR.n574 VGND 0.00956f
C40875 VPWR.n575 VGND 0.00466f
C40876 VPWR.n576 VGND 0.00687f
C40877 VPWR.n577 VGND 0.01115f
C40878 VPWR.n578 VGND 0.01081f
C40879 VPWR.n579 VGND 0.00759f
C40880 VPWR.n580 VGND 0.0078f
C40881 VPWR.n581 VGND 0.00883f
C40882 VPWR.n582 VGND 0.015f
C40883 VPWR.n583 VGND 0.00883f
C40884 VPWR.n584 VGND 0.01281f
C40885 VPWR.n585 VGND 0.00795f
C40886 VPWR.n586 VGND 0.00973f
C40887 VPWR.n587 VGND 0.00532f
C40888 VPWR.n588 VGND 0.01089f
C40889 VPWR.n589 VGND 0.00651f
C40890 VPWR.n590 VGND 0.00727f
C40891 VPWR.n591 VGND 0.00727f
C40892 VPWR.n592 VGND 0.00928f
C40893 VPWR.n593 VGND 0.00878f
C40894 VPWR.n594 VGND 0.01044f
C40895 VPWR.n595 VGND 0.01101f
C40896 VPWR.n596 VGND 0.00697f
C40897 VPWR.n597 VGND 0.01062f
C40898 VPWR.n598 VGND 0.01077f
C40899 VPWR.n599 VGND 0.00803f
C40900 VPWR.n600 VGND 0.00777f
C40901 VPWR.n601 VGND 0.13412f
C40902 VPWR.t6803 VGND 0.00152f
C40903 VPWR.t6796 VGND 0.00152f
C40904 VPWR.n602 VGND 0.00306f
C40905 VPWR.n603 VGND 0.00454f
C40906 VPWR.t1263 VGND 0.0039f
C40907 VPWR.t3773 VGND 0.00394f
C40908 VPWR.n604 VGND 0.02872f
C40909 VPWR.t3304 VGND 0.002f
C40910 VPWR.t3306 VGND 0.00165f
C40911 VPWR.n605 VGND 0.00366f
C40912 VPWR.t6712 VGND 0.00226f
C40913 VPWR.t6714 VGND 0.00163f
C40914 VPWR.n606 VGND 0.00392f
C40915 VPWR.t1 VGND 0.00433f
C40916 VPWR.t1327 VGND 0.00159f
C40917 VPWR.t850 VGND 0.00158f
C40918 VPWR.n607 VGND 0.00497f
C40919 VPWR.t258 VGND 0.00296f
C40920 VPWR.t252 VGND 0.0011f
C40921 VPWR.t246 VGND 0.00153f
C40922 VPWR.n608 VGND 0.00265f
C40923 VPWR.t254 VGND 0.0011f
C40924 VPWR.t248 VGND 0.00153f
C40925 VPWR.n609 VGND 0.00265f
C40926 VPWR.t1265 VGND 0.00516f
C40927 VPWR.t268 VGND 0.0011f
C40928 VPWR.t272 VGND 0.00153f
C40929 VPWR.n610 VGND 0.00265f
C40930 VPWR.t6801 VGND 0.00434f
C40931 VPWR.t266 VGND 0.00229f
C40932 VPWR.t6930 VGND 0.00173f
C40933 VPWR.n611 VGND 0.00485f
C40934 VPWR.t3303 VGND 0.03538f
C40935 VPWR.t1473 VGND 0.025f
C40936 VPWR.t3305 VGND 0.02277f
C40937 VPWR.t4237 VGND 0.025f
C40938 VPWR.t5586 VGND 0.02322f
C40939 VPWR.t4236 VGND 0.02277f
C40940 VPWR.t896 VGND 0.025f
C40941 VPWR.t1472 VGND 0.02277f
C40942 VPWR.t4791 VGND 0.02277f
C40943 VPWR.t6711 VGND 0.02322f
C40944 VPWR.t4796 VGND 0.025f
C40945 VPWR.t6713 VGND 0.02277f
C40946 VPWR.t895 VGND 0.01317f
C40947 VPWR.t849 VGND 0.03271f
C40948 VPWR.t0 VGND 0.01976f
C40949 VPWR.t1326 VGND 0.0154f
C40950 VPWR.t257 VGND 0.01886f
C40951 VPWR.t122 VGND 0.025f
C40952 VPWR.t251 VGND 0.025f
C40953 VPWR.t6507 VGND 0.025f
C40954 VPWR.t245 VGND 0.02679f
C40955 VPWR.t19 VGND 0.02288f
C40956 VPWR.t253 VGND 0.0154f
C40957 VPWR.t247 VGND 0.01395f
C40958 VPWR.t1264 VGND 0.025f
C40959 VPWR.t267 VGND 0.04778f
C40960 VPWR.t271 VGND 0.02724f
C40961 VPWR.t6800 VGND 0.025f
C40962 VPWR.t265 VGND 0.04085f
C40963 VPWR.n612 VGND 0.03274f
C40964 VPWR.t6932 VGND 0.00164f
C40965 VPWR.t6928 VGND 0.00227f
C40966 VPWR.n613 VGND 0.00392f
C40967 VPWR.n614 VGND 0.00116f
C40968 VPWR.t6924 VGND 0.00164f
C40969 VPWR.t6916 VGND 0.00227f
C40970 VPWR.n615 VGND 0.00392f
C40971 VPWR.t6912 VGND 0.00164f
C40972 VPWR.t6914 VGND 0.00227f
C40973 VPWR.n616 VGND 0.00392f
C40974 VPWR.t6910 VGND 0.00164f
C40975 VPWR.t6936 VGND 0.00227f
C40976 VPWR.n617 VGND 0.00392f
C40977 VPWR.t4982 VGND 0.00123f
C40978 VPWR.n618 VGND 0.00172f
C40979 VPWR.t6940 VGND 0.00164f
C40980 VPWR.t6934 VGND 0.00227f
C40981 VPWR.n619 VGND 0.00392f
C40982 VPWR.t6938 VGND 0.00164f
C40983 VPWR.t6922 VGND 0.00227f
C40984 VPWR.n620 VGND 0.00392f
C40985 VPWR.t3732 VGND 0.00529f
C40986 VPWR.n621 VGND 0.00208f
C40987 VPWR.t6920 VGND 0.00164f
C40988 VPWR.t6926 VGND 0.00227f
C40989 VPWR.n622 VGND 0.00392f
C40990 VPWR.t5629 VGND 0.00281f
C40991 VPWR.t6963 VGND 0.00149f
C40992 VPWR.n623 VGND 0.00388f
C40993 VPWR.t6918 VGND 0.00425f
C40994 VPWR.t6929 VGND 0.0173f
C40995 VPWR.t6931 VGND 0.025f
C40996 VPWR.t6927 VGND 0.0173f
C40997 VPWR.t2541 VGND 0.025f
C40998 VPWR.t6923 VGND 0.025f
C40999 VPWR.t1788 VGND 0.025f
C41000 VPWR.t6915 VGND 0.01875f
C41001 VPWR.t1787 VGND 0.025f
C41002 VPWR.t6911 VGND 0.04219f
C41003 VPWR.t6913 VGND 0.03148f
C41004 VPWR.t4980 VGND 0.025f
C41005 VPWR.t6909 VGND 0.01875f
C41006 VPWR.t4978 VGND 0.025f
C41007 VPWR.t6935 VGND 0.0317f
C41008 VPWR.t4981 VGND 0.025f
C41009 VPWR.t6939 VGND 0.01875f
C41010 VPWR.t4983 VGND 0.025f
C41011 VPWR.t6933 VGND 0.04867f
C41012 VPWR.t3360 VGND 0.025f
C41013 VPWR.t6937 VGND 0.01875f
C41014 VPWR.t3361 VGND 0.025f
C41015 VPWR.t6921 VGND 0.03192f
C41016 VPWR.t6919 VGND 0.02992f
C41017 VPWR.t3731 VGND 0.025f
C41018 VPWR.t6925 VGND 0.04108f
C41019 VPWR.t5628 VGND 0.025f
C41020 VPWR.t6917 VGND 0.02902f
C41021 VPWR.t6962 VGND 0.03137f
C41022 VPWR.t3915 VGND 0.0202f
C41023 VPWR.n624 VGND 0.02649f
C41024 VPWR.n625 VGND 0.00162f
C41025 VPWR.t6603 VGND 0.00203f
C41026 VPWR.t2649 VGND 0.00431f
C41027 VPWR.t1764 VGND 0.00438f
C41028 VPWR.t1762 VGND 0.00431f
C41029 VPWR.t5255 VGND 0.00394f
C41030 VPWR.t6600 VGND 0.00431f
C41031 VPWR.t1289 VGND 0.00431f
C41032 VPWR.t4820 VGND 0.00132f
C41033 VPWR.t4232 VGND 0.00132f
C41034 VPWR.n626 VGND 0.00267f
C41035 VPWR.t3345 VGND 0.00307f
C41036 VPWR.t6108 VGND 0.00334f
C41037 VPWR.t6605 VGND 0.00114f
C41038 VPWR.t6594 VGND 0.00114f
C41039 VPWR.n627 VGND 0.00229f
C41040 VPWR.t2378 VGND 0.04175f
C41041 VPWR.t6602 VGND 0.02411f
C41042 VPWR.t6825 VGND 0.01306f
C41043 VPWR.t3914 VGND 0.02579f
C41044 VPWR.t6957 VGND 0.03751f
C41045 VPWR.t224 VGND 0.02277f
C41046 VPWR.t2648 VGND 0.02422f
C41047 VPWR.t3913 VGND 0.02579f
C41048 VPWR.t5713 VGND 0.04018f
C41049 VPWR.t1763 VGND 0.02277f
C41050 VPWR.t1761 VGND 0.02154f
C41051 VPWR.t4309 VGND 0.03608f
C41052 VPWR.t2953 VGND 0.04214f
C41053 VPWR.t5116 VGND 0.02052f
C41054 VPWR.t5254 VGND 0.03672f
C41055 VPWR.t972 VGND 0.0154f
C41056 VPWR.t6599 VGND 0.02065f
C41057 VPWR.t1288 VGND 0.02288f
C41058 VPWR.t3350 VGND 0.02724f
C41059 VPWR.t4819 VGND 0.04677f
C41060 VPWR.t4231 VGND 0.02679f
C41061 VPWR.t3344 VGND 0.02277f
C41062 VPWR.t6107 VGND 0.02277f
C41063 VPWR.t6604 VGND 0.01473f
C41064 VPWR.t6593 VGND 0.0125f
C41065 VPWR.n628 VGND 0.02604f
C41066 VPWR.t6884 VGND 0.00307f
C41067 VPWR.t3591 VGND 0.00433f
C41068 VPWR.t5366 VGND 0.00433f
C41069 VPWR.t6588 VGND 0.00431f
C41070 VPWR.t1664 VGND 0.00433f
C41071 VPWR.t1454 VGND 0.00433f
C41072 VPWR.t5192 VGND 0.00433f
C41073 VPWR.t5540 VGND 0.00431f
C41074 VPWR.t5673 VGND 0.00427f
C41075 VPWR.t3224 VGND 0.00181f
C41076 VPWR.t6376 VGND 0.0018f
C41077 VPWR.n629 VGND 0.00494f
C41078 VPWR.t688 VGND 0.00107f
C41079 VPWR.n630 VGND 0.00292f
C41080 VPWR.t6608 VGND 0.00203f
C41081 VPWR.t6374 VGND 0.00431f
C41082 VPWR.n631 VGND 0.00115f
C41083 VPWR.t6883 VGND 0.0173f
C41084 VPWR.t3590 VGND 0.03717f
C41085 VPWR.t6860 VGND 0.04309f
C41086 VPWR.t6587 VGND 0.03304f
C41087 VPWR.t5365 VGND 0.01172f
C41088 VPWR.t1663 VGND 0.04521f
C41089 VPWR.t1453 VGND 0.0173f
C41090 VPWR.t207 VGND 0.04521f
C41091 VPWR.t5191 VGND 0.02422f
C41092 VPWR.t4472 VGND 0.02355f
C41093 VPWR.t5539 VGND 0.03483f
C41094 VPWR.t5672 VGND 0.01395f
C41095 VPWR.t3223 VGND 0.03695f
C41096 VPWR.t687 VGND 0.02902f
C41097 VPWR.t5674 VGND 0.02858f
C41098 VPWR.t6375 VGND 0.01741f
C41099 VPWR.t1913 VGND 0.02277f
C41100 VPWR.t6607 VGND 0.01797f
C41101 VPWR.t156 VGND 0.0154f
C41102 VPWR.t6373 VGND 0.03181f
C41103 VPWR.t527 VGND 0.02612f
C41104 VPWR.t6601 VGND 0.02411f
C41105 VPWR.t3899 VGND 0.0346f
C41106 VPWR.t153 VGND 0.02389f
C41107 VPWR.n632 VGND 0.01198f
C41108 VPWR.t3092 VGND 0.00433f
C41109 VPWR.t1912 VGND 0.00255f
C41110 VPWR.t4668 VGND 0.00433f
C41111 VPWR.t155 VGND 0.00116f
C41112 VPWR.t6660 VGND 0.00116f
C41113 VPWR.n633 VGND 0.00236f
C41114 VPWR.t583 VGND 0.00433f
C41115 VPWR.t1951 VGND 0.00433f
C41116 VPWR.t718 VGND 0.00433f
C41117 VPWR.t2480 VGND 0.00433f
C41118 VPWR.t704 VGND 0.00433f
C41119 VPWR.t5862 VGND 0.00433f
C41120 VPWR.t2948 VGND 0.00433f
C41121 VPWR.t994 VGND 0.00433f
C41122 VPWR.t4955 VGND 0.00433f
C41123 VPWR.t4936 VGND 0.00433f
C41124 VPWR.t4985 VGND 0.00433f
C41125 VPWR.t4341 VGND 0.00433f
C41126 VPWR.t1033 VGND 0.01775f
C41127 VPWR.n634 VGND 0.02471f
C41128 VPWR.t3091 VGND 0.0374f
C41129 VPWR.t1911 VGND 0.0173f
C41130 VPWR.t4667 VGND 0.03829f
C41131 VPWR.t154 VGND 0.02835f
C41132 VPWR.t6659 VGND 0.03672f
C41133 VPWR.t582 VGND 0.0125f
C41134 VPWR.t1950 VGND 0.03271f
C41135 VPWR.t717 VGND 0.0298f
C41136 VPWR.t2479 VGND 0.03271f
C41137 VPWR.t703 VGND 0.05001f
C41138 VPWR.t5861 VGND 0.05001f
C41139 VPWR.t2947 VGND 0.05001f
C41140 VPWR.t993 VGND 0.05001f
C41141 VPWR.t4954 VGND 0.05001f
C41142 VPWR.t4935 VGND 0.05001f
C41143 VPWR.t4984 VGND 0.0298f
C41144 VPWR.t5380 VGND 0.0298f
C41145 VPWR.t2678 VGND 0.05001f
C41146 VPWR.t1385 VGND 0.05001f
C41147 VPWR.t4097 VGND 0.05001f
C41148 VPWR.t823 VGND 0.05001f
C41149 VPWR.t1159 VGND 0.04521f
C41150 VPWR.t6268 VGND 0.0173f
C41151 VPWR.t570 VGND 0.05001f
C41152 VPWR.t1712 VGND 0.05001f
C41153 VPWR.t1553 VGND 0.04521f
C41154 VPWR.t5757 VGND 0.01172f
C41155 VPWR.t4205 VGND 0.02969f
C41156 VPWR.t165 VGND 0.04309f
C41157 VPWR.t4527 VGND 0.02992f
C41158 VPWR.t3848 VGND 0.04521f
C41159 VPWR.t4441 VGND 0.0173f
C41160 VPWR.t4888 VGND 0.05001f
C41161 VPWR.t4340 VGND 0.06143f
C41162 VPWR.t4889 VGND 0.00433f
C41163 VPWR.t4442 VGND 0.00433f
C41164 VPWR.t4528 VGND 0.00433f
C41165 VPWR.t166 VGND 0.00183f
C41166 VPWR.t3849 VGND 0.00157f
C41167 VPWR.n635 VGND 0.00508f
C41168 VPWR.t5758 VGND 0.00433f
C41169 VPWR.t4206 VGND 0.00203f
C41170 VPWR.t1554 VGND 0.00433f
C41171 VPWR.t1713 VGND 0.00433f
C41172 VPWR.t571 VGND 0.00433f
C41173 VPWR.t6269 VGND 0.00433f
C41174 VPWR.t1160 VGND 0.00433f
C41175 VPWR.t824 VGND 0.00433f
C41176 VPWR.n636 VGND 0.01085f
C41177 VPWR.n637 VGND 0.01085f
C41178 VPWR.n638 VGND 0.01085f
C41179 VPWR.n639 VGND 0.00676f
C41180 VPWR.n640 VGND 0.00974f
C41181 VPWR.n641 VGND 0.00788f
C41182 VPWR.n642 VGND 0.00684f
C41183 VPWR.n643 VGND 0.00974f
C41184 VPWR.n644 VGND 0.00659f
C41185 VPWR.n645 VGND 0.01284f
C41186 VPWR.n646 VGND 0.00544f
C41187 VPWR.n647 VGND 0.00758f
C41188 VPWR.n648 VGND 0.01189f
C41189 VPWR.n649 VGND 0.01144f
C41190 VPWR.n650 VGND 0.01085f
C41191 VPWR.n651 VGND 0.01085f
C41192 VPWR.n652 VGND 0.01023f
C41193 VPWR.n653 VGND 0.00974f
C41194 VPWR.n654 VGND 0.01085f
C41195 VPWR.n655 VGND 0.01085f
C41196 VPWR.n656 VGND 0.01085f
C41197 VPWR.n657 VGND 0.0085f
C41198 VPWR.n658 VGND 0.008f
C41199 VPWR.n659 VGND 0.00661f
C41200 VPWR.n660 VGND 0.00913f
C41201 VPWR.n661 VGND 0.00735f
C41202 VPWR.n662 VGND 0.00992f
C41203 VPWR.n663 VGND 0.00778f
C41204 VPWR.n664 VGND 0.00912f
C41205 VPWR.n665 VGND 0.01189f
C41206 VPWR.n666 VGND 0.01008f
C41207 VPWR.n667 VGND 0.01015f
C41208 VPWR.n668 VGND 0.00411f
C41209 VPWR.n669 VGND 0.01066f
C41210 VPWR.n670 VGND 0.00375f
C41211 VPWR.n671 VGND 0.00782f
C41212 VPWR.n672 VGND 0.0105f
C41213 VPWR.n673 VGND 0.01102f
C41214 VPWR.n674 VGND 0.01433f
C41215 VPWR.n675 VGND 0.00564f
C41216 VPWR.n676 VGND 0.00676f
C41217 VPWR.n677 VGND 0.00904f
C41218 VPWR.n678 VGND 0.008f
C41219 VPWR.n679 VGND 0.01071f
C41220 VPWR.n680 VGND 0.00467f
C41221 VPWR.n681 VGND 0.01091f
C41222 VPWR.n682 VGND 0.0017f
C41223 VPWR.n683 VGND 0.00883f
C41224 VPWR.n684 VGND 0.0036f
C41225 VPWR.n685 VGND 0.00798f
C41226 VPWR.n686 VGND 0.00986f
C41227 VPWR.n687 VGND 0.01015f
C41228 VPWR.n688 VGND 0.00665f
C41229 VPWR.n689 VGND 0.01152f
C41230 VPWR.n690 VGND 0.01158f
C41231 VPWR.n691 VGND 0.01251f
C41232 VPWR.n692 VGND 0.0071f
C41233 VPWR.n693 VGND 0.00551f
C41234 VPWR.n694 VGND 0.01009f
C41235 VPWR.n695 VGND 0.00671f
C41236 VPWR.n696 VGND 0.00808f
C41237 VPWR.n697 VGND 0.13412f
C41238 VPWR.t5595 VGND 0.00132f
C41239 VPWR.t5597 VGND 0.00132f
C41240 VPWR.n698 VGND 0.00266f
C41241 VPWR.n699 VGND 0.01081f
C41242 VPWR.t2544 VGND 0.00132f
C41243 VPWR.t2540 VGND 0.00132f
C41244 VPWR.n700 VGND 0.00266f
C41245 VPWR.t2458 VGND 0.00226f
C41246 VPWR.t2456 VGND 0.00163f
C41247 VPWR.n701 VGND 0.00392f
C41248 VPWR.t5593 VGND 0.00332f
C41249 VPWR.t279 VGND 0.0202f
C41250 VPWR.t286 VGND 0.00164f
C41251 VPWR.t280 VGND 0.00227f
C41252 VPWR.n702 VGND 0.00392f
C41253 VPWR.t2919 VGND 0.00433f
C41254 VPWR.t288 VGND 0.00164f
C41255 VPWR.t282 VGND 0.00227f
C41256 VPWR.n703 VGND 0.00392f
C41257 VPWR.t296 VGND 0.00164f
C41258 VPWR.t284 VGND 0.00227f
C41259 VPWR.n704 VGND 0.00392f
C41260 VPWR.t126 VGND 0.00431f
C41261 VPWR.t298 VGND 0.00164f
C41262 VPWR.t238 VGND 0.00227f
C41263 VPWR.n705 VGND 0.00392f
C41264 VPWR.t5588 VGND 0.00187f
C41265 VPWR.t2806 VGND 0.00139f
C41266 VPWR.n706 VGND 0.00471f
C41267 VPWR.t6831 VGND 0.00229f
C41268 VPWR.t240 VGND 0.00173f
C41269 VPWR.n707 VGND 0.00485f
C41270 VPWR.t244 VGND 0.00296f
C41271 VPWR.t6845 VGND 0.0011f
C41272 VPWR.t6843 VGND 0.00153f
C41273 VPWR.n708 VGND 0.00265f
C41274 VPWR.t256 VGND 0.00153f
C41275 VPWR.t250 VGND 0.0011f
C41276 VPWR.n709 VGND 0.00265f
C41277 VPWR.t6835 VGND 0.0011f
C41278 VPWR.t6839 VGND 0.00153f
C41279 VPWR.n710 VGND 0.00265f
C41280 VPWR.t264 VGND 0.00153f
C41281 VPWR.t262 VGND 0.0011f
C41282 VPWR.n711 VGND 0.00265f
C41283 VPWR.t6833 VGND 0.0011f
C41284 VPWR.t6837 VGND 0.00153f
C41285 VPWR.n712 VGND 0.00265f
C41286 VPWR.t274 VGND 0.00153f
C41287 VPWR.t260 VGND 0.0011f
C41288 VPWR.n713 VGND 0.00265f
C41289 VPWR.t6841 VGND 0.00296f
C41290 VPWR.t285 VGND 0.0173f
C41291 VPWR.t2918 VGND 0.025f
C41292 VPWR.t281 VGND 0.03907f
C41293 VPWR.t287 VGND 0.04041f
C41294 VPWR.t3307 VGND 0.025f
C41295 VPWR.t283 VGND 0.02612f
C41296 VPWR.t125 VGND 0.025f
C41297 VPWR.t295 VGND 0.01172f
C41298 VPWR.t237 VGND 0.0317f
C41299 VPWR.t2805 VGND 0.025f
C41300 VPWR.t297 VGND 0.03036f
C41301 VPWR.t5587 VGND 0.025f
C41302 VPWR.t239 VGND 0.02277f
C41303 VPWR.t4794 VGND 0.02824f
C41304 VPWR.t6830 VGND 0.0154f
C41305 VPWR.t6842 VGND 0.01172f
C41306 VPWR.t243 VGND 0.025f
C41307 VPWR.t6844 VGND 0.025f
C41308 VPWR.t249 VGND 0.025f
C41309 VPWR.t6838 VGND 0.025f
C41310 VPWR.t255 VGND 0.025f
C41311 VPWR.t6834 VGND 0.025f
C41312 VPWR.t261 VGND 0.025f
C41313 VPWR.t6836 VGND 0.025f
C41314 VPWR.t263 VGND 0.025f
C41315 VPWR.t6832 VGND 0.025f
C41316 VPWR.t259 VGND 0.025f
C41317 VPWR.t6840 VGND 0.025f
C41318 VPWR.t273 VGND 0.01172f
C41319 VPWR.t269 VGND 0.0202f
C41320 VPWR.n714 VGND 0.03274f
C41321 VPWR.t6571 VGND 0.00173f
C41322 VPWR.t270 VGND 0.00229f
C41323 VPWR.n715 VGND 0.00485f
C41324 VPWR.t124 VGND 0.00159f
C41325 VPWR.t1795 VGND 0.00158f
C41326 VPWR.n716 VGND 0.00497f
C41327 VPWR.t6549 VGND 0.00227f
C41328 VPWR.t6543 VGND 0.00164f
C41329 VPWR.n717 VGND 0.00392f
C41330 VPWR.t6551 VGND 0.00227f
C41331 VPWR.t6545 VGND 0.00164f
C41332 VPWR.n718 VGND 0.00392f
C41333 VPWR.t6559 VGND 0.00227f
C41334 VPWR.t6557 VGND 0.00164f
C41335 VPWR.n719 VGND 0.00392f
C41336 VPWR.t5962 VGND 0.00498f
C41337 VPWR.t6561 VGND 0.00227f
C41338 VPWR.t6563 VGND 0.00164f
C41339 VPWR.n720 VGND 0.00392f
C41340 VPWR.t6565 VGND 0.00227f
C41341 VPWR.t6567 VGND 0.00164f
C41342 VPWR.n721 VGND 0.00392f
C41343 VPWR.t192 VGND 0.00473f
C41344 VPWR.t6573 VGND 0.00227f
C41345 VPWR.t6569 VGND 0.00164f
C41346 VPWR.n722 VGND 0.00392f
C41347 VPWR.t4909 VGND 0.00434f
C41348 VPWR.t6555 VGND 0.00227f
C41349 VPWR.t6553 VGND 0.00164f
C41350 VPWR.n723 VGND 0.00392f
C41351 VPWR.t3962 VGND 0.00516f
C41352 VPWR.t6547 VGND 0.00425f
C41353 VPWR.t6570 VGND 0.03505f
C41354 VPWR.t1794 VGND 0.025f
C41355 VPWR.t6542 VGND 0.02902f
C41356 VPWR.t123 VGND 0.025f
C41357 VPWR.t6548 VGND 0.02902f
C41358 VPWR.t6981 VGND 0.025f
C41359 VPWR.t6544 VGND 0.025f
C41360 VPWR.t3310 VGND 0.025f
C41361 VPWR.t6550 VGND 0.01172f
C41362 VPWR.t6556 VGND 0.025f
C41363 VPWR.t6558 VGND 0.01395f
C41364 VPWR.t5961 VGND 0.025f
C41365 VPWR.t6562 VGND 0.025f
C41366 VPWR.t6617 VGND 0.025f
C41367 VPWR.t6560 VGND 0.025f
C41368 VPWR.t3840 VGND 0.025f
C41369 VPWR.t6566 VGND 0.02277f
C41370 VPWR.t191 VGND 0.025f
C41371 VPWR.t6564 VGND 0.03829f
C41372 VPWR.t6568 VGND 0.02824f
C41373 VPWR.t6572 VGND 0.02992f
C41374 VPWR.t4908 VGND 0.025f
C41375 VPWR.t6552 VGND 0.02724f
C41376 VPWR.t3311 VGND 0.025f
C41377 VPWR.t6554 VGND 0.02277f
C41378 VPWR.t3961 VGND 0.01886f
C41379 VPWR.t6546 VGND 0.0154f
C41380 VPWR.t5404 VGND 0.0298f
C41381 VPWR.n724 VGND 0.03642f
C41382 VPWR.t5405 VGND 0.00433f
C41383 VPWR.t503 VGND 0.00433f
C41384 VPWR.t6128 VGND 0.00433f
C41385 VPWR.t3256 VGND 0.00433f
C41386 VPWR.t1442 VGND 0.00433f
C41387 VPWR.t2163 VGND 0.00433f
C41388 VPWR.t1144 VGND 0.00433f
C41389 VPWR.t2920 VGND 0.00433f
C41390 VPWR.t1610 VGND 0.00433f
C41391 VPWR.t4538 VGND 0.00433f
C41392 VPWR.t5097 VGND 0.00433f
C41393 VPWR.t5071 VGND 0.00433f
C41394 VPWR.t1049 VGND 0.00473f
C41395 VPWR.t1588 VGND 0.00427f
C41396 VPWR.t1051 VGND 0.00427f
C41397 VPWR.t1590 VGND 0.00473f
C41398 VPWR.t4434 VGND 0.00473f
C41399 VPWR.t502 VGND 0.06731f
C41400 VPWR.t1441 VGND 0.10001f
C41401 VPWR.t1143 VGND 0.08271f
C41402 VPWR.t1609 VGND 0.05001f
C41403 VPWR.t4537 VGND 0.05001f
C41404 VPWR.t5070 VGND 0.025f
C41405 VPWR.t1048 VGND 0.0125f
C41406 VPWR.t1587 VGND 0.02288f
C41407 VPWR.t1050 VGND 0.02288f
C41408 VPWR.t1589 VGND 0.03538f
C41409 VPWR.t4433 VGND 0.03538f
C41410 VPWR.t4437 VGND 0.0298f
C41411 VPWR.n725 VGND 0.01544f
C41412 VPWR.t4438 VGND 0.00427f
C41413 VPWR.t1317 VGND 0.00427f
C41414 VPWR.t445 VGND 0.00433f
C41415 VPWR.t1315 VGND 0.00473f
C41416 VPWR.t1319 VGND 0.00427f
C41417 VPWR.n726 VGND 0.00766f
C41418 VPWR.n727 VGND 0.13412f
C41419 VPWR.t4335 VGND 0.00433f
C41420 VPWR.n728 VGND 0.0072f
C41421 VPWR.t4432 VGND 0.00473f
C41422 VPWR.t5739 VGND 0.00431f
C41423 VPWR.t4430 VGND 0.00427f
C41424 VPWR.n729 VGND 0.0276f
C41425 VPWR.t5741 VGND 0.00164f
C41426 VPWR.t4836 VGND 0.0029f
C41427 VPWR.n730 VGND 0.0047f
C41428 VPWR.t335 VGND 0.00431f
C41429 VPWR.t337 VGND 0.00164f
C41430 VPWR.t1592 VGND 0.0029f
C41431 VPWR.n731 VGND 0.0047f
C41432 VPWR.t3881 VGND 0.00164f
C41433 VPWR.t7024 VGND 0.00164f
C41434 VPWR.n732 VGND 0.00331f
C41435 VPWR.t2747 VGND 0.00427f
C41436 VPWR.t4436 VGND 0.00164f
C41437 VPWR.t7009 VGND 0.00164f
C41438 VPWR.n733 VGND 0.00331f
C41439 VPWR.t4834 VGND 0.00427f
C41440 VPWR.t2745 VGND 0.00473f
C41441 VPWR.t595 VGND 0.00433f
C41442 VPWR.t4832 VGND 0.00473f
C41443 VPWR.t5516 VGND 0.00433f
C41444 VPWR.t4568 VGND 0.00433f
C41445 VPWR.t4044 VGND 0.00433f
C41446 VPWR.t6755 VGND 0.00116f
C41447 VPWR.t6370 VGND 0.00116f
C41448 VPWR.n734 VGND 0.00236f
C41449 VPWR.t4080 VGND 0.00433f
C41450 VPWR.t3284 VGND 0.00255f
C41451 VPWR.t5740 VGND 0.0202f
C41452 VPWR.t334 VGND 0.01395f
C41453 VPWR.t4835 VGND 0.02389f
C41454 VPWR.t336 VGND 0.02858f
C41455 VPWR.t5737 VGND 0.02724f
C41456 VPWR.t1591 VGND 0.02277f
C41457 VPWR.t7020 VGND 0.01786f
C41458 VPWR.t3880 VGND 0.02724f
C41459 VPWR.t2499 VGND 0.02277f
C41460 VPWR.t7023 VGND 0.02277f
C41461 VPWR.t7013 VGND 0.02724f
C41462 VPWR.t4435 VGND 0.02221f
C41463 VPWR.t2746 VGND 0.01708f
C41464 VPWR.t7008 VGND 0.02791f
C41465 VPWR.t2744 VGND 0.03293f
C41466 VPWR.t4833 VGND 0.03963f
C41467 VPWR.t4831 VGND 0.03058f
C41468 VPWR.t594 VGND 0.03248f
C41469 VPWR.t5515 VGND 0.03271f
C41470 VPWR.t4567 VGND 0.0298f
C41471 VPWR.t4043 VGND 0.01395f
C41472 VPWR.t6754 VGND 0.03192f
C41473 VPWR.t6369 VGND 0.04085f
C41474 VPWR.t4079 VGND 0.03538f
C41475 VPWR.t3283 VGND 0.0202f
C41476 VPWR.n735 VGND 0.01968f
C41477 VPWR.t5508 VGND 0.00433f
C41478 VPWR.n736 VGND 0.00115f
C41479 VPWR.t18 VGND 0.00433f
C41480 VPWR.t2258 VGND 0.00107f
C41481 VPWR.n737 VGND 0.00292f
C41482 VPWR.t5847 VGND 0.00431f
C41483 VPWR.t2260 VGND 0.00427f
C41484 VPWR.t3309 VGND 0.00203f
C41485 VPWR.t182 VGND 0.00183f
C41486 VPWR.t4126 VGND 0.00157f
C41487 VPWR.n738 VGND 0.00508f
C41488 VPWR.t2478 VGND 0.00219f
C41489 VPWR.t13 VGND 0.00185f
C41490 VPWR.n739 VGND 0.00433f
C41491 VPWR.t4693 VGND 0.00159f
C41492 VPWR.t1022 VGND 0.00158f
C41493 VPWR.n740 VGND 0.00497f
C41494 VPWR.t5256 VGND 0.01733f
C41495 VPWR.n742 VGND 0.04381f
C41496 VPWR.t6371 VGND 0.01909f
C41497 VPWR.t5790 VGND 0.03014f
C41498 VPWR.t5507 VGND 0.02411f
C41499 VPWR.t5342 VGND 0.0173f
C41500 VPWR.t6372 VGND 0.01172f
C41501 VPWR.t17 VGND 0.03181f
C41502 VPWR.t3285 VGND 0.04867f
C41503 VPWR.t2261 VGND 0.0288f
C41504 VPWR.t906 VGND 0.02768f
C41505 VPWR.t2257 VGND 0.02612f
C41506 VPWR.t5846 VGND 0.02154f
C41507 VPWR.t2259 VGND 0.01172f
C41508 VPWR.t3308 VGND 0.03259f
C41509 VPWR.t181 VGND 0.04688f
C41510 VPWR.t119 VGND 0.02992f
C41511 VPWR.t4125 VGND 0.02277f
C41512 VPWR.t14 VGND 0.03974f
C41513 VPWR.t2477 VGND 0.03349f
C41514 VPWR.t1021 VGND 0.03125f
C41515 VPWR.t12 VGND 0.02902f
C41516 VPWR.t4692 VGND 0.02277f
C41517 VPWR.t118 VGND 0.02824f
C41518 VPWR.t6732 VGND 0.0125f
C41519 VPWR.t3841 VGND 0.0202f
C41520 VPWR.n743 VGND 0.01544f
C41521 VPWR.t3004 VGND 0.00425f
C41522 VPWR.t6980 VGND 0.00375f
C41523 VPWR.t3002 VGND 0.00227f
C41524 VPWR.t3008 VGND 0.00164f
C41525 VPWR.n744 VGND 0.00393f
C41526 VPWR.t3006 VGND 0.00401f
C41527 VPWR.t6743 VGND 0.0011f
C41528 VPWR.n745 VGND 0.00375f
C41529 VPWR.t6753 VGND 0.00296f
C41530 VPWR.t6983 VGND 0.00224f
C41531 VPWR.t775 VGND 0.00145f
C41532 VPWR.n746 VGND 0.00443f
C41533 VPWR.t117 VGND 0.00431f
C41534 VPWR.t777 VGND 0.00399f
C41535 VPWR.t5999 VGND 0.00394f
C41536 VPWR.t4227 VGND 0.00394f
C41537 VPWR.t6725 VGND 0.00394f
C41538 VPWR.t6727 VGND 0.00394f
C41539 VPWR.t6767 VGND 0.00116f
C41540 VPWR.t176 VGND 0.00116f
C41541 VPWR.n747 VGND 0.00236f
C41542 VPWR.t188 VGND 0.00287f
C41543 VPWR.t1620 VGND 0.00224f
C41544 VPWR.n748 VGND 0.00514f
C41545 VPWR.t6298 VGND 0.00255f
C41546 VPWR.t1622 VGND 0.00472f
C41547 VPWR.t3003 VGND 0.04097f
C41548 VPWR.t6979 VGND 0.02532f
C41549 VPWR.t3001 VGND 0.0283f
C41550 VPWR.t6500 VGND 0.02428f
C41551 VPWR.t3007 VGND 0.02428f
C41552 VPWR.t16 VGND 0.02428f
C41553 VPWR.t3005 VGND 0.02211f
C41554 VPWR.t20 VGND 0.02818f
C41555 VPWR.t6742 VGND 0.02428f
C41556 VPWR.t6503 VGND 0.02428f
C41557 VPWR.t6752 VGND 0.02832f
C41558 VPWR.t6982 VGND 0.01232f
C41559 VPWR.t774 VGND 0.01172f
C41560 VPWR.t116 VGND 0.02277f
C41561 VPWR.t776 VGND 0.02612f
C41562 VPWR.t3839 VGND 0.01395f
C41563 VPWR.t5998 VGND 0.025f
C41564 VPWR.t4226 VGND 0.02277f
C41565 VPWR.t6724 VGND 0.02277f
C41566 VPWR.t6726 VGND 0.025f
C41567 VPWR.t6766 VGND 0.01172f
C41568 VPWR.t187 VGND 0.02277f
C41569 VPWR.t175 VGND 0.02925f
C41570 VPWR.t1619 VGND 0.04175f
C41571 VPWR.t1621 VGND 0.03148f
C41572 VPWR.t6297 VGND 0.02244f
C41573 VPWR.t3630 VGND 0.01772f
C41574 VPWR.n749 VGND 0.03707f
C41575 VPWR.n750 VGND 0.00115f
C41576 VPWR.t3374 VGND 0.00427f
C41577 VPWR.t2960 VGND 0.00107f
C41578 VPWR.n751 VGND 0.00292f
C41579 VPWR.t4106 VGND 0.00107f
C41580 VPWR.n752 VGND 0.00292f
C41581 VPWR.t4108 VGND 0.00427f
C41582 VPWR.n753 VGND 0.00115f
C41583 VPWR.t4112 VGND 0.00603f
C41584 VPWR.t4691 VGND 0.00394f
C41585 VPWR.t6007 VGND 0.00255f
C41586 VPWR.t6430 VGND 0.00394f
C41587 VPWR.t144 VGND 0.00116f
C41588 VPWR.t6654 VGND 0.00116f
C41589 VPWR.n754 VGND 0.00236f
C41590 VPWR.t3268 VGND 0.00394f
C41591 VPWR.t6813 VGND 0.00394f
C41592 VPWR.t177 VGND 0.02478f
C41593 VPWR.t2650 VGND 0.02054f
C41594 VPWR.t3373 VGND 0.02411f
C41595 VPWR.t3631 VGND 0.03885f
C41596 VPWR.t2959 VGND 0.03338f
C41597 VPWR.t178 VGND 0.02768f
C41598 VPWR.t3371 VGND 0.03047f
C41599 VPWR.t6008 VGND 0.01875f
C41600 VPWR.t6296 VGND 0.01875f
C41601 VPWR.t4109 VGND 0.03047f
C41602 VPWR.t141 VGND 0.02768f
C41603 VPWR.t4105 VGND 0.03338f
C41604 VPWR.t4569 VGND 0.03885f
C41605 VPWR.t4107 VGND 0.02411f
C41606 VPWR.t2957 VGND 0.02054f
C41607 VPWR.t142 VGND 0.01875f
C41608 VPWR.t4111 VGND 0.00826f
C41609 VPWR.t5514 VGND 0.01775f
C41610 VPWR.n755 VGND 0.05865f
C41611 VPWR.t6006 VGND 0.0163f
C41612 VPWR.t4690 VGND 0.02311f
C41613 VPWR.t6429 VGND 0.0346f
C41614 VPWR.t143 VGND 0.0154f
C41615 VPWR.t6653 VGND 0.01183f
C41616 VPWR.t3267 VGND 0.01395f
C41617 VPWR.t6812 VGND 0.025f
C41618 VPWR.t819 VGND 0.0202f
C41619 VPWR.n756 VGND 0.04256f
C41620 VPWR.t820 VGND 0.00427f
C41621 VPWR.t5093 VGND 0.00433f
C41622 VPWR.t5463 VGND 0.00107f
C41623 VPWR.n757 VGND 0.00292f
C41624 VPWR.t3684 VGND 0.00433f
C41625 VPWR.t6032 VGND 0.00433f
C41626 VPWR.n758 VGND 0.00115f
C41627 VPWR.t7118 VGND 0.00433f
C41628 VPWR.t4149 VGND 0.00433f
C41629 VPWR.t3266 VGND 0.00255f
C41630 VPWR.t3971 VGND 0.00433f
C41631 VPWR.t223 VGND 0.00116f
C41632 VPWR.t6652 VGND 0.00116f
C41633 VPWR.n759 VGND 0.00236f
C41634 VPWR.t209 VGND 0.00431f
C41635 VPWR.t6864 VGND 0.00431f
C41636 VPWR.t3171 VGND 0.00433f
C41637 VPWR.t5462 VGND 0.03751f
C41638 VPWR.t5092 VGND 0.02768f
C41639 VPWR.t817 VGND 0.03684f
C41640 VPWR.t3264 VGND 0.03058f
C41641 VPWR.t3683 VGND 0.03047f
C41642 VPWR.t221 VGND 0.03271f
C41643 VPWR.t6031 VGND 0.03338f
C41644 VPWR.t525 VGND 0.02612f
C41645 VPWR.t5460 VGND 0.04063f
C41646 VPWR.t220 VGND 0.02389f
C41647 VPWR.t7117 VGND 0.02969f
C41648 VPWR.t2940 VGND 0.01775f
C41649 VPWR.n760 VGND 0.03208f
C41650 VPWR.t3265 VGND 0.0211f
C41651 VPWR.t4148 VGND 0.04822f
C41652 VPWR.t222 VGND 0.05001f
C41653 VPWR.t3970 VGND 0.02277f
C41654 VPWR.t6651 VGND 0.0173f
C41655 VPWR.t5117 VGND 0.025f
C41656 VPWR.t6863 VGND 0.01172f
C41657 VPWR.t208 VGND 0.01172f
C41658 VPWR.t6862 VGND 0.025f
C41659 VPWR.t2357 VGND 0.0202f
C41660 VPWR.t479 VGND 0.01574f
C41661 VPWR.t6540 VGND 0.02277f
C41662 VPWR.t3476 VGND 0.02277f
C41663 VPWR.t3482 VGND 0.02768f
C41664 VPWR.t6769 VGND 0.05626f
C41665 VPWR.t3182 VGND 0.03784f
C41666 VPWR.t3357 VGND 0.02735f
C41667 VPWR.t480 VGND 0.03282f
C41668 VPWR.t3477 VGND 0.03996f
C41669 VPWR.t2091 VGND 0.02277f
C41670 VPWR.t6525 VGND 0.0173f
C41671 VPWR.t928 VGND 0.06731f
C41672 VPWR.t1573 VGND 0.08271f
C41673 VPWR.t397 VGND 0.06731f
C41674 VPWR.t490 VGND 0.08271f
C41675 VPWR.t3170 VGND 0.05372f
C41676 VPWR.t6149 VGND 0.00433f
C41677 VPWR.t491 VGND 0.00433f
C41678 VPWR.t398 VGND 0.00433f
C41679 VPWR.t2684 VGND 0.00433f
C41680 VPWR.t6247 VGND 0.00433f
C41681 VPWR.t1574 VGND 0.00433f
C41682 VPWR.t2304 VGND 0.00433f
C41683 VPWR.t929 VGND 0.00433f
C41684 VPWR.t2092 VGND 0.00433f
C41685 VPWR.n761 VGND 0.00145f
C41686 VPWR.t3358 VGND 0.00433f
C41687 VPWR.n762 VGND 0.00831f
C41688 VPWR.n763 VGND 0.00811f
C41689 VPWR.n764 VGND 0.00819f
C41690 VPWR.n765 VGND 0.02059f
C41691 VPWR.n766 VGND 0.01588f
C41692 VPWR.n767 VGND 0.01476f
C41693 VPWR.n768 VGND 0.01562f
C41694 VPWR.n769 VGND 0.00893f
C41695 VPWR.n770 VGND 0.00792f
C41696 VPWR.n771 VGND 0.00792f
C41697 VPWR.n772 VGND 0.00561f
C41698 VPWR.n773 VGND 0.00992f
C41699 VPWR.n774 VGND 0.01013f
C41700 VPWR.n775 VGND 0.00893f
C41701 VPWR.n776 VGND 0.01247f
C41702 VPWR.n777 VGND 0.01011f
C41703 VPWR.n778 VGND 0.01507f
C41704 VPWR.n779 VGND 0.01197f
C41705 VPWR.n780 VGND 0.00809f
C41706 VPWR.n781 VGND 0.0093f
C41707 VPWR.n782 VGND 0.00647f
C41708 VPWR.n783 VGND 0.00928f
C41709 VPWR.n784 VGND 0.00727f
C41710 VPWR.n785 VGND 0.00804f
C41711 VPWR.n786 VGND 0.00432f
C41712 VPWR.n787 VGND 0.00411f
C41713 VPWR.n788 VGND 0.00834f
C41714 VPWR.n789 VGND 0.0064f
C41715 VPWR.n790 VGND 0.00993f
C41716 VPWR.n791 VGND 0.01492f
C41717 VPWR.n792 VGND 0.01029f
C41718 VPWR.n793 VGND 0.00938f
C41719 VPWR.n794 VGND 0.01721f
C41720 VPWR.n795 VGND 0.01721f
C41721 VPWR.n796 VGND 0.00938f
C41722 VPWR.n797 VGND 0.01035f
C41723 VPWR.n798 VGND 0.04341f
C41724 VPWR.n799 VGND 0.00971f
C41725 VPWR.n800 VGND 0.00833f
C41726 VPWR.n801 VGND 0.00593f
C41727 VPWR.n802 VGND 0.00466f
C41728 VPWR.n803 VGND 0.00936f
C41729 VPWR.n804 VGND 0.007f
C41730 VPWR.n805 VGND 0.007f
C41731 VPWR.n806 VGND 0.00803f
C41732 VPWR.n807 VGND 0.00868f
C41733 VPWR.n808 VGND 0.00811f
C41734 VPWR.n809 VGND 0.00431f
C41735 VPWR.n810 VGND 0.01025f
C41736 VPWR.n811 VGND 0.00551f
C41737 VPWR.n812 VGND 0.01054f
C41738 VPWR.n813 VGND 0.01201f
C41739 VPWR.n814 VGND 0.00812f
C41740 VPWR.n815 VGND 0.01288f
C41741 VPWR.n816 VGND 0.00615f
C41742 VPWR.n817 VGND 0.20174f
C41743 VPWR.t6506 VGND 0.00433f
C41744 VPWR.n818 VGND 0.00722f
C41745 VPWR.t226 VGND 0.00394f
C41746 VPWR.t218 VGND 0.00473f
C41747 VPWR.t4360 VGND 0.00394f
C41748 VPWR.t7038 VGND 0.00394f
C41749 VPWR.n819 VGND 0.03162f
C41750 VPWR.t3828 VGND 0.00394f
C41751 VPWR.t6730 VGND 0.00374f
C41752 VPWR.t909 VGND 0.00431f
C41753 VPWR.t4221 VGND 0.00132f
C41754 VPWR.t6502 VGND 0.00132f
C41755 VPWR.n820 VGND 0.00266f
C41756 VPWR.t7036 VGND 0.00132f
C41757 VPWR.t4223 VGND 0.00132f
C41758 VPWR.n821 VGND 0.00266f
C41759 VPWR.t6721 VGND 0.0033f
C41760 VPWR.t644 VGND 0.00431f
C41761 VPWR.t2448 VGND 0.00431f
C41762 VPWR.t646 VGND 0.00431f
C41763 VPWR.t4225 VGND 0.00433f
C41764 VPWR.t1323 VGND 0.00394f
C41765 VPWR.t6799 VGND 0.00394f
C41766 VPWR.t7037 VGND 0.0298f
C41767 VPWR.t3827 VGND 0.0125f
C41768 VPWR.t6729 VGND 0.0125f
C41769 VPWR.t908 VGND 0.02244f
C41770 VPWR.t4220 VGND 0.02277f
C41771 VPWR.t3949 VGND 0.02277f
C41772 VPWR.t6501 VGND 0.025f
C41773 VPWR.t1056 VGND 0.02277f
C41774 VPWR.t7035 VGND 0.025f
C41775 VPWR.t15 VGND 0.02277f
C41776 VPWR.t4222 VGND 0.02679f
C41777 VPWR.t6720 VGND 0.03427f
C41778 VPWR.t643 VGND 0.03672f
C41779 VPWR.t3950 VGND 0.03393f
C41780 VPWR.t7039 VGND 0.025f
C41781 VPWR.t4219 VGND 0.025f
C41782 VPWR.t3825 VGND 0.025f
C41783 VPWR.t6504 VGND 0.025f
C41784 VPWR.t4698 VGND 0.03393f
C41785 VPWR.t645 VGND 0.02712f
C41786 VPWR.t2447 VGND 0.02712f
C41787 VPWR.t5305 VGND 0.03393f
C41788 VPWR.t4224 VGND 0.02288f
C41789 VPWR.t1490 VGND 0.0154f
C41790 VPWR.t1322 VGND 0.0346f
C41791 VPWR.n822 VGND 0.04725f
C41792 VPWR.t4229 VGND 0.00433f
C41793 VPWR.t5633 VGND 0.00433f
C41794 VPWR.t3730 VGND 0.00163f
C41795 VPWR.t212 VGND 0.00163f
C41796 VPWR.n823 VGND 0.00329f
C41797 VPWR.t6815 VGND 0.00472f
C41798 VPWR.t5398 VGND 0.00433f
C41799 VPWR.t6809 VGND 0.00431f
C41800 VPWR.t5706 VGND 0.00433f
C41801 VPWR.t6304 VGND 0.00427f
C41802 VPWR.t3749 VGND 0.00433f
C41803 VPWR.t1652 VGND 0.00107f
C41804 VPWR.n824 VGND 0.00292f
C41805 VPWR.t3147 VGND 0.00433f
C41806 VPWR.t6126 VGND 0.00433f
C41807 VPWR.n825 VGND 0.00115f
C41808 VPWR.t3417 VGND 0.00433f
C41809 VPWR.t299 VGND 0.01733f
C41810 VPWR.t803 VGND 0.03751f
C41811 VPWR.t4228 VGND 0.02277f
C41812 VPWR.t3826 VGND 0.03137f
C41813 VPWR.t3729 VGND 0.04141f
C41814 VPWR.t5632 VGND 0.02277f
C41815 VPWR.t211 VGND 0.0173f
C41816 VPWR.t6814 VGND 0.03271f
C41817 VPWR.t5397 VGND 0.025f
C41818 VPWR.t6808 VGND 0.0298f
C41819 VPWR.t5705 VGND 0.03561f
C41820 VPWR.t6303 VGND 0.0173f
C41821 VPWR.t3748 VGND 0.03695f
C41822 VPWR.t1651 VGND 0.03192f
C41823 VPWR.t6305 VGND 0.0451f
C41824 VPWR.t1519 VGND 0.01808f
C41825 VPWR.t3146 VGND 0.03181f
C41826 VPWR.t7098 VGND 0.05001f
C41827 VPWR.t6125 VGND 0.03338f
C41828 VPWR.t2979 VGND 0.03862f
C41829 VPWR.t1625 VGND 0.0355f
C41830 VPWR.t3416 VGND 0.01652f
C41831 VPWR.t7099 VGND 0.01339f
C41832 VPWR.n827 VGND 0.02734f
C41833 VPWR.t1521 VGND 0.00255f
C41834 VPWR.t5497 VGND 0.00433f
C41835 VPWR.t7097 VGND 0.00116f
C41836 VPWR.t6499 VGND 0.00116f
C41837 VPWR.n828 VGND 0.00236f
C41838 VPWR.t5169 VGND 0.00433f
C41839 VPWR.t3599 VGND 0.00164f
C41840 VPWR.t3141 VGND 0.00347f
C41841 VPWR.n829 VGND 0.00515f
C41842 VPWR.t5870 VGND 0.00433f
C41843 VPWR.t3139 VGND 0.00164f
C41844 VPWR.t3143 VGND 0.00227f
C41845 VPWR.n830 VGND 0.00395f
C41846 VPWR.t5356 VGND 0.00433f
C41847 VPWR.t5806 VGND 0.00427f
C41848 VPWR.t4050 VGND 0.00219f
C41849 VPWR.t6719 VGND 0.00185f
C41850 VPWR.n831 VGND 0.00433f
C41851 VPWR.t1012 VGND 0.00107f
C41852 VPWR.n832 VGND 0.00292f
C41853 VPWR.t1520 VGND 0.025f
C41854 VPWR.t7096 VGND 0.03271f
C41855 VPWR.t5496 VGND 0.02277f
C41856 VPWR.t6498 VGND 0.0298f
C41857 VPWR.t5168 VGND 0.01172f
C41858 VPWR.t3598 VGND 0.0173f
C41859 VPWR.t3140 VGND 0.03829f
C41860 VPWR.t5869 VGND 0.025f
C41861 VPWR.t3138 VGND 0.01172f
C41862 VPWR.t3142 VGND 0.03271f
C41863 VPWR.t5355 VGND 0.03114f
C41864 VPWR.t6859 VGND 0.03561f
C41865 VPWR.t5805 VGND 0.02277f
C41866 VPWR.t6728 VGND 0.03393f
C41867 VPWR.t4049 VGND 0.02768f
C41868 VPWR.t1011 VGND 0.03125f
C41869 VPWR.t6718 VGND 0.02768f
C41870 VPWR.t5807 VGND 0.01875f
C41871 VPWR.t5487 VGND 0.02143f
C41872 VPWR.t6861 VGND 0.01797f
C41873 VPWR.t6612 VGND 0.025f
C41874 VPWR.t910 VGND 0.0202f
C41875 VPWR.n833 VGND 0.02783f
C41876 VPWR.n834 VGND 0.00115f
C41877 VPWR.t6536 VGND 0.00309f
C41878 VPWR.t5486 VGND 0.00255f
C41879 VPWR.t2349 VGND 0.00114f
C41880 VPWR.t2353 VGND 0.00306f
C41881 VPWR.n835 VGND 0.00423f
C41882 VPWR.t6614 VGND 0.00116f
C41883 VPWR.t6648 VGND 0.00116f
C41884 VPWR.n836 VGND 0.00236f
C41885 VPWR.t6532 VGND 0.00114f
C41886 VPWR.t6539 VGND 0.00114f
C41887 VPWR.n837 VGND 0.00231f
C41888 VPWR.t2362 VGND 0.00114f
C41889 VPWR.t2347 VGND 0.00306f
C41890 VPWR.n838 VGND 0.00423f
C41891 VPWR.t42 VGND 0.00374f
C41892 VPWR.t6534 VGND 0.00114f
C41893 VPWR.t3475 VGND 0.00114f
C41894 VPWR.n839 VGND 0.00231f
C41895 VPWR.t2355 VGND 0.00156f
C41896 VPWR.n840 VGND 0.00505f
C41897 VPWR.t6965 VGND 0.00114f
C41898 VPWR.t6974 VGND 0.00114f
C41899 VPWR.n841 VGND 0.00231f
C41900 VPWR.t47 VGND 0.0019f
C41901 VPWR.t3485 VGND 0.00114f
C41902 VPWR.t3480 VGND 0.00114f
C41903 VPWR.n842 VGND 0.00231f
C41904 VPWR.t111 VGND 0.00431f
C41905 VPWR.t6978 VGND 0.00114f
C41906 VPWR.t6976 VGND 0.00114f
C41907 VPWR.n843 VGND 0.00231f
C41908 VPWR.t4039 VGND 0.01733f
C41909 VPWR.t5009 VGND 0.0173f
C41910 VPWR.t6615 VGND 0.0211f
C41911 VPWR.n845 VGND 0.0181f
C41912 VPWR.t6535 VGND 0.03866f
C41913 VPWR.t5485 VGND 0.02277f
C41914 VPWR.t2348 VGND 0.0433f
C41915 VPWR.t2352 VGND 0.0357f
C41916 VPWR.t6613 VGND 0.02211f
C41917 VPWR.t6531 VGND 0.02211f
C41918 VPWR.t6647 VGND 0.01919f
C41919 VPWR.t6538 VGND 0.01214f
C41920 VPWR.t2361 VGND 0.03718f
C41921 VPWR.t41 VGND 0.03166f
C41922 VPWR.t2346 VGND 0.02873f
C41923 VPWR.t6533 VGND 0.03306f
C41924 VPWR.t2359 VGND 0.01605f
C41925 VPWR.t3474 VGND 0.02389f
C41926 VPWR.t2085 VGND 0.02277f
C41927 VPWR.t6964 VGND 0.02902f
C41928 VPWR.t2354 VGND 0.02277f
C41929 VPWR.t6973 VGND 0.02277f
C41930 VPWR.t46 VGND 0.02277f
C41931 VPWR.t3484 VGND 0.01485f
C41932 VPWR.t3479 VGND 0.01172f
C41933 VPWR.t110 VGND 0.02277f
C41934 VPWR.t6977 VGND 0.02612f
C41935 VPWR.t6537 VGND 0.02277f
C41936 VPWR.t6975 VGND 0.03505f
C41937 VPWR.t3468 VGND 0.02969f
C41938 VPWR.n846 VGND 0.01544f
C41939 VPWR.t3469 VGND 0.0031f
C41940 VPWR.t6999 VGND 0.00332f
C41941 VPWR.t2030 VGND 0.00456f
C41942 VPWR.t794 VGND 0.00132f
C41943 VPWR.t798 VGND 0.00132f
C41944 VPWR.n847 VGND 0.00266f
C41945 VPWR.t7001 VGND 0.00132f
C41946 VPWR.t6997 VGND 0.00132f
C41947 VPWR.n848 VGND 0.00266f
C41948 VPWR.t2034 VGND 0.00227f
C41949 VPWR.t2032 VGND 0.00227f
C41950 VPWR.n849 VGND 0.00463f
C41951 VPWR.t796 VGND 0.00132f
C41952 VPWR.t800 VGND 0.00132f
C41953 VPWR.n850 VGND 0.00266f
C41954 VPWR.t7003 VGND 0.00183f
C41955 VPWR.t5145 VGND 0.00166f
C41956 VPWR.n851 VGND 0.0043f
C41957 VPWR.t2028 VGND 0.00456f
C41958 VPWR.t5143 VGND 0.00147f
C41959 VPWR.t5139 VGND 0.00147f
C41960 VPWR.n852 VGND 0.00295f
C41961 VPWR.t7113 VGND 0.00433f
C41962 VPWR.t5141 VGND 0.00379f
C41963 VPWR.t6998 VGND 0.0154f
C41964 VPWR.t793 VGND 0.01395f
C41965 VPWR.t2029 VGND 0.02277f
C41966 VPWR.t797 VGND 0.02277f
C41967 VPWR.t6792 VGND 0.02277f
C41968 VPWR.t7000 VGND 0.02724f
C41969 VPWR.t6783 VGND 0.02277f
C41970 VPWR.t6996 VGND 0.02277f
C41971 VPWR.t2033 VGND 0.02277f
C41972 VPWR.t795 VGND 0.02724f
C41973 VPWR.t2031 VGND 0.02277f
C41974 VPWR.t799 VGND 0.02277f
C41975 VPWR.t6784 VGND 0.02277f
C41976 VPWR.t7002 VGND 0.02724f
C41977 VPWR.t6777 VGND 0.02724f
C41978 VPWR.t5144 VGND 0.02342f
C41979 VPWR.t2027 VGND 0.02828f
C41980 VPWR.t6508 VGND 0.03436f
C41981 VPWR.t6511 VGND 0.03241f
C41982 VPWR.t5142 VGND 0.03122f
C41983 VPWR.t7112 VGND 0.01615f
C41984 VPWR.t5138 VGND 0.01496f
C41985 VPWR.t6574 VGND 0.01745f
C41986 VPWR.t6513 VGND 0.02211f
C41987 VPWR.t6625 VGND 0.02211f
C41988 VPWR.t6509 VGND 0.02211f
C41989 VPWR.t6623 VGND 0.02749f
C41990 VPWR.t5140 VGND 0.02429f
C41991 VPWR.t6577 VGND 0.01395f
C41992 VPWR.t2560 VGND 0.0202f
C41993 VPWR.t881 VGND 0.0211f
C41994 VPWR.t4085 VGND 0.02657f
C41995 VPWR.t6848 VGND 0.04554f
C41996 VPWR.t6410 VGND 0.01629f
C41997 VPWR.t5752 VGND 0.0404f
C41998 VPWR.t6412 VGND 0.03038f
C41999 VPWR.t6852 VGND 0.02428f
C42000 VPWR.t6846 VGND 0.01355f
C42001 VPWR.t979 VGND 0.02211f
C42002 VPWR.t6404 VGND 0.02211f
C42003 VPWR.t3581 VGND 0.02955f
C42004 VPWR.t6512 VGND 0.03352f
C42005 VPWR.t6408 VGND 0.01673f
C42006 VPWR.t6850 VGND 0.04911f
C42007 VPWR.t3582 VGND 0.02712f
C42008 VPWR.t3577 VGND 0.025f
C42009 VPWR.t3575 VGND 0.03751f
C42010 VPWR.t6774 VGND 0.02277f
C42011 VPWR.t3579 VGND 0.025f
C42012 VPWR.t5730 VGND 0.02902f
C42013 VPWR.t6576 VGND 0.025f
C42014 VPWR.t6995 VGND 0.02277f
C42015 VPWR.t6626 VGND 0.02277f
C42016 VPWR.t3101 VGND 0.02277f
C42017 VPWR.t6624 VGND 0.01183f
C42018 VPWR.t6575 VGND 0.0202f
C42019 VPWR.n853 VGND 0.02638f
C42020 VPWR.t3580 VGND 0.00161f
C42021 VPWR.t3576 VGND 0.00161f
C42022 VPWR.n854 VGND 0.00325f
C42023 VPWR.t6775 VGND 0.00429f
C42024 VPWR.t3578 VGND 0.00161f
C42025 VPWR.t3583 VGND 0.00161f
C42026 VPWR.n855 VGND 0.00325f
C42027 VPWR.t6851 VGND 0.00309f
C42028 VPWR.t6409 VGND 0.00114f
C42029 VPWR.t6405 VGND 0.00306f
C42030 VPWR.n856 VGND 0.00423f
C42031 VPWR.t980 VGND 0.00431f
C42032 VPWR.t6847 VGND 0.00114f
C42033 VPWR.t6853 VGND 0.00114f
C42034 VPWR.n857 VGND 0.00231f
C42035 VPWR.n858 VGND 0.0039f
C42036 VPWR.n859 VGND 0.01028f
C42037 VPWR.n860 VGND 0.00916f
C42038 VPWR.n861 VGND 0.0114f
C42039 VPWR.n862 VGND 0.00476f
C42040 VPWR.n863 VGND 0.00837f
C42041 VPWR.n864 VGND 0.01207f
C42042 VPWR.n865 VGND 0.01511f
C42043 VPWR.n866 VGND 0.01504f
C42044 VPWR.n867 VGND 0.01007f
C42045 VPWR.n868 VGND 0.00439f
C42046 VPWR.n869 VGND 0.0119f
C42047 VPWR.n870 VGND 0.00892f
C42048 VPWR.n871 VGND 0.00911f
C42049 VPWR.n872 VGND 0.00776f
C42050 VPWR.n873 VGND 0.0119f
C42051 VPWR.n874 VGND 0.0105f
C42052 VPWR.n875 VGND 0.0103f
C42053 VPWR.n876 VGND 0.0066f
C42054 VPWR.n877 VGND 0.00576f
C42055 VPWR.n878 VGND 0.00965f
C42056 VPWR.n879 VGND 0.00851f
C42057 VPWR.n880 VGND 0.00891f
C42058 VPWR.n881 VGND 0.00407f
C42059 VPWR.n882 VGND 0.0065f
C42060 VPWR.n883 VGND 0.0049f
C42061 VPWR.n884 VGND 0.00879f
C42062 VPWR.n885 VGND 0.00871f
C42063 VPWR.n886 VGND 0.00587f
C42064 VPWR.n887 VGND 0.01064f
C42065 VPWR.n888 VGND 0.00511f
C42066 VPWR.n889 VGND 0.00682f
C42067 VPWR.n890 VGND 0.00797f
C42068 VPWR.n891 VGND 0.00761f
C42069 VPWR.n892 VGND 0.00951f
C42070 VPWR.n893 VGND 0.01072f
C42071 VPWR.n894 VGND 0.00578f
C42072 VPWR.n895 VGND 0.00916f
C42073 VPWR.n896 VGND 0.01208f
C42074 VPWR.n897 VGND 0.00499f
C42075 VPWR.n898 VGND 0.01577f
C42076 VPWR.n899 VGND 0.00772f
C42077 VPWR.n900 VGND 0.00469f
C42078 VPWR.n901 VGND 0.00706f
C42079 VPWR.n902 VGND 0.01089f
C42080 VPWR.n903 VGND 0.00992f
C42081 VPWR.n904 VGND 0.00561f
C42082 VPWR.n905 VGND 0.00958f
C42083 VPWR.n906 VGND 0.00593f
C42084 VPWR.n907 VGND 0.03918f
C42085 VPWR.n908 VGND 0.01244f
C42086 VPWR.n909 VGND 0.00809f
C42087 VPWR.n910 VGND 0.01899f
C42088 VPWR.t6705 VGND 0.00186f
C42089 VPWR.t6695 VGND 0.00139f
C42090 VPWR.n911 VGND 0.00435f
C42091 VPWR.n912 VGND 0.02548f
C42092 VPWR.t1693 VGND 0.00296f
C42093 VPWR.t6697 VGND 0.00164f
C42094 VPWR.t6689 VGND 0.00164f
C42095 VPWR.n913 VGND 0.0033f
C42096 VPWR.t1691 VGND 0.0011f
C42097 VPWR.t4186 VGND 0.00401f
C42098 VPWR.n914 VGND 0.00375f
C42099 VPWR.t6683 VGND 0.00164f
C42100 VPWR.t6687 VGND 0.00164f
C42101 VPWR.n915 VGND 0.0033f
C42102 VPWR.t4184 VGND 0.00164f
C42103 VPWR.t4188 VGND 0.00227f
C42104 VPWR.n916 VGND 0.00393f
C42105 VPWR.t6693 VGND 0.00164f
C42106 VPWR.t6685 VGND 0.00164f
C42107 VPWR.n917 VGND 0.0033f
C42108 VPWR.t4182 VGND 0.00425f
C42109 VPWR.t6691 VGND 0.00425f
C42110 VPWR.t5924 VGND 0.00456f
C42111 VPWR.t5930 VGND 0.00141f
C42112 VPWR.t3230 VGND 0.00251f
C42113 VPWR.n918 VGND 0.0044f
C42114 VPWR.t5922 VGND 0.00227f
C42115 VPWR.t5920 VGND 0.00227f
C42116 VPWR.n919 VGND 0.00463f
C42117 VPWR.t6696 VGND 0.01172f
C42118 VPWR.t1692 VGND 0.02277f
C42119 VPWR.t6688 VGND 0.025f
C42120 VPWR.t1690 VGND 0.02724f
C42121 VPWR.t6682 VGND 0.02902f
C42122 VPWR.t4185 VGND 0.02277f
C42123 VPWR.t6686 VGND 0.025f
C42124 VPWR.t4183 VGND 0.02724f
C42125 VPWR.t6692 VGND 0.025f
C42126 VPWR.t4187 VGND 0.02277f
C42127 VPWR.t6684 VGND 0.025f
C42128 VPWR.t4181 VGND 0.02724f
C42129 VPWR.t6690 VGND 0.03427f
C42130 VPWR.t5923 VGND 0.0154f
C42131 VPWR.t6515 VGND 0.01395f
C42132 VPWR.t5929 VGND 0.02724f
C42133 VPWR.t6518 VGND 0.02679f
C42134 VPWR.t3229 VGND 0.02277f
C42135 VPWR.t5921 VGND 0.03907f
C42136 VPWR.n920 VGND 0.03095f
C42137 VPWR.t6523 VGND 0.00296f
C42138 VPWR.t6520 VGND 0.0011f
C42139 VPWR.t4961 VGND 0.00401f
C42140 VPWR.n921 VGND 0.00375f
C42141 VPWR.t5926 VGND 0.00456f
C42142 VPWR.t4963 VGND 0.00164f
C42143 VPWR.t4959 VGND 0.00227f
C42144 VPWR.n922 VGND 0.00393f
C42145 VPWR.t5919 VGND 0.0202f
C42146 VPWR.t6517 VGND 0.03672f
C42147 VPWR.t6519 VGND 0.02724f
C42148 VPWR.t6522 VGND 0.025f
C42149 VPWR.t5925 VGND 0.02679f
C42150 VPWR.t4960 VGND 0.02902f
C42151 VPWR.t4962 VGND 0.03907f
C42152 VPWR.n923 VGND 0.02872f
C42153 VPWR.t2045 VGND 0.00603f
C42154 VPWR.t4965 VGND 0.00425f
C42155 VPWR.t2049 VGND 0.00427f
C42156 VPWR.t6332 VGND 0.00456f
C42157 VPWR.t672 VGND 0.00107f
C42158 VPWR.n924 VGND 0.00292f
C42159 VPWR.t6334 VGND 0.00227f
C42160 VPWR.t6336 VGND 0.00227f
C42161 VPWR.n925 VGND 0.00463f
C42162 VPWR.n926 VGND 0.00115f
C42163 VPWR.t6330 VGND 0.00456f
C42164 VPWR.t107 VGND 0.00431f
C42165 VPWR.t669 VGND 0.00255f
C42166 VPWR.t7057 VGND 0.00116f
C42167 VPWR.t6469 VGND 0.00116f
C42168 VPWR.n927 VGND 0.00236f
C42169 VPWR.t146 VGND 0.00456f
C42170 VPWR.t6329 VGND 0.02147f
C42171 VPWR.t3561 VGND 0.01772f
C42172 VPWR.t4958 VGND 0.03594f
C42173 VPWR.t4964 VGND 0.0317f
C42174 VPWR.t2044 VGND 0.02947f
C42175 VPWR.t2048 VGND 0.02467f
C42176 VPWR.t6331 VGND 0.02154f
C42177 VPWR.t671 VGND 0.02277f
C42178 VPWR.t6789 VGND 0.02768f
C42179 VPWR.t2046 VGND 0.02724f
C42180 VPWR.t6780 VGND 0.01741f
C42181 VPWR.t670 VGND 0.02277f
C42182 VPWR.t6333 VGND 0.03181f
C42183 VPWR.t7054 VGND 0.02724f
C42184 VPWR.t6335 VGND 0.03338f
C42185 VPWR.t4937 VGND 0.02277f
C42186 VPWR.t6787 VGND 0.02411f
C42187 VPWR.t4655 VGND 0.02724f
C42188 VPWR.t6791 VGND 0.01652f
C42189 VPWR.t7055 VGND 0.01674f
C42190 VPWR.n928 VGND 0.03945f
C42191 VPWR.t668 VGND 0.0163f
C42192 VPWR.t106 VGND 0.03784f
C42193 VPWR.t3481 VGND 0.03617f
C42194 VPWR.t7056 VGND 0.03282f
C42195 VPWR.t6468 VGND 0.02712f
C42196 VPWR.t145 VGND 0.0125f
C42197 VPWR.t6788 VGND 0.0202f
C42198 VPWR.n929 VGND 0.03095f
C42199 VPWR.t3536 VGND 0.00603f
C42200 VPWR.t150 VGND 0.00227f
C42201 VPWR.t152 VGND 0.00227f
C42202 VPWR.n930 VGND 0.00463f
C42203 VPWR.t3534 VGND 0.00427f
C42204 VPWR.t3530 VGND 0.00107f
C42205 VPWR.n931 VGND 0.00292f
C42206 VPWR.t148 VGND 0.00456f
C42207 VPWR.t44 VGND 0.00431f
C42208 VPWR.n932 VGND 0.00115f
C42209 VPWR.t3292 VGND 0.00255f
C42210 VPWR.t851 VGND 0.01733f
C42211 VPWR.t6778 VGND 0.04264f
C42212 VPWR.t3535 VGND 0.02277f
C42213 VPWR.t149 VGND 0.02277f
C42214 VPWR.t3533 VGND 0.02724f
C42215 VPWR.t151 VGND 0.02902f
C42216 VPWR.t6779 VGND 0.03259f
C42217 VPWR.t3529 VGND 0.02724f
C42218 VPWR.t6790 VGND 0.02768f
C42219 VPWR.t3531 VGND 0.02277f
C42220 VPWR.t147 VGND 0.01741f
C42221 VPWR.t3290 VGND 0.03672f
C42222 VPWR.t94 VGND 0.03338f
C42223 VPWR.t43 VGND 0.03181f
C42224 VPWR.t4996 VGND 0.02277f
C42225 VPWR.t5777 VGND 0.02411f
C42226 VPWR.t4514 VGND 0.025f
C42227 VPWR.t6768 VGND 0.01652f
C42228 VPWR.t95 VGND 0.01898f
C42229 VPWR.n934 VGND 0.05118f
C42230 VPWR.t3291 VGND 0.0202f
C42231 VPWR.n935 VGND 0.05194f
C42232 VPWR.t97 VGND 0.00116f
C42233 VPWR.t6487 VGND 0.00116f
C42234 VPWR.n936 VGND 0.00236f
C42235 VPWR.t7137 VGND 0.00427f
C42236 VPWR.t2284 VGND 0.00107f
C42237 VPWR.n937 VGND 0.00292f
C42238 VPWR.t96 VGND 0.04041f
C42239 VPWR.t7136 VGND 0.02277f
C42240 VPWR.t6486 VGND 0.0269f
C42241 VPWR.t2283 VGND 0.0125f
C42242 VPWR.n938 VGND 0.03084f
C42243 VPWR.t3218 VGND 0.00427f
C42244 VPWR.n939 VGND 0.00115f
C42245 VPWR.t5052 VGND 0.00107f
C42246 VPWR.n940 VGND 0.00292f
C42247 VPWR.t1032 VGND 0.00255f
C42248 VPWR.n941 VGND 0.00115f
C42249 VPWR.t6368 VGND 0.00116f
C42250 VPWR.t6483 VGND 0.00116f
C42251 VPWR.n942 VGND 0.00236f
C42252 VPWR.t6773 VGND 0.00287f
C42253 VPWR.t888 VGND 0.00224f
C42254 VPWR.n943 VGND 0.00514f
C42255 VPWR.t1930 VGND 0.00255f
C42256 VPWR.t890 VGND 0.00472f
C42257 VPWR.t6868 VGND 0.00116f
C42258 VPWR.t6479 VGND 0.00116f
C42259 VPWR.n944 VGND 0.00236f
C42260 VPWR.t1423 VGND 0.01733f
C42261 VPWR.t6772 VGND 0.02147f
C42262 VPWR.t7134 VGND 0.0173f
C42263 VPWR.t1030 VGND 0.025f
C42264 VPWR.t6366 VGND 0.03561f
C42265 VPWR.t3217 VGND 0.03338f
C42266 VPWR.t1932 VGND 0.03572f
C42267 VPWR.t433 VGND 0.02724f
C42268 VPWR.t5051 VGND 0.01652f
C42269 VPWR.t6365 VGND 0.02771f
C42270 VPWR.t3219 VGND 0.03082f
C42271 VPWR.t1928 VGND 0.01304f
C42272 VPWR.t1927 VGND 0.0276f
C42273 VPWR.t1031 VGND 0.02836f
C42274 VPWR.t6865 VGND 0.04465f
C42275 VPWR.t1617 VGND 0.03695f
C42276 VPWR.t6367 VGND 0.02411f
C42277 VPWR.t1777 VGND 0.02277f
C42278 VPWR.t6482 VGND 0.01619f
C42279 VPWR.t6866 VGND 0.0086f
C42280 VPWR.n946 VGND 0.03228f
C42281 VPWR.t1929 VGND 0.01976f
C42282 VPWR.t887 VGND 0.0288f
C42283 VPWR.t889 VGND 0.04443f
C42284 VPWR.t6867 VGND 0.04219f
C42285 VPWR.t6478 VGND 0.02422f
C42286 VPWR.n947 VGND 0.02682f
C42287 VPWR.t4400 VGND 0.00427f
C42288 VPWR.t1162 VGND 0.00431f
C42289 VPWR.t5219 VGND 0.00107f
C42290 VPWR.n948 VGND 0.00292f
C42291 VPWR.t4882 VGND 0.00431f
C42292 VPWR.n949 VGND 0.00115f
C42293 VPWR.t2554 VGND 0.00203f
C42294 VPWR.t4880 VGND 0.0018f
C42295 VPWR.t5063 VGND 0.00181f
C42296 VPWR.n950 VGND 0.00494f
C42297 VPWR.t4038 VGND 0.00255f
C42298 VPWR.t159 VGND 0.00116f
C42299 VPWR.t6481 VGND 0.00116f
C42300 VPWR.n951 VGND 0.00236f
C42301 VPWR.t4296 VGND 0.01733f
C42302 VPWR.t2553 VGND 0.02341f
C42303 VPWR.t4399 VGND 0.0202f
C42304 VPWR.t1161 VGND 0.02154f
C42305 VPWR.t5218 VGND 0.02612f
C42306 VPWR.t6675 VGND 0.02768f
C42307 VPWR.t4397 VGND 0.0288f
C42308 VPWR.t4036 VGND 0.02288f
C42309 VPWR.t160 VGND 0.0154f
C42310 VPWR.t4881 VGND 0.01931f
C42311 VPWR.t5231 VGND 0.02612f
C42312 VPWR.t2559 VGND 0.02411f
C42313 VPWR.t2380 VGND 0.0221f
C42314 VPWR.t157 VGND 0.02478f
C42315 VPWR.n953 VGND 0.02762f
C42316 VPWR.t4879 VGND 0.01596f
C42317 VPWR.t4037 VGND 0.02992f
C42318 VPWR.t5062 VGND 0.04822f
C42319 VPWR.t158 VGND 0.04376f
C42320 VPWR.t6480 VGND 0.03672f
C42321 VPWR.t6680 VGND 0.0202f
C42322 VPWR.n954 VGND 0.02872f
C42323 VPWR.t1259 VGND 0.00431f
C42324 VPWR.t6447 VGND 0.00433f
C42325 VPWR.t1158 VGND 0.02835f
C42326 VPWR.t1258 VGND 0.02422f
C42327 VPWR.t6446 VGND 0.0202f
C42328 VPWR.n955 VGND 0.03352f
C42329 VPWR.t4495 VGND 0.00433f
C42330 VPWR.t3015 VGND 0.00433f
C42331 VPWR.t5261 VGND 0.00433f
C42332 VPWR.t6497 VGND 0.0014f
C42333 VPWR.t1361 VGND 0.00223f
C42334 VPWR.n956 VGND 0.00369f
C42335 VPWR.t6190 VGND 0.00433f
C42336 VPWR.t5019 VGND 0.00426f
C42337 VPWR.t2171 VGND 0.00433f
C42338 VPWR.t5015 VGND 0.00164f
C42339 VPWR.t5023 VGND 0.00164f
C42340 VPWR.n957 VGND 0.00329f
C42341 VPWR.t414 VGND 0.00132f
C42342 VPWR.t5671 VGND 0.00132f
C42343 VPWR.n958 VGND 0.00267f
C42344 VPWR.t5017 VGND 0.00224f
C42345 VPWR.t1949 VGND 0.00156f
C42346 VPWR.n959 VGND 0.00428f
C42347 VPWR.t2736 VGND 0.00334f
C42348 VPWR.t1947 VGND 0.00127f
C42349 VPWR.n960 VGND 0.00342f
C42350 VPWR.t6902 VGND 0.00187f
C42351 VPWR.t6066 VGND 0.00139f
C42352 VPWR.n961 VGND 0.00471f
C42353 VPWR.n962 VGND 0.00115f
C42354 VPWR.t4494 VGND 0.03271f
C42355 VPWR.t3014 VGND 0.0173f
C42356 VPWR.t6496 VGND 0.0298f
C42357 VPWR.t5260 VGND 0.02768f
C42358 VPWR.t1360 VGND 0.05001f
C42359 VPWR.t6189 VGND 0.05313f
C42360 VPWR.t5018 VGND 0.04219f
C42361 VPWR.t5014 VGND 0.03505f
C42362 VPWR.t2170 VGND 0.02277f
C42363 VPWR.t5022 VGND 0.0173f
C42364 VPWR.t5016 VGND 0.02724f
C42365 VPWR.t413 VGND 0.02512f
C42366 VPWR.t5670 VGND 0.02445f
C42367 VPWR.t1948 VGND 0.02277f
C42368 VPWR.t2735 VGND 0.02277f
C42369 VPWR.t1946 VGND 0.01473f
C42370 VPWR.t5020 VGND 0.0317f
C42371 VPWR.t6065 VGND 0.01741f
C42372 VPWR.t6099 VGND 0.03036f
C42373 VPWR.t6901 VGND 0.03181f
C42374 VPWR.t140 VGND 0.02277f
C42375 VPWR.t6900 VGND 0.03338f
C42376 VPWR.t1354 VGND 0.01518f
C42377 VPWR.t1177 VGND 0.01733f
C42378 VPWR.t2403 VGND 0.05001f
C42379 VPWR.t3074 VGND 0.06731f
C42380 VPWR.t6361 VGND 0.05447f
C42381 VPWR.t6674 VGND 0.03058f
C42382 VPWR.t2586 VGND 0.03784f
C42383 VPWR.t4117 VGND 0.0365f
C42384 VPWR.t2733 VGND 0.03271f
C42385 VPWR.t6490 VGND 0.01886f
C42386 VPWR.t6896 VGND 0.02277f
C42387 VPWR.t138 VGND 0.02277f
C42388 VPWR.t4389 VGND 0.03617f
C42389 VPWR.t6894 VGND 0.04331f
C42390 VPWR.t6097 VGND 0.02277f
C42391 VPWR.t2734 VGND 0.03954f
C42392 VPWR.n964 VGND 0.01942f
C42393 VPWR.t137 VGND 0.02478f
C42394 VPWR.t1356 VGND 0.01764f
C42395 VPWR.n965 VGND 0.02504f
C42396 VPWR.n966 VGND 0.01266f
C42397 VPWR.n967 VGND 0.01181f
C42398 VPWR.n968 VGND 0.01087f
C42399 VPWR.n969 VGND 0.00848f
C42400 VPWR.n970 VGND 0.00851f
C42401 VPWR.n971 VGND 0.00382f
C42402 VPWR.n972 VGND 0.00902f
C42403 VPWR.n973 VGND 0.01129f
C42404 VPWR.n974 VGND 0.01085f
C42405 VPWR.n975 VGND 0.01038f
C42406 VPWR.n976 VGND 0.00788f
C42407 VPWR.n977 VGND 0.00518f
C42408 VPWR.n978 VGND 0.01321f
C42409 VPWR.n979 VGND 0.01259f
C42410 VPWR.n980 VGND 0.00588f
C42411 VPWR.n981 VGND 0.01077f
C42412 VPWR.n982 VGND 0.00622f
C42413 VPWR.n983 VGND 0.00653f
C42414 VPWR.n984 VGND 0.00865f
C42415 VPWR.n985 VGND 0.00926f
C42416 VPWR.n986 VGND 0.00398f
C42417 VPWR.n987 VGND 0.01366f
C42418 VPWR.n988 VGND 0.00949f
C42419 VPWR.n989 VGND 0.01062f
C42420 VPWR.n990 VGND 0.00836f
C42421 VPWR.n991 VGND 0.00795f
C42422 VPWR.n992 VGND 0.00569f
C42423 VPWR.n993 VGND 0.00644f
C42424 VPWR.n994 VGND 0.01102f
C42425 VPWR.n995 VGND 0.00533f
C42426 VPWR.n996 VGND 0.00899f
C42427 VPWR.n997 VGND 0.00833f
C42428 VPWR.n998 VGND 0.01312f
C42429 VPWR.n999 VGND 0.00313f
C42430 VPWR.n1000 VGND 0.00918f
C42431 VPWR.n1001 VGND 0.0185f
C42432 VPWR.n1002 VGND 0.01584f
C42433 VPWR.n1003 VGND 0.00856f
C42434 VPWR.n1004 VGND 0.01227f
C42435 VPWR.n1005 VGND 0.01165f
C42436 VPWR.n1006 VGND 0.00482f
C42437 VPWR.n1007 VGND 0.00884f
C42438 VPWR.n1008 VGND 0.00846f
C42439 VPWR.n1009 VGND 0.01486f
C42440 VPWR.n1010 VGND 0.00647f
C42441 VPWR.n1011 VGND 0.01099f
C42442 VPWR.n1012 VGND 0.01328f
C42443 VPWR.n1013 VGND 0.01412f
C42444 VPWR.n1014 VGND 0.0134f
C42445 VPWR.n1015 VGND 0.011f
C42446 VPWR.n1016 VGND 0.00789f
C42447 VPWR.n1017 VGND 0.01283f
C42448 VPWR.n1018 VGND 0.00941f
C42449 VPWR.t1207 VGND 0.00456f
C42450 VPWR.t1205 VGND 0.00227f
C42451 VPWR.t1203 VGND 0.00227f
C42452 VPWR.n1019 VGND 0.00463f
C42453 VPWR.t1201 VGND 0.00456f
C42454 VPWR.t7108 VGND 0.00425f
C42455 VPWR.t2288 VGND 0.00433f
C42456 VPWR.t3660 VGND 0.03948f
C42457 VPWR.t3661 VGND 0.00456f
C42458 VPWR.t3665 VGND 0.00227f
C42459 VPWR.t3663 VGND 0.00227f
C42460 VPWR.n1020 VGND 0.00463f
C42461 VPWR.t3667 VGND 0.00456f
C42462 VPWR.t4315 VGND 0.0019f
C42463 VPWR.t4678 VGND 0.00156f
C42464 VPWR.n1021 VGND 0.00505f
C42465 VPWR.t4313 VGND 0.00374f
C42466 VPWR.t5549 VGND 0.00433f
C42467 VPWR.t1953 VGND 0.00433f
C42468 VPWR.t5298 VGND 0.00433f
C42469 VPWR.t5430 VGND 0.00433f
C42470 VPWR.t5530 VGND 0.00433f
C42471 VPWR.t2969 VGND 0.00433f
C42472 VPWR.t3065 VGND 0.00433f
C42473 VPWR.t1152 VGND 0.00433f
C42474 VPWR.t5548 VGND 0.04035f
C42475 VPWR.t1952 VGND 0.05996f
C42476 VPWR.t5297 VGND 0.05996f
C42477 VPWR.t5429 VGND 0.05996f
C42478 VPWR.t5529 VGND 0.05996f
C42479 VPWR.t2968 VGND 0.05996f
C42480 VPWR.t3064 VGND 0.05996f
C42481 VPWR.t1151 VGND 0.05247f
C42482 VPWR.n1022 VGND 0.03832f
C42483 VPWR.t2114 VGND 0.00251f
C42484 VPWR.t89 VGND 0.00141f
C42485 VPWR.n1023 VGND 0.0044f
C42486 VPWR.t2771 VGND 0.00431f
C42487 VPWR.n1024 VGND 0.00116f
C42488 VPWR.t4138 VGND 0.00529f
C42489 VPWR.n1025 VGND 0.00208f
C42490 VPWR.t6749 VGND 0.00433f
C42491 VPWR.t88 VGND 0.02443f
C42492 VPWR.t2113 VGND 0.03661f
C42493 VPWR.t2770 VGND 0.02998f
C42494 VPWR.t179 VGND 0.0257f
C42495 VPWR.t5455 VGND 0.02623f
C42496 VPWR.t5454 VGND 0.04176f
C42497 VPWR.t5969 VGND 0.04176f
C42498 VPWR.t5970 VGND 0.03333f
C42499 VPWR.t4137 VGND 0.05494f
C42500 VPWR.t6748 VGND 0.03989f
C42501 VPWR.n1026 VGND 0.02794f
C42502 VPWR.t9 VGND 0.00296f
C42503 VPWR.t4672 VGND 0.00401f
C42504 VPWR.t11 VGND 0.0011f
C42505 VPWR.n1027 VGND 0.00375f
C42506 VPWR.t4674 VGND 0.00227f
C42507 VPWR.t4676 VGND 0.00164f
C42508 VPWR.n1028 VGND 0.00393f
C42509 VPWR.t4670 VGND 0.00425f
C42510 VPWR.t3356 VGND 0.00433f
C42511 VPWR.t4829 VGND 0.00433f
C42512 VPWR.t6765 VGND 0.00431f
C42513 VPWR.t8 VGND 0.02202f
C42514 VPWR.t10 VGND 0.03239f
C42515 VPWR.t4671 VGND 0.03239f
C42516 VPWR.t4675 VGND 0.02998f
C42517 VPWR.t4673 VGND 0.02998f
C42518 VPWR.t4669 VGND 0.04926f
C42519 VPWR.t3355 VGND 0.04129f
C42520 VPWR.t4828 VGND 0.02998f
C42521 VPWR.t6764 VGND 0.02269f
C42522 VPWR.t7021 VGND 0.03795f
C42523 VPWR.n1029 VGND 0.0337f
C42524 VPWR.n1030 VGND 0.00116f
C42525 VPWR.t2922 VGND 0.00529f
C42526 VPWR.n1031 VGND 0.00208f
C42527 VPWR.n1032 VGND 0.03099f
C42528 VPWR.t324 VGND 0.00433f
C42529 VPWR.n1033 VGND 0.00677f
C42530 VPWR.t5271 VGND 0.00434f
C42531 VPWR.t6876 VGND 0.0298f
C42532 VPWR.t6637 VGND 0.00374f
C42533 VPWR.t2482 VGND 0.00473f
C42534 VPWR.t2484 VGND 0.00427f
C42535 VPWR.t6875 VGND 0.00156f
C42536 VPWR.n1034 VGND 0.00505f
C42537 VPWR.t5934 VGND 0.00473f
C42538 VPWR.t6630 VGND 0.0019f
C42539 VPWR.t5936 VGND 0.00427f
C42540 VPWR.t6636 VGND 0.03637f
C42541 VPWR.t2481 VGND 0.03097f
C42542 VPWR.t6873 VGND 0.02824f
C42543 VPWR.t2483 VGND 0.02389f
C42544 VPWR.t3409 VGND 0.01172f
C42545 VPWR.t6874 VGND 0.03538f
C42546 VPWR.t5933 VGND 0.02277f
C42547 VPWR.t6629 VGND 0.02712f
C42548 VPWR.t5935 VGND 0.0125f
C42549 VPWR.t6879 VGND 0.0173f
C42550 VPWR.n1035 VGND 0.02649f
C42551 VPWR.t4871 VGND 0.00163f
C42552 VPWR.t6880 VGND 0.00163f
C42553 VPWR.n1036 VGND 0.00328f
C42554 VPWR.t4869 VGND 0.00427f
C42555 VPWR.t4873 VGND 0.00473f
C42556 VPWR.t3790 VGND 0.00427f
C42557 VPWR.t5657 VGND 0.00433f
C42558 VPWR.t6342 VGND 0.00296f
C42559 VPWR.t3792 VGND 0.00473f
C42560 VPWR.t1106 VGND 0.00401f
C42561 VPWR.t6344 VGND 0.0011f
C42562 VPWR.n1037 VGND 0.00375f
C42563 VPWR.t4870 VGND 0.0202f
C42564 VPWR.t4868 VGND 0.02422f
C42565 VPWR.t7016 VGND 0.02791f
C42566 VPWR.t4872 VGND 0.02366f
C42567 VPWR.t1532 VGND 0.03326f
C42568 VPWR.t6635 VGND 0.02712f
C42569 VPWR.t5656 VGND 0.025f
C42570 VPWR.t3789 VGND 0.025f
C42571 VPWR.t3791 VGND 0.01172f
C42572 VPWR.t6341 VGND 0.0346f
C42573 VPWR.t6343 VGND 0.02579f
C42574 VPWR.t1105 VGND 0.0298f
C42575 VPWR.n1038 VGND 0.02548f
C42576 VPWR.t5661 VGND 0.00427f
C42577 VPWR.t1112 VGND 0.00227f
C42578 VPWR.t1108 VGND 0.00164f
C42579 VPWR.n1039 VGND 0.00393f
C42580 VPWR.t5663 VGND 0.00473f
C42581 VPWR.t1110 VGND 0.00425f
C42582 VPWR.t1742 VGND 0.00427f
C42583 VPWR.t2570 VGND 0.00427f
C42584 VPWR.t1744 VGND 0.00473f
C42585 VPWR.t2572 VGND 0.00473f
C42586 VPWR.t1213 VGND 0.00427f
C42587 VPWR.t5719 VGND 0.00427f
C42588 VPWR.t1217 VGND 0.00473f
C42589 VPWR.t5717 VGND 0.00473f
C42590 VPWR.t1531 VGND 0.00473f
C42591 VPWR.t1525 VGND 0.00427f
C42592 VPWR.t1529 VGND 0.00427f
C42593 VPWR.t1527 VGND 0.00473f
C42594 VPWR.t1107 VGND 0.01172f
C42595 VPWR.t5660 VGND 0.025f
C42596 VPWR.t1111 VGND 0.02791f
C42597 VPWR.t5662 VGND 0.025f
C42598 VPWR.t1109 VGND 0.03538f
C42599 VPWR.t1741 VGND 0.0125f
C42600 VPWR.t2569 VGND 0.02712f
C42601 VPWR.t1743 VGND 0.02791f
C42602 VPWR.t2571 VGND 0.03538f
C42603 VPWR.t1212 VGND 0.0125f
C42604 VPWR.t5718 VGND 0.02712f
C42605 VPWR.t1216 VGND 0.02791f
C42606 VPWR.t5716 VGND 0.04789f
C42607 VPWR.t1530 VGND 0.01172f
C42608 VPWR.t1524 VGND 0.02791f
C42609 VPWR.t1528 VGND 0.02791f
C42610 VPWR.t1526 VGND 0.01172f
C42611 VPWR.n1040 VGND 0.00443f
C42612 VPWR.n1041 VGND 0.00655f
C42613 VPWR.n1042 VGND 0.00655f
C42614 VPWR.n1043 VGND 0.00584f
C42615 VPWR.n1044 VGND 0.00698f
C42616 VPWR.n1045 VGND 0.0054f
C42617 VPWR.n1046 VGND 0.0077f
C42618 VPWR.n1047 VGND 0.00698f
C42619 VPWR.n1048 VGND 0.00584f
C42620 VPWR.n1049 VGND 0.0054f
C42621 VPWR.n1050 VGND 0.0077f
C42622 VPWR.n1051 VGND 0.00683f
C42623 VPWR.n1052 VGND 0.00679f
C42624 VPWR.n1053 VGND 0.00481f
C42625 VPWR.t1738 VGND 0.00427f
C42626 VPWR.n1054 VGND 0.00791f
C42627 VPWR.t1740 VGND 0.00473f
C42628 VPWR.n1055 VGND 0.00116f
C42629 VPWR.t1380 VGND 0.00529f
C42630 VPWR.n1056 VGND 0.00208f
C42631 VPWR.n1057 VGND 0.02508f
C42632 VPWR.n1058 VGND 0.01771f
C42633 VPWR.t6817 VGND 0.0257f
C42634 VPWR.t3321 VGND 0.02623f
C42635 VPWR.t3323 VGND 0.04176f
C42636 VPWR.t3324 VGND 0.04176f
C42637 VPWR.t3325 VGND 0.03333f
C42638 VPWR.t1379 VGND 0.03948f
C42639 VPWR.t1737 VGND 0.02376f
C42640 VPWR.t1739 VGND 0.04082f
C42641 VPWR.n1059 VGND 0.05029f
C42642 VPWR.t5284 VGND 0.00433f
C42643 VPWR.t6142 VGND 0.00425f
C42644 VPWR.t6140 VGND 0.00227f
C42645 VPWR.t6144 VGND 0.00164f
C42646 VPWR.n1060 VGND 0.00393f
C42647 VPWR.t6146 VGND 0.00401f
C42648 VPWR.t7051 VGND 0.0011f
C42649 VPWR.n1061 VGND 0.00375f
C42650 VPWR.t7053 VGND 0.00296f
C42651 VPWR.t2530 VGND 0.00223f
C42652 VPWR.t24 VGND 0.0014f
C42653 VPWR.n1062 VGND 0.00369f
C42654 VPWR.t5653 VGND 0.00223f
C42655 VPWR.t7 VGND 0.0014f
C42656 VPWR.n1063 VGND 0.00369f
C42657 VPWR.t5283 VGND 0.03286f
C42658 VPWR.t6141 VGND 0.03554f
C42659 VPWR.t6139 VGND 0.02998f
C42660 VPWR.t6143 VGND 0.02998f
C42661 VPWR.t6145 VGND 0.03239f
C42662 VPWR.t7050 VGND 0.03239f
C42663 VPWR.t7052 VGND 0.02202f
C42664 VPWR.t2529 VGND 0.03661f
C42665 VPWR.t23 VGND 0.02496f
C42666 VPWR.t5652 VGND 0.03661f
C42667 VPWR.t6 VGND 0.02496f
C42668 VPWR.t7048 VGND 0.0257f
C42669 VPWR.t3239 VGND 0.02623f
C42670 VPWR.t3241 VGND 0.04176f
C42671 VPWR.t5521 VGND 0.04176f
C42672 VPWR.t5519 VGND 0.03333f
C42673 VPWR.t2921 VGND 0.05113f
C42674 VPWR.t340 VGND 0.05113f
C42675 VPWR.t359 VGND 0.03333f
C42676 VPWR.t358 VGND 0.04176f
C42677 VPWR.t1436 VGND 0.04176f
C42678 VPWR.t1437 VGND 0.02623f
C42679 VPWR.t52 VGND 0.0257f
C42680 VPWR.n1064 VGND 0.02794f
C42681 VPWR.n1065 VGND 0.00116f
C42682 VPWR.t341 VGND 0.00529f
C42683 VPWR.n1066 VGND 0.00208f
C42684 VPWR.n1067 VGND 0.0311f
C42685 VPWR.n1068 VGND 0.01771f
C42686 VPWR.n1069 VGND 0.01511f
C42687 VPWR.n1070 VGND 0.01212f
C42688 VPWR.n1071 VGND 0.00849f
C42689 VPWR.n1072 VGND 0.01141f
C42690 VPWR.n1073 VGND 0.01202f
C42691 VPWR.n1074 VGND 0.01147f
C42692 VPWR.n1075 VGND 0.01594f
C42693 VPWR.n1076 VGND 0.00912f
C42694 VPWR.n1077 VGND 0.01189f
C42695 VPWR.n1078 VGND 0.00937f
C42696 VPWR.n1079 VGND 0.01555f
C42697 VPWR.t5908 VGND 0.00473f
C42698 VPWR.n1080 VGND 0.00519f
C42699 VPWR.t4509 VGND 0.00427f
C42700 VPWR.t3496 VGND 0.00433f
C42701 VPWR.t761 VGND 0.00433f
C42702 VPWR.t6177 VGND 0.00473f
C42703 VPWR.t2524 VGND 0.00473f
C42704 VPWR.t6176 VGND 0.00427f
C42705 VPWR.t2526 VGND 0.00427f
C42706 VPWR.t5906 VGND 0.00427f
C42707 VPWR.t3737 VGND 0.00427f
C42708 VPWR.t5905 VGND 0.00473f
C42709 VPWR.t3735 VGND 0.00473f
C42710 VPWR.t5910 VGND 0.00427f
C42711 VPWR.t4511 VGND 0.00473f
C42712 VPWR.n1081 VGND 0.00655f
C42713 VPWR.n1082 VGND 0.00672f
C42714 VPWR.n1083 VGND 0.01101f
C42715 VPWR.n1084 VGND 0.01353f
C42716 VPWR.n1085 VGND 0.01353f
C42717 VPWR.n1086 VGND 0.0117f
C42718 VPWR.t2523 VGND 0.06329f
C42719 VPWR.t2525 VGND 0.03963f
C42720 VPWR.t3736 VGND 0.03963f
C42721 VPWR.t3734 VGND 0.06039f
C42722 VPWR.t5909 VGND 0.03248f
C42723 VPWR.t4510 VGND 0.02791f
C42724 VPWR.t5907 VGND 0.02791f
C42725 VPWR.t4508 VGND 0.03248f
C42726 VPWR.t3495 VGND 0.03271f
C42727 VPWR.t760 VGND 0.0173f
C42728 VPWR.n1087 VGND 0.04122f
C42729 VPWR.t1536 VGND 0.00433f
C42730 VPWR.t4971 VGND 0.00433f
C42731 VPWR.t63 VGND 0.00433f
C42732 VPWR.t4410 VGND 0.00433f
C42733 VPWR.t4844 VGND 0.00433f
C42734 VPWR.t3969 VGND 0.00433f
C42735 VPWR.t1037 VGND 0.00433f
C42736 VPWR.t6138 VGND 0.00433f
C42737 VPWR.t5292 VGND 0.00433f
C42738 VPWR.t1860 VGND 0.00427f
C42739 VPWR.t3798 VGND 0.00433f
C42740 VPWR.t2779 VGND 0.00433f
C42741 VPWR.t1864 VGND 0.00473f
C42742 VPWR.t1400 VGND 0.00433f
C42743 VPWR.t3042 VGND 0.00433f
C42744 VPWR.t2753 VGND 0.00433f
C42745 VPWR.t5152 VGND 0.00433f
C42746 VPWR.t1535 VGND 0.025f
C42747 VPWR.t62 VGND 0.05001f
C42748 VPWR.t4409 VGND 0.08271f
C42749 VPWR.t1036 VGND 0.10001f
C42750 VPWR.t5291 VGND 0.06731f
C42751 VPWR.t1859 VGND 0.0173f
C42752 VPWR.t3797 VGND 0.02791f
C42753 VPWR.t1863 VGND 0.05001f
C42754 VPWR.t2778 VGND 0.05269f
C42755 VPWR.t1399 VGND 0.05001f
C42756 VPWR.t3041 VGND 0.05001f
C42757 VPWR.t2752 VGND 0.04231f
C42758 VPWR.t5151 VGND 0.0202f
C42759 VPWR.n1088 VGND 0.03352f
C42760 VPWR.t765 VGND 0.00433f
C42761 VPWR.t1582 VGND 0.00473f
C42762 VPWR.t3975 VGND 0.00427f
C42763 VPWR.t1586 VGND 0.00427f
C42764 VPWR.t3973 VGND 0.00473f
C42765 VPWR.t1685 VGND 0.00473f
C42766 VPWR.t1683 VGND 0.00427f
C42767 VPWR.t5111 VGND 0.00433f
C42768 VPWR.t2843 VGND 0.00433f
C42769 VPWR.t2498 VGND 0.00433f
C42770 VPWR.t538 VGND 0.00473f
C42771 VPWR.t6167 VGND 0.00433f
C42772 VPWR.t542 VGND 0.00427f
C42773 VPWR.t536 VGND 0.00427f
C42774 VPWR.t5614 VGND 0.00427f
C42775 VPWR.t540 VGND 0.00473f
C42776 VPWR.t5612 VGND 0.00473f
C42777 VPWR.t1223 VGND 0.00433f
C42778 VPWR.t764 VGND 0.03538f
C42779 VPWR.t1581 VGND 0.0173f
C42780 VPWR.t1585 VGND 0.01172f
C42781 VPWR.t3974 VGND 0.01172f
C42782 VPWR.t3972 VGND 0.03538f
C42783 VPWR.t1684 VGND 0.03248f
C42784 VPWR.t1682 VGND 0.0125f
C42785 VPWR.t5110 VGND 0.025f
C42786 VPWR.t2497 VGND 0.05001f
C42787 VPWR.t537 VGND 0.03829f
C42788 VPWR.t6166 VGND 0.01462f
C42789 VPWR.t535 VGND 0.0154f
C42790 VPWR.t541 VGND 0.0154f
C42791 VPWR.t5613 VGND 0.01462f
C42792 VPWR.t539 VGND 0.02791f
C42793 VPWR.t5611 VGND 0.03248f
C42794 VPWR.t1222 VGND 0.06623f
C42795 VPWR.t5025 VGND 0.00433f
C42796 VPWR.t3676 VGND 0.00433f
C42797 VPWR.t5801 VGND 0.00433f
C42798 VPWR.t876 VGND 0.00433f
C42799 VPWR.t3388 VGND 0.00433f
C42800 VPWR.t515 VGND 0.00433f
C42801 VPWR.t2177 VGND 0.00433f
C42802 VPWR.t6747 VGND 0.00116f
C42803 VPWR.t26 VGND 0.00116f
C42804 VPWR.n1089 VGND 0.00236f
C42805 VPWR.t2534 VGND 0.00433f
C42806 VPWR.t3984 VGND 0.00255f
C42807 VPWR.t2108 VGND 0.00433f
C42808 VPWR.t554 VGND 0.00433f
C42809 VPWR.n1090 VGND 0.00115f
C42810 VPWR.t937 VGND 0.00431f
C42811 VPWR.t2107 VGND 0.01566f
C42812 VPWR.t6069 VGND 0.02353f
C42813 VPWR.t5024 VGND 0.03271f
C42814 VPWR.t3675 VGND 0.0298f
C42815 VPWR.t5800 VGND 0.03271f
C42816 VPWR.t875 VGND 0.05001f
C42817 VPWR.t3387 VGND 0.05001f
C42818 VPWR.t514 VGND 0.0298f
C42819 VPWR.t2176 VGND 0.01395f
C42820 VPWR.t6746 VGND 0.03192f
C42821 VPWR.t25 VGND 0.04085f
C42822 VPWR.t2533 VGND 0.04822f
C42823 VPWR.t3983 VGND 0.0461f
C42824 VPWR.n1092 VGND 0.03945f
C42825 VPWR.t28 VGND 0.02478f
C42826 VPWR.t2932 VGND 0.01764f
C42827 VPWR.t553 VGND 0.01842f
C42828 VPWR.t2930 VGND 0.0154f
C42829 VPWR.t936 VGND 0.02366f
C42830 VPWR.t27 VGND 0.04085f
C42831 VPWR.t5589 VGND 0.0202f
C42832 VPWR.t3772 VGND 0.025f
C42833 VPWR.t907 VGND 0.01227f
C42834 VPWR.t1262 VGND 0.03024f
C42835 VPWR.t6795 VGND 0.03258f
C42836 VPWR.t5848 VGND 0.0154f
C42837 VPWR.t6802 VGND 0.02277f
C42838 VPWR.t5488 VGND 0.02277f
C42839 VPWR.t1268 VGND 0.04097f
C42840 VPWR.t938 VGND 0.01395f
C42841 VPWR.t129 VGND 0.02679f
C42842 VPWR.t183 VGND 0.02277f
C42843 VPWR.t186 VGND 0.025f
C42844 VPWR.t6616 VGND 0.02724f
C42845 VPWR.t1266 VGND 0.025f
C42846 VPWR.t134 VGND 0.02277f
C42847 VPWR.t6806 VGND 0.02902f
C42848 VPWR.t440 VGND 0.03829f
C42849 VPWR.t189 VGND 0.0125f
C42850 VPWR.t727 VGND 0.04521f
C42851 VPWR.t1294 VGND 0.02992f
C42852 VPWR.t5393 VGND 0.03885f
C42853 VPWR.t2285 VGND 0.03561f
C42854 VPWR.t1292 VGND 0.025f
C42855 VPWR.t3985 VGND 0.0173f
C42856 VPWR.n1093 VGND 0.03553f
C42857 VPWR.t2286 VGND 0.00107f
C42858 VPWR.n1094 VGND 0.00292f
C42859 VPWR.t1295 VGND 0.00427f
C42860 VPWR.t728 VGND 0.00183f
C42861 VPWR.t5394 VGND 0.00157f
C42862 VPWR.n1095 VGND 0.00508f
C42863 VPWR.t190 VGND 0.00203f
C42864 VPWR.t135 VGND 0.00159f
C42865 VPWR.t441 VGND 0.00158f
C42866 VPWR.n1096 VGND 0.00497f
C42867 VPWR.t6807 VGND 0.00132f
C42868 VPWR.t1267 VGND 0.00132f
C42869 VPWR.n1097 VGND 0.00266f
C42870 VPWR.t130 VGND 0.00516f
C42871 VPWR.t1269 VGND 0.00425f
C42872 VPWR.t5489 VGND 0.00438f
C42873 VPWR.n1098 VGND 0.01027f
C42874 VPWR.n1099 VGND 0.0079f
C42875 VPWR.n1100 VGND 0.01322f
C42876 VPWR.n1101 VGND 0.00601f
C42877 VPWR.n1102 VGND 0.00944f
C42878 VPWR.n1103 VGND 0.00793f
C42879 VPWR.n1104 VGND 0.00622f
C42880 VPWR.n1105 VGND 0.01065f
C42881 VPWR.n1106 VGND 0.00501f
C42882 VPWR.n1107 VGND 0.01165f
C42883 VPWR.n1108 VGND 0.00916f
C42884 VPWR.n1109 VGND 0.01042f
C42885 VPWR.n1110 VGND 0.01482f
C42886 VPWR.n1111 VGND 0.01352f
C42887 VPWR.n1112 VGND 0.01013f
C42888 VPWR.n1113 VGND 0.00992f
C42889 VPWR.n1114 VGND 0.00437f
C42890 VPWR.n1115 VGND 0.00988f
C42891 VPWR.n1116 VGND 0.00923f
C42892 VPWR.n1117 VGND 0.00974f
C42893 VPWR.n1118 VGND 0.01085f
C42894 VPWR.n1119 VGND 0.0085f
C42895 VPWR.n1120 VGND 0.008f
C42896 VPWR.n1121 VGND 0.00661f
C42897 VPWR.n1122 VGND 0.01266f
C42898 VPWR.n1123 VGND 0.00788f
C42899 VPWR.n1124 VGND 0.00443f
C42900 VPWR.n1125 VGND 0.00593f
C42901 VPWR.n1126 VGND 0.00545f
C42902 VPWR.n1127 VGND 0.00642f
C42903 VPWR.n1128 VGND 0.00708f
C42904 VPWR.n1129 VGND 0.00708f
C42905 VPWR.n1130 VGND 0.00678f
C42906 VPWR.n1131 VGND 0.00853f
C42907 VPWR.n1132 VGND 0.01129f
C42908 VPWR.n1133 VGND 0.00591f
C42909 VPWR.n1134 VGND 0.0063f
C42910 VPWR.n1135 VGND 0.0056f
C42911 VPWR.n1136 VGND 0.00557f
C42912 VPWR.n1137 VGND 0.0077f
C42913 VPWR.n1138 VGND 0.0077f
C42914 VPWR.n1139 VGND 0.00829f
C42915 VPWR.n1140 VGND 0.00702f
C42916 VPWR.n1141 VGND 0.01165f
C42917 VPWR.n1142 VGND 0.01144f
C42918 VPWR.n1143 VGND 0.0085f
C42919 VPWR.n1144 VGND 0.00974f
C42920 VPWR.n1145 VGND 0.01076f
C42921 VPWR.n1146 VGND 0.00593f
C42922 VPWR.n1147 VGND 0.00501f
C42923 VPWR.n1148 VGND 0.01855f
C42924 VPWR.n1149 VGND 0.02171f
C42925 VPWR.n1150 VGND 0.01588f
C42926 VPWR.n1151 VGND 0.01824f
C42927 VPWR.n1152 VGND 0.01287f
C42928 VPWR.n1153 VGND 0.00653f
C42929 VPWR.n1154 VGND 0.00627f
C42930 VPWR.n1155 VGND 0.00614f
C42931 VPWR.n1156 VGND 0.00546f
C42932 VPWR.n1157 VGND 0.00771f
C42933 VPWR.n1158 VGND 0.13412f
C42934 VPWR.t1080 VGND 0.00473f
C42935 VPWR.n1159 VGND 0.00407f
C42936 VPWR.t903 VGND 0.00473f
C42937 VPWR.t1078 VGND 0.00427f
C42938 VPWR.t4281 VGND 0.00427f
C42939 VPWR.t844 VGND 0.00473f
C42940 VPWR.t5186 VGND 0.00433f
C42941 VPWR.t842 VGND 0.00427f
C42942 VPWR.t7106 VGND 0.00427f
C42943 VPWR.t4480 VGND 0.00473f
C42944 VPWR.t7104 VGND 0.00473f
C42945 VPWR.t4478 VGND 0.00427f
C42946 VPWR.t4484 VGND 0.00427f
C42947 VPWR.t6173 VGND 0.00473f
C42948 VPWR.t4482 VGND 0.00473f
C42949 VPWR.t6175 VGND 0.00427f
C42950 VPWR.t905 VGND 0.00427f
C42951 VPWR.n1160 VGND 0.00698f
C42952 VPWR.n1161 VGND 0.00698f
C42953 VPWR.n1162 VGND 0.00655f
C42954 VPWR.n1163 VGND 0.00655f
C42955 VPWR.n1164 VGND 0.00698f
C42956 VPWR.n1165 VGND 0.00698f
C42957 VPWR.n1166 VGND 0.00655f
C42958 VPWR.n1167 VGND 0.00655f
C42959 VPWR.n1168 VGND 0.00698f
C42960 VPWR.n1169 VGND 0.00819f
C42961 VPWR.n1170 VGND 0.00685f
C42962 VPWR.n1171 VGND 0.00515f
C42963 VPWR.t843 VGND 0.03271f
C42964 VPWR.t5185 VGND 0.02791f
C42965 VPWR.t841 VGND 0.0173f
C42966 VPWR.t7105 VGND 0.01998f
C42967 VPWR.t4479 VGND 0.02791f
C42968 VPWR.t7103 VGND 0.02791f
C42969 VPWR.t4477 VGND 0.01998f
C42970 VPWR.t4483 VGND 0.01998f
C42971 VPWR.t6172 VGND 0.02791f
C42972 VPWR.t4481 VGND 0.02791f
C42973 VPWR.t6174 VGND 0.01998f
C42974 VPWR.t904 VGND 0.01998f
C42975 VPWR.t1079 VGND 0.02791f
C42976 VPWR.t902 VGND 0.02791f
C42977 VPWR.t1077 VGND 0.01998f
C42978 VPWR.n1172 VGND 0.01544f
C42979 VPWR.t3587 VGND 0.00427f
C42980 VPWR.t4279 VGND 0.00473f
C42981 VPWR.t3585 VGND 0.00473f
C42982 VPWR.t5413 VGND 0.00473f
C42983 VPWR.t1866 VGND 0.00473f
C42984 VPWR.t5411 VGND 0.00427f
C42985 VPWR.t1273 VGND 0.00427f
C42986 VPWR.t1868 VGND 0.00427f
C42987 VPWR.t2401 VGND 0.00473f
C42988 VPWR.t1271 VGND 0.00473f
C42989 VPWR.t2399 VGND 0.00427f
C42990 VPWR.t7026 VGND 0.00164f
C42991 VPWR.t1862 VGND 0.00164f
C42992 VPWR.n1173 VGND 0.00331f
C42993 VPWR.t2397 VGND 0.00473f
C42994 VPWR.t2395 VGND 0.00427f
C42995 VPWR.t6244 VGND 0.00473f
C42996 VPWR.t5409 VGND 0.0029f
C42997 VPWR.t2594 VGND 0.00164f
C42998 VPWR.n1174 VGND 0.0047f
C42999 VPWR.t6246 VGND 0.00427f
C43000 VPWR.t2596 VGND 0.00431f
C43001 VPWR.t1689 VGND 0.00473f
C43002 VPWR.t4280 VGND 0.0202f
C43003 VPWR.t3586 VGND 0.01462f
C43004 VPWR.t4278 VGND 0.02791f
C43005 VPWR.t3584 VGND 0.04498f
C43006 VPWR.t5412 VGND 0.03538f
C43007 VPWR.t1865 VGND 0.02791f
C43008 VPWR.t5410 VGND 0.01462f
C43009 VPWR.t1867 VGND 0.0154f
C43010 VPWR.t1272 VGND 0.03003f
C43011 VPWR.t1270 VGND 0.03326f
C43012 VPWR.t2400 VGND 0.03326f
C43013 VPWR.t2398 VGND 0.03963f
C43014 VPWR.t7025 VGND 0.0307f
C43015 VPWR.t1861 VGND 0.02746f
C43016 VPWR.t2396 VGND 0.01652f
C43017 VPWR.t7022 VGND 0.02791f
C43018 VPWR.t2394 VGND 0.02277f
C43019 VPWR.t2592 VGND 0.01172f
C43020 VPWR.t5408 VGND 0.03538f
C43021 VPWR.t6243 VGND 0.02724f
C43022 VPWR.t2593 VGND 0.02791f
C43023 VPWR.t6245 VGND 0.02389f
C43024 VPWR.t2595 VGND 0.01172f
C43025 VPWR.t1316 VGND 0.0173f
C43026 VPWR.t444 VGND 0.02791f
C43027 VPWR.t1314 VGND 0.05001f
C43028 VPWR.t683 VGND 0.03538f
C43029 VPWR.t1318 VGND 0.025f
C43030 VPWR.t1320 VGND 0.04677f
C43031 VPWR.t7012 VGND 0.03538f
C43032 VPWR.t3058 VGND 0.02288f
C43033 VPWR.t4719 VGND 0.02288f
C43034 VPWR.t3060 VGND 0.03293f
C43035 VPWR.t7018 VGND 0.05068f
C43036 VPWR.t4159 VGND 0.02746f
C43037 VPWR.t2123 VGND 0.01652f
C43038 VPWR.t7010 VGND 0.02791f
C43039 VPWR.t2125 VGND 0.02277f
C43040 VPWR.t737 VGND 0.01172f
C43041 VPWR.t1583 VGND 0.01172f
C43042 VPWR.t4155 VGND 0.02724f
C43043 VPWR.t2729 VGND 0.02791f
C43044 VPWR.t4157 VGND 0.02389f
C43045 VPWR.t2727 VGND 0.03248f
C43046 VPWR.t1686 VGND 0.0125f
C43047 VPWR.t1688 VGND 0.0298f
C43048 VPWR.n1175 VGND 0.0266f
C43049 VPWR.t1687 VGND 0.00427f
C43050 VPWR.t2728 VGND 0.00431f
C43051 VPWR.t4158 VGND 0.00473f
C43052 VPWR.t2730 VGND 0.00164f
C43053 VPWR.t1584 VGND 0.0029f
C43054 VPWR.n1176 VGND 0.0047f
C43055 VPWR.t4156 VGND 0.00427f
C43056 VPWR.t2126 VGND 0.00427f
C43057 VPWR.t2124 VGND 0.00473f
C43058 VPWR.t4160 VGND 0.00164f
C43059 VPWR.t7019 VGND 0.00164f
C43060 VPWR.n1177 VGND 0.00331f
C43061 VPWR.t3061 VGND 0.00473f
C43062 VPWR.t4720 VGND 0.00431f
C43063 VPWR.t3059 VGND 0.00427f
C43064 VPWR.t1321 VGND 0.00473f
C43065 VPWR.t684 VGND 0.00433f
C43066 VPWR.n1178 VGND 0.00785f
C43067 VPWR.n1179 VGND 0.00878f
C43068 VPWR.n1180 VGND 0.0076f
C43069 VPWR.n1181 VGND 0.00677f
C43070 VPWR.n1182 VGND 0.00866f
C43071 VPWR.n1183 VGND 0.00679f
C43072 VPWR.n1184 VGND 0.00605f
C43073 VPWR.n1185 VGND 0.00794f
C43074 VPWR.n1186 VGND 0.00887f
C43075 VPWR.n1187 VGND 0.00652f
C43076 VPWR.n1188 VGND 0.00813f
C43077 VPWR.n1189 VGND 0.00721f
C43078 VPWR.n1190 VGND 0.00646f
C43079 VPWR.n1191 VGND 0.01077f
C43080 VPWR.n1192 VGND 0.00543f
C43081 VPWR.n1193 VGND 0.00721f
C43082 VPWR.n1194 VGND 0.00928f
C43083 VPWR.n1195 VGND 0.00538f
C43084 VPWR.n1196 VGND 0.00773f
C43085 VPWR.n1197 VGND 0.00794f
C43086 VPWR.n1198 VGND 0.00605f
C43087 VPWR.n1199 VGND 0.00565f
C43088 VPWR.n1200 VGND 0.01042f
C43089 VPWR.n1201 VGND 0.0054f
C43090 VPWR.n1202 VGND 0.0054f
C43091 VPWR.n1203 VGND 0.0077f
C43092 VPWR.n1204 VGND 0.00708f
C43093 VPWR.n1205 VGND 0.00646f
C43094 VPWR.n1206 VGND 0.00593f
C43095 VPWR.n1207 VGND 0.00577f
C43096 VPWR.n1208 VGND 0.00608f
C43097 VPWR.n1209 VGND 0.00593f
C43098 VPWR.n1210 VGND 0.00708f
C43099 VPWR.n1211 VGND 0.01189f
C43100 VPWR.n1212 VGND 0.00642f
C43101 VPWR.n1213 VGND 0.00698f
C43102 VPWR.n1214 VGND 0.00655f
C43103 VPWR.n1215 VGND 0.00777f
C43104 VPWR.n1216 VGND 0.13412f
C43105 VPWR.t2488 VGND 0.00473f
C43106 VPWR.t4235 VGND 0.00433f
C43107 VPWR.t2486 VGND 0.00427f
C43108 VPWR.t5621 VGND 0.00473f
C43109 VPWR.t2881 VGND 0.00473f
C43110 VPWR.t5623 VGND 0.00427f
C43111 VPWR.t5627 VGND 0.00427f
C43112 VPWR.t2879 VGND 0.00427f
C43113 VPWR.t2184 VGND 0.00427f
C43114 VPWR.t5625 VGND 0.00473f
C43115 VPWR.t1104 VGND 0.00427f
C43116 VPWR.t2182 VGND 0.00473f
C43117 VPWR.t2278 VGND 0.00427f
C43118 VPWR.t1102 VGND 0.00473f
C43119 VPWR.t2276 VGND 0.00473f
C43120 VPWR.n1217 VGND 0.0052f
C43121 VPWR.n1218 VGND 0.00593f
C43122 VPWR.n1219 VGND 0.0076f
C43123 VPWR.n1220 VGND 0.00593f
C43124 VPWR.n1221 VGND 0.00655f
C43125 VPWR.n1222 VGND 0.00593f
C43126 VPWR.n1223 VGND 0.00646f
C43127 VPWR.n1224 VGND 0.00708f
C43128 VPWR.n1225 VGND 0.00708f
C43129 VPWR.n1226 VGND 0.00646f
C43130 VPWR.n1227 VGND 0.00593f
C43131 VPWR.n1228 VGND 0.00577f
C43132 VPWR.t5620 VGND 0.03538f
C43133 VPWR.t2880 VGND 0.02791f
C43134 VPWR.t5622 VGND 0.01462f
C43135 VPWR.t2878 VGND 0.0154f
C43136 VPWR.t5626 VGND 0.0154f
C43137 VPWR.t2183 VGND 0.01462f
C43138 VPWR.t5624 VGND 0.02791f
C43139 VPWR.t2181 VGND 0.03538f
C43140 VPWR.t1103 VGND 0.025f
C43141 VPWR.t2277 VGND 0.01462f
C43142 VPWR.t1101 VGND 0.02791f
C43143 VPWR.t2275 VGND 0.03248f
C43144 VPWR.t2487 VGND 0.03271f
C43145 VPWR.t4234 VGND 0.02712f
C43146 VPWR.t2485 VGND 0.0125f
C43147 VPWR.n1229 VGND 0.02872f
C43148 VPWR.t2428 VGND 0.00433f
C43149 VPWR.t706 VGND 0.00433f
C43150 VPWR.t3889 VGND 0.00473f
C43151 VPWR.t6064 VGND 0.00473f
C43152 VPWR.t3891 VGND 0.00427f
C43153 VPWR.t6062 VGND 0.00427f
C43154 VPWR.t2224 VGND 0.00427f
C43155 VPWR.t6060 VGND 0.00427f
C43156 VPWR.t2226 VGND 0.00473f
C43157 VPWR.t6058 VGND 0.00473f
C43158 VPWR.t4967 VGND 0.00433f
C43159 VPWR.t1070 VGND 0.00427f
C43160 VPWR.t3435 VGND 0.00433f
C43161 VPWR.t1068 VGND 0.00473f
C43162 VPWR.t1235 VGND 0.00433f
C43163 VPWR.t4193 VGND 0.00433f
C43164 VPWR.t5029 VGND 0.00433f
C43165 VPWR.t1876 VGND 0.00433f
C43166 VPWR.t3907 VGND 0.00433f
C43167 VPWR.t2427 VGND 0.03271f
C43168 VPWR.t705 VGND 0.0173f
C43169 VPWR.t3888 VGND 0.03538f
C43170 VPWR.t6063 VGND 0.02791f
C43171 VPWR.t3890 VGND 0.02712f
C43172 VPWR.t6061 VGND 0.0125f
C43173 VPWR.t2223 VGND 0.0125f
C43174 VPWR.t6059 VGND 0.02712f
C43175 VPWR.t2225 VGND 0.02791f
C43176 VPWR.t6057 VGND 0.04789f
C43177 VPWR.t4966 VGND 0.01172f
C43178 VPWR.t1069 VGND 0.03483f
C43179 VPWR.t1067 VGND 0.04309f
C43180 VPWR.t3434 VGND 0.05269f
C43181 VPWR.t1234 VGND 0.05001f
C43182 VPWR.t4192 VGND 0.0173f
C43183 VPWR.t5028 VGND 0.04521f
C43184 VPWR.t1875 VGND 0.0298f
C43185 VPWR.t5738 VGND 0.0202f
C43186 VPWR.t4429 VGND 0.0154f
C43187 VPWR.t4431 VGND 0.0173f
C43188 VPWR.t4334 VGND 0.03538f
C43189 VPWR.t922 VGND 0.04789f
C43190 VPWR.t6633 VGND 0.04231f
C43191 VPWR.t2588 VGND 0.0154f
C43192 VPWR.t5468 VGND 0.025f
C43193 VPWR.t4365 VGND 0.025f
C43194 VPWR.t7017 VGND 0.01395f
C43195 VPWR.t5212 VGND 0.025f
C43196 VPWR.t790 VGND 0.025f
C43197 VPWR.t6087 VGND 0.025f
C43198 VPWR.t1169 VGND 0.025f
C43199 VPWR.t789 VGND 0.02712f
C43200 VPWR.t1873 VGND 0.03605f
C43201 VPWR.t715 VGND 0.025f
C43202 VPWR.t5352 VGND 0.04231f
C43203 VPWR.t934 VGND 0.03271f
C43204 VPWR.t3906 VGND 0.04122f
C43205 VPWR.t935 VGND 0.00433f
C43206 VPWR.t5353 VGND 0.00433f
C43207 VPWR.t716 VGND 0.00433f
C43208 VPWR.t1874 VGND 0.00473f
C43209 VPWR.t1170 VGND 0.00429f
C43210 VPWR.t5213 VGND 0.00498f
C43211 VPWR.t5469 VGND 0.00433f
C43212 VPWR.t2589 VGND 0.00433f
C43213 VPWR.t6634 VGND 0.00433f
C43214 VPWR.t923 VGND 0.00433f
C43215 VPWR.n1230 VGND 0.0084f
C43216 VPWR.n1231 VGND 0.00976f
C43217 VPWR.n1232 VGND 0.0085f
C43218 VPWR.n1233 VGND 0.00825f
C43219 VPWR.n1234 VGND 0.0121f
C43220 VPWR.n1235 VGND 0.00984f
C43221 VPWR.n1236 VGND 0.01118f
C43222 VPWR.n1237 VGND 0.01005f
C43223 VPWR.n1238 VGND 0.00896f
C43224 VPWR.n1239 VGND 0.0058f
C43225 VPWR.n1240 VGND 0.01165f
C43226 VPWR.n1241 VGND 0.01144f
C43227 VPWR.n1242 VGND 0.01085f
C43228 VPWR.n1243 VGND 0.01023f
C43229 VPWR.n1244 VGND 0.00564f
C43230 VPWR.n1245 VGND 0.00791f
C43231 VPWR.n1246 VGND 0.00767f
C43232 VPWR.n1247 VGND 0.00685f
C43233 VPWR.n1248 VGND 0.00943f
C43234 VPWR.n1249 VGND 0.00729f
C43235 VPWR.n1250 VGND 0.00584f
C43236 VPWR.n1251 VGND 0.0054f
C43237 VPWR.n1252 VGND 0.0077f
C43238 VPWR.n1253 VGND 0.00584f
C43239 VPWR.n1254 VGND 0.00584f
C43240 VPWR.n1255 VGND 0.0077f
C43241 VPWR.n1256 VGND 0.0054f
C43242 VPWR.n1257 VGND 0.00819f
C43243 VPWR.n1258 VGND 0.00627f
C43244 VPWR.n1259 VGND 0.00661f
C43245 VPWR.n1260 VGND 0.01093f
C43246 VPWR.n1261 VGND 0.00878f
C43247 VPWR.n1262 VGND 0.00685f
C43248 VPWR.n1263 VGND 0.00432f
C43249 VPWR.n1264 VGND 0.00693f
C43250 VPWR.n1265 VGND 0.13412f
C43251 VPWR.t4382 VGND 0.00427f
C43252 VPWR.t6025 VGND 0.00433f
C43253 VPWR.t4380 VGND 0.00473f
C43254 VPWR.t3278 VGND 0.00427f
C43255 VPWR.t1943 VGND 0.00473f
C43256 VPWR.t3280 VGND 0.00473f
C43257 VPWR.t1941 VGND 0.00427f
C43258 VPWR.t2913 VGND 0.00427f
C43259 VPWR.t2274 VGND 0.00427f
C43260 VPWR.t2912 VGND 0.00473f
C43261 VPWR.t2272 VGND 0.00473f
C43262 VPWR.t5723 VGND 0.00427f
C43263 VPWR.t3711 VGND 0.00427f
C43264 VPWR.t5721 VGND 0.00473f
C43265 VPWR.t3709 VGND 0.00473f
C43266 VPWR.n1266 VGND 0.0056f
C43267 VPWR.n1267 VGND 0.0054f
C43268 VPWR.n1268 VGND 0.0077f
C43269 VPWR.n1269 VGND 0.00557f
C43270 VPWR.n1270 VGND 0.01101f
C43271 VPWR.n1271 VGND 0.01353f
C43272 VPWR.n1272 VGND 0.00698f
C43273 VPWR.n1273 VGND 0.00655f
C43274 VPWR.n1274 VGND 0.00655f
C43275 VPWR.n1275 VGND 0.00745f
C43276 VPWR.t3277 VGND 0.01998f
C43277 VPWR.t1942 VGND 0.02791f
C43278 VPWR.t3279 VGND 0.02791f
C43279 VPWR.t1940 VGND 0.01998f
C43280 VPWR.t2273 VGND 0.03963f
C43281 VPWR.t2271 VGND 0.06039f
C43282 VPWR.t5722 VGND 0.0125f
C43283 VPWR.t3710 VGND 0.02712f
C43284 VPWR.t5720 VGND 0.02791f
C43285 VPWR.t3708 VGND 0.03248f
C43286 VPWR.t4381 VGND 0.0173f
C43287 VPWR.t6024 VGND 0.02288f
C43288 VPWR.t4379 VGND 0.0202f
C43289 VPWR.n1276 VGND 0.0391f
C43290 VPWR.t921 VGND 0.00427f
C43291 VPWR.t4867 VGND 0.00473f
C43292 VPWR.t919 VGND 0.00473f
C43293 VPWR.t4865 VGND 0.00427f
C43294 VPWR.t3098 VGND 0.00473f
C43295 VPWR.t5385 VGND 0.00433f
C43296 VPWR.t3096 VGND 0.00427f
C43297 VPWR.t3151 VGND 0.00427f
C43298 VPWR.t3149 VGND 0.00473f
C43299 VPWR.t1215 VGND 0.00163f
C43300 VPWR.t6872 VGND 0.00163f
C43301 VPWR.n1277 VGND 0.00329f
C43302 VPWR.t901 VGND 0.00433f
C43303 VPWR.t1826 VGND 0.00433f
C43304 VPWR.t2051 VGND 0.00433f
C43305 VPWR.t5059 VGND 0.00429f
C43306 VPWR.t4524 VGND 0.00433f
C43307 VPWR.t920 VGND 0.01998f
C43308 VPWR.t4866 VGND 0.02791f
C43309 VPWR.t918 VGND 0.02791f
C43310 VPWR.t4864 VGND 0.01998f
C43311 VPWR.t3097 VGND 0.03271f
C43312 VPWR.t5384 VGND 0.02791f
C43313 VPWR.t3095 VGND 0.0173f
C43314 VPWR.t3150 VGND 0.01563f
C43315 VPWR.t4282 VGND 0.02668f
C43316 VPWR.t6638 VGND 0.024f
C43317 VPWR.t3148 VGND 0.02277f
C43318 VPWR.t1214 VGND 0.04431f
C43319 VPWR.t6871 VGND 0.02344f
C43320 VPWR.t900 VGND 0.01183f
C43321 VPWR.t4851 VGND 0.0173f
C43322 VPWR.t7011 VGND 0.03271f
C43323 VPWR.t1825 VGND 0.025f
C43324 VPWR.t2507 VGND 0.0298f
C43325 VPWR.t5058 VGND 0.04521f
C43326 VPWR.t2050 VGND 0.03751f
C43327 VPWR.t4523 VGND 0.05372f
C43328 VPWR.t5659 VGND 0.00433f
C43329 VPWR.t3316 VGND 0.00433f
C43330 VPWR.t2902 VGND 0.00433f
C43331 VPWR.t5057 VGND 0.00433f
C43332 VPWR.t353 VGND 0.00433f
C43333 VPWR.t6640 VGND 0.00394f
C43334 VPWR.t6878 VGND 0.00394f
C43335 VPWR.t4094 VGND 0.00425f
C43336 VPWR.t2239 VGND 0.00433f
C43337 VPWR.t6870 VGND 0.00433f
C43338 VPWR.t5476 VGND 0.00498f
C43339 VPWR.t3836 VGND 0.00433f
C43340 VPWR.t3565 VGND 0.00473f
C43341 VPWR.t1957 VGND 0.00473f
C43342 VPWR.t5658 VGND 0.03271f
C43343 VPWR.t3315 VGND 0.05001f
C43344 VPWR.t2901 VGND 0.05001f
C43345 VPWR.t5056 VGND 0.0298f
C43346 VPWR.t352 VGND 0.01183f
C43347 VPWR.t6639 VGND 0.0173f
C43348 VPWR.t6877 VGND 0.03784f
C43349 VPWR.t4093 VGND 0.05079f
C43350 VPWR.t2238 VGND 0.02768f
C43351 VPWR.t788 VGND 0.01172f
C43352 VPWR.t4042 VGND 0.0154f
C43353 VPWR.t6869 VGND 0.0125f
C43354 VPWR.t5475 VGND 0.0154f
C43355 VPWR.t3835 VGND 0.01395f
C43356 VPWR.t2508 VGND 0.02724f
C43357 VPWR.t6037 VGND 0.04565f
C43358 VPWR.t3564 VGND 0.03538f
C43359 VPWR.t1956 VGND 0.03538f
C43360 VPWR.n1278 VGND 0.0295f
C43361 VPWR.t1955 VGND 0.00427f
C43362 VPWR.t3810 VGND 0.00433f
C43363 VPWR.t3508 VGND 0.00427f
C43364 VPWR.t3883 VGND 0.00427f
C43365 VPWR.t3506 VGND 0.00473f
C43366 VPWR.t3879 VGND 0.00473f
C43367 VPWR.t3698 VGND 0.00433f
C43368 VPWR.t3457 VGND 0.00433f
C43369 VPWR.t2522 VGND 0.00433f
C43370 VPWR.t5598 VGND 0.00433f
C43371 VPWR.t3764 VGND 0.00433f
C43372 VPWR.t1150 VGND 0.00433f
C43373 VPWR.t5203 VGND 0.00429f
C43374 VPWR.t1427 VGND 0.00429f
C43375 VPWR.t5201 VGND 0.00164f
C43376 VPWR.t5204 VGND 0.00164f
C43377 VPWR.n1279 VGND 0.0033f
C43378 VPWR.t1431 VGND 0.00164f
C43379 VPWR.t1429 VGND 0.00164f
C43380 VPWR.n1280 VGND 0.0033f
C43381 VPWR.t5202 VGND 0.00429f
C43382 VPWR.t1425 VGND 0.00429f
C43383 VPWR.t4469 VGND 0.00433f
C43384 VPWR.t1954 VGND 0.0173f
C43385 VPWR.t3809 VGND 0.01172f
C43386 VPWR.t3507 VGND 0.0173f
C43387 VPWR.t3505 VGND 0.01172f
C43388 VPWR.t3882 VGND 0.03248f
C43389 VPWR.t3878 VGND 0.025f
C43390 VPWR.t3456 VGND 0.05001f
C43391 VPWR.t2521 VGND 0.08271f
C43392 VPWR.t1149 VGND 0.06731f
C43393 VPWR.t1426 VGND 0.03896f
C43394 VPWR.t1430 VGND 0.05001f
C43395 VPWR.t1428 VGND 0.05001f
C43396 VPWR.t1424 VGND 0.06039f
C43397 VPWR.t4359 VGND 0.02288f
C43398 VPWR.t217 VGND 0.02277f
C43399 VPWR.t225 VGND 0.02277f
C43400 VPWR.t522 VGND 0.02791f
C43401 VPWR.t6618 VGND 0.01172f
C43402 VPWR.t6505 VGND 0.025f
C43403 VPWR.t1958 VGND 0.03538f
C43404 VPWR.t5193 VGND 0.01183f
C43405 VPWR.t1324 VGND 0.0298f
C43406 VPWR.t523 VGND 0.02567f
C43407 VPWR.t114 VGND 0.01395f
C43408 VPWR.t2772 VGND 0.02277f
C43409 VPWR.t2837 VGND 0.03315f
C43410 VPWR.t3679 VGND 0.0173f
C43411 VPWR.t5803 VGND 0.03605f
C43412 VPWR.t5817 VGND 0.0298f
C43413 VPWR.t5442 VGND 0.02277f
C43414 VPWR.t3752 VGND 0.0298f
C43415 VPWR.t4610 VGND 0.03605f
C43416 VPWR.t3677 VGND 0.0298f
C43417 VPWR.t4468 VGND 0.04412f
C43418 VPWR.t3678 VGND 0.00431f
C43419 VPWR.t4611 VGND 0.00433f
C43420 VPWR.t3753 VGND 0.00394f
C43421 VPWR.t5443 VGND 0.00433f
C43422 VPWR.t5818 VGND 0.00394f
C43423 VPWR.t5804 VGND 0.00433f
C43424 VPWR.t3680 VGND 0.00431f
C43425 VPWR.t2838 VGND 0.00394f
C43426 VPWR.t2773 VGND 0.00431f
C43427 VPWR.t115 VGND 0.00394f
C43428 VPWR.t524 VGND 0.00394f
C43429 VPWR.t5194 VGND 0.00433f
C43430 VPWR.t1325 VGND 0.00394f
C43431 VPWR.t1959 VGND 0.00498f
C43432 VPWR.n1281 VGND 0.00975f
C43433 VPWR.n1282 VGND 0.00665f
C43434 VPWR.n1283 VGND 0.00651f
C43435 VPWR.n1284 VGND 0.00691f
C43436 VPWR.n1285 VGND 0.00645f
C43437 VPWR.n1286 VGND 0.00608f
C43438 VPWR.n1287 VGND 0.00783f
C43439 VPWR.n1288 VGND 0.0067f
C43440 VPWR.n1289 VGND 0.00823f
C43441 VPWR.n1290 VGND 0.00902f
C43442 VPWR.n1291 VGND 0.00651f
C43443 VPWR.n1292 VGND 0.009f
C43444 VPWR.n1293 VGND 0.00596f
C43445 VPWR.n1294 VGND 0.00842f
C43446 VPWR.n1295 VGND 0.0122f
C43447 VPWR.n1296 VGND 0.00647f
C43448 VPWR.n1297 VGND 0.01684f
C43449 VPWR.n1298 VGND 0.00986f
C43450 VPWR.n1299 VGND 0.02118f
C43451 VPWR.n1300 VGND 0.01588f
C43452 VPWR.n1301 VGND 0.01824f
C43453 VPWR.n1302 VGND 0.01287f
C43454 VPWR.n1303 VGND 0.0052f
C43455 VPWR.n1304 VGND 0.00655f
C43456 VPWR.n1305 VGND 0.00655f
C43457 VPWR.n1306 VGND 0.00596f
C43458 VPWR.n1307 VGND 0.00614f
C43459 VPWR.n1308 VGND 0.00646f
C43460 VPWR.n1309 VGND 0.01139f
C43461 VPWR.n1310 VGND 0.00601f
C43462 VPWR.n1311 VGND 0.00623f
C43463 VPWR.n1312 VGND 0.00845f
C43464 VPWR.n1313 VGND 0.00912f
C43465 VPWR.n1314 VGND 0.00775f
C43466 VPWR.n1315 VGND 0.00914f
C43467 VPWR.n1316 VGND 0.0074f
C43468 VPWR.n1317 VGND 0.00732f
C43469 VPWR.n1318 VGND 0.00727f
C43470 VPWR.n1319 VGND 0.00876f
C43471 VPWR.n1320 VGND 0.01087f
C43472 VPWR.n1321 VGND 0.01023f
C43473 VPWR.n1322 VGND 0.00564f
C43474 VPWR.n1323 VGND 0.00974f
C43475 VPWR.n1324 VGND 0.00661f
C43476 VPWR.n1325 VGND 0.01266f
C43477 VPWR.n1326 VGND 0.0072f
C43478 VPWR.n1327 VGND 0.00981f
C43479 VPWR.n1328 VGND 0.00616f
C43480 VPWR.n1329 VGND 0.01172f
C43481 VPWR.n1330 VGND 0.00896f
C43482 VPWR.n1331 VGND 0.00448f
C43483 VPWR.n1332 VGND 0.00839f
C43484 VPWR.n1333 VGND 0.00993f
C43485 VPWR.n1334 VGND 0.00819f
C43486 VPWR.n1335 VGND 0.00685f
C43487 VPWR.n1336 VGND 0.00515f
C43488 VPWR.n1337 VGND 0.00776f
C43489 VPWR.n1338 VGND 0.00655f
C43490 VPWR.n1339 VGND 0.00655f
C43491 VPWR.n1340 VGND 0.0076f
C43492 VPWR.n1341 VGND 0.01189f
C43493 VPWR.n1342 VGND 0.0059f
C43494 VPWR.n1343 VGND 0.01173f
C43495 VPWR.n1344 VGND 0.00679f
C43496 VPWR.n1345 VGND 0.13412f
C43497 VPWR.n1346 VGND 0.20174f
C43498 VPWR.n1347 VGND 0.00777f
C43499 VPWR.n1348 VGND 0.00542f
C43500 VPWR.n1349 VGND 0.0068f
C43501 VPWR.n1350 VGND 0.0117f
C43502 VPWR.n1351 VGND 0.00471f
C43503 VPWR.n1352 VGND 0.00813f
C43504 VPWR.n1353 VGND 0.00471f
C43505 VPWR.n1354 VGND 0.00712f
C43506 VPWR.n1355 VGND 0.00596f
C43507 VPWR.n1356 VGND 0.01114f
C43508 VPWR.n1357 VGND 0.00943f
C43509 VPWR.n1358 VGND 0.00306f
C43510 VPWR.n1359 VGND 0.01189f
C43511 VPWR.n1360 VGND 0.00863f
C43512 VPWR.n1361 VGND 0.00415f
C43513 VPWR.n1362 VGND 0.00773f
C43514 VPWR.n1363 VGND 0.00576f
C43515 VPWR.n1364 VGND 0.00875f
C43516 VPWR.n1365 VGND 0.00847f
C43517 VPWR.n1366 VGND 0.01089f
C43518 VPWR.t6632 VGND 0.00187f
C43519 VPWR.t6082 VGND 0.00139f
C43520 VPWR.n1367 VGND 0.00471f
C43521 VPWR.t5209 VGND 0.00187f
C43522 VPWR.t5123 VGND 0.00139f
C43523 VPWR.n1368 VGND 0.00471f
C43524 VPWR.t6271 VGND 0.00159f
C43525 VPWR.t971 VGND 0.00158f
C43526 VPWR.n1369 VGND 0.00497f
C43527 VPWR.t1910 VGND 0.00516f
C43528 VPWR.n1370 VGND 0.00145f
C43529 VPWR.t3834 VGND 0.00196f
C43530 VPWR.t5 VGND 0.00157f
C43531 VPWR.n1371 VGND 0.00539f
C43532 VPWR.t315 VGND 0.00132f
C43533 VPWR.t3755 VGND 0.00132f
C43534 VPWR.n1372 VGND 0.00266f
C43535 VPWR.t7015 VGND 0.00433f
C43536 VPWR.t1129 VGND 0.00394f
C43537 VPWR.t4076 VGND 0.00516f
C43538 VPWR.t5211 VGND 0.00394f
C43539 VPWR.n1373 VGND 0.00711f
C43540 VPWR.n1374 VGND 0.00589f
C43541 VPWR.n1375 VGND 0.00702f
C43542 VPWR.n1376 VGND 0.01098f
C43543 VPWR.n1377 VGND 0.00768f
C43544 VPWR.n1378 VGND 0.00535f
C43545 VPWR.n1379 VGND 0.00684f
C43546 VPWR.n1380 VGND 0.00994f
C43547 VPWR.n1381 VGND 0.01042f
C43548 VPWR.n1382 VGND 0.00573f
C43549 VPWR.n1383 VGND 0.00537f
C43550 VPWR.n1384 VGND 0.01077f
C43551 VPWR.n1385 VGND 0.02649f
C43552 VPWR.t6631 VGND 0.0173f
C43553 VPWR.t6081 VGND 0.025f
C43554 VPWR.t2237 VGND 0.0125f
C43555 VPWR.t1130 VGND 0.02422f
C43556 VPWR.t897 VGND 0.02277f
C43557 VPWR.t5208 VGND 0.02902f
C43558 VPWR.t6270 VGND 0.03036f
C43559 VPWR.t5122 VGND 0.02902f
C43560 VPWR.t970 VGND 0.0317f
C43561 VPWR.t6793 VGND 0.0125f
C43562 VPWR.t1909 VGND 0.02199f
C43563 VPWR.t7094 VGND 0.02277f
C43564 VPWR.t6178 VGND 0.02277f
C43565 VPWR.t3833 VGND 0.02724f
C43566 VPWR.t314 VGND 0.03259f
C43567 VPWR.t4 VGND 0.02277f
C43568 VPWR.t3754 VGND 0.03516f
C43569 VPWR.t7014 VGND 0.025f
C43570 VPWR.t1128 VGND 0.03605f
C43571 VPWR.t5210 VGND 0.025f
C43572 VPWR.t4075 VGND 0.0154f
C43573 VPWR.t323 VGND 0.03896f
C43574 VPWR.t5270 VGND 0.04309f
C43575 VPWR.n1386 VGND 0.03687f
C43576 VPWR.t2153 VGND 0.00427f
C43577 VPWR.t5269 VGND 0.00163f
C43578 VPWR.t5810 VGND 0.00163f
C43579 VPWR.n1387 VGND 0.00328f
C43580 VPWR.t2151 VGND 0.00473f
C43581 VPWR.t4273 VGND 0.00433f
C43582 VPWR.t2658 VGND 0.00429f
C43583 VPWR.t5816 VGND 0.00431f
C43584 VPWR.t2653 VGND 0.00164f
C43585 VPWR.t2660 VGND 0.00164f
C43586 VPWR.n1388 VGND 0.0033f
C43587 VPWR.t5268 VGND 0.01172f
C43588 VPWR.t2152 VGND 0.02277f
C43589 VPWR.t5809 VGND 0.02791f
C43590 VPWR.t2150 VGND 0.025f
C43591 VPWR.t7064 VGND 0.03248f
C43592 VPWR.t5895 VGND 0.02579f
C43593 VPWR.t322 VGND 0.03192f
C43594 VPWR.t4272 VGND 0.02422f
C43595 VPWR.t2657 VGND 0.0154f
C43596 VPWR.t5815 VGND 0.02288f
C43597 VPWR.t2652 VGND 0.0317f
C43598 VPWR.t2659 VGND 0.03192f
C43599 VPWR.n1389 VGND 0.03017f
C43600 VPWR.t2656 VGND 0.00429f
C43601 VPWR.t4603 VGND 0.00429f
C43602 VPWR.t6281 VGND 0.00429f
C43603 VPWR.t4599 VGND 0.00164f
C43604 VPWR.t4605 VGND 0.00164f
C43605 VPWR.n1390 VGND 0.0033f
C43606 VPWR.t6277 VGND 0.00164f
C43607 VPWR.t6275 VGND 0.00164f
C43608 VPWR.n1391 VGND 0.0033f
C43609 VPWR.t4601 VGND 0.00429f
C43610 VPWR.t6279 VGND 0.00429f
C43611 VPWR.t6734 VGND 0.00203f
C43612 VPWR.t2655 VGND 0.0125f
C43613 VPWR.t4602 VGND 0.03605f
C43614 VPWR.t6280 VGND 0.02724f
C43615 VPWR.t4598 VGND 0.02724f
C43616 VPWR.t6276 VGND 0.02277f
C43617 VPWR.t4604 VGND 0.02277f
C43618 VPWR.t6274 VGND 0.02724f
C43619 VPWR.t4600 VGND 0.02645f
C43620 VPWR.t6278 VGND 0.0125f
C43621 VPWR.t6733 VGND 0.0173f
C43622 VPWR.n1392 VGND 0.02649f
C43623 VPWR.t5040 VGND 0.00429f
C43624 VPWR.n1393 VGND 0.00162f
C43625 VPWR.t3751 VGND 0.00149f
C43626 VPWR.t5585 VGND 0.00281f
C43627 VPWR.n1394 VGND 0.00388f
C43628 VPWR.t6737 VGND 0.00454f
C43629 VPWR.t3490 VGND 0.00431f
C43630 VPWR.t6761 VGND 0.00431f
C43631 VPWR.t1035 VGND 0.00163f
C43632 VPWR.t2609 VGND 0.00163f
C43633 VPWR.n1395 VGND 0.00329f
C43634 VPWR.t2769 VGND 0.00431f
C43635 VPWR.t6751 VGND 0.00116f
C43636 VPWR.t6948 VGND 0.00116f
C43637 VPWR.n1396 VGND 0.00236f
C43638 VPWR.t2336 VGND 0.00255f
C43639 VPWR.t7062 VGND 0.0202f
C43640 VPWR.t5039 VGND 0.0211f
C43641 VPWR.t6216 VGND 0.02724f
C43642 VPWR.t5896 VGND 0.02277f
C43643 VPWR.t3750 VGND 0.02277f
C43644 VPWR.t2654 VGND 0.02902f
C43645 VPWR.t5584 VGND 0.02724f
C43646 VPWR.t7066 VGND 0.03885f
C43647 VPWR.t6736 VGND 0.03282f
C43648 VPWR.t6738 VGND 0.03617f
C43649 VPWR.t6760 VGND 0.02824f
C43650 VPWR.t3489 VGND 0.02712f
C43651 VPWR.t7065 VGND 0.02668f
C43652 VPWR.t2573 VGND 0.025f
C43653 VPWR.t6735 VGND 0.02277f
C43654 VPWR.t203 VGND 0.02445f
C43655 VPWR.t1034 VGND 0.03371f
C43656 VPWR.t2608 VGND 0.025f
C43657 VPWR.t2768 VGND 0.01395f
C43658 VPWR.t6750 VGND 0.025f
C43659 VPWR.t6947 VGND 0.02389f
C43660 VPWR.t205 VGND 0.03538f
C43661 VPWR.t2335 VGND 0.025f
C43662 VPWR.t4911 VGND 0.01775f
C43663 VPWR.n1397 VGND 0.02234f
C43664 VPWR.t4256 VGND 0.00433f
C43665 VPWR.n1398 VGND 0.00115f
C43666 VPWR.t6723 VGND 0.00433f
C43667 VPWR.t6027 VGND 0.00394f
C43668 VPWR.t5050 VGND 0.00107f
C43669 VPWR.n1399 VGND 0.00292f
C43670 VPWR.t3181 VGND 0.00394f
C43671 VPWR.t2440 VGND 0.00427f
C43672 VPWR.t2681 VGND 0.00429f
C43673 VPWR.t2438 VGND 0.00603f
C43674 VPWR.t6946 VGND 0.01909f
C43675 VPWR.t879 VGND 0.03014f
C43676 VPWR.t4255 VGND 0.02411f
C43677 VPWR.t4247 VGND 0.0173f
C43678 VPWR.t6945 VGND 0.01172f
C43679 VPWR.t6722 VGND 0.03181f
C43680 VPWR.t2337 VGND 0.03829f
C43681 VPWR.t2435 VGND 0.01183f
C43682 VPWR.t6026 VGND 0.02422f
C43683 VPWR.t3180 VGND 0.02623f
C43684 VPWR.t5049 VGND 0.04231f
C43685 VPWR.t2439 VGND 0.04945f
C43686 VPWR.t2680 VGND 0.02277f
C43687 VPWR.t2437 VGND 0.025f
C43688 VPWR.t4316 VGND 0.03784f
C43689 VPWR.t3179 VGND 0.0298f
C43690 VPWR.n1400 VGND 0.02649f
C43691 VPWR.t6759 VGND 0.00116f
C43692 VPWR.t7061 VGND 0.00116f
C43693 VPWR.n1401 VGND 0.00236f
C43694 VPWR.t22 VGND 0.00394f
C43695 VPWR.t2159 VGND 0.00255f
C43696 VPWR.t1055 VGND 0.00394f
C43697 VPWR.t3157 VGND 0.01733f
C43698 VPWR.t1881 VGND 0.0202f
C43699 VPWR.t6758 VGND 0.0125f
C43700 VPWR.t7060 VGND 0.025f
C43701 VPWR.t21 VGND 0.03784f
C43702 VPWR.t2158 VGND 0.02277f
C43703 VPWR.t1054 VGND 0.03711f
C43704 VPWR.n1403 VGND 0.01237f
C43705 VPWR.t5084 VGND 0.01733f
C43706 VPWR.t6694 VGND 0.0202f
C43707 VPWR.t6704 VGND 0.01395f
C43708 VPWR.t6492 VGND 0.02724f
C43709 VPWR.t6700 VGND 0.02277f
C43710 VPWR.t7041 VGND 0.02277f
C43711 VPWR.t6698 VGND 0.04822f
C43712 VPWR.t805 VGND 0.02724f
C43713 VPWR.t6702 VGND 0.01217f
C43714 VPWR.n1405 VGND 0.01275f
C43715 VPWR.t3124 VGND 0.02973f
C43716 VPWR.t7040 VGND 0.02389f
C43717 VPWR.t1478 VGND 0.02534f
C43718 VPWR.t5085 VGND 0.04521f
C43719 VPWR.t835 VGND 0.03338f
C43720 VPWR.t7043 VGND 0.03527f
C43721 VPWR.t804 VGND 0.03538f
C43722 VPWR.t2161 VGND 0.01741f
C43723 VPWR.t4448 VGND 0.02768f
C43724 VPWR.t837 VGND 0.02768f
C43725 VPWR.t5479 VGND 0.01741f
C43726 VPWR.t2160 VGND 0.03538f
C43727 VPWR.t7059 VGND 0.03527f
C43728 VPWR.t4450 VGND 0.03338f
C43729 VPWR.t3158 VGND 0.03561f
C43730 VPWR.t5257 VGND 0.025f
C43731 VPWR.t7058 VGND 0.0173f
C43732 VPWR.n1406 VGND 0.01198f
C43733 VPWR.n1407 VGND 0.00115f
C43734 VPWR.t4451 VGND 0.00427f
C43735 VPWR.t5480 VGND 0.00107f
C43736 VPWR.n1408 VGND 0.00292f
C43737 VPWR.t2162 VGND 0.00107f
C43738 VPWR.n1409 VGND 0.00292f
C43739 VPWR.t836 VGND 0.00427f
C43740 VPWR.n1410 VGND 0.00115f
C43741 VPWR.t3125 VGND 0.00433f
C43742 VPWR.t6703 VGND 0.00296f
C43743 VPWR.t806 VGND 0.00255f
C43744 VPWR.t6699 VGND 0.0011f
C43745 VPWR.t6701 VGND 0.0011f
C43746 VPWR.n1411 VGND 0.00223f
C43747 VPWR.t7042 VGND 0.00116f
C43748 VPWR.t6493 VGND 0.00116f
C43749 VPWR.n1412 VGND 0.00236f
C43750 VPWR.n1413 VGND 0.00561f
C43751 VPWR.n1414 VGND 0.00734f
C43752 VPWR.n1415 VGND 0.01013f
C43753 VPWR.n1416 VGND 0.01019f
C43754 VPWR.n1417 VGND 0.00896f
C43755 VPWR.n1418 VGND 0.01051f
C43756 VPWR.n1419 VGND 0.01633f
C43757 VPWR.n1420 VGND 0.01026f
C43758 VPWR.n1421 VGND 0.01026f
C43759 VPWR.n1422 VGND 0.01605f
C43760 VPWR.n1423 VGND 0.00591f
C43761 VPWR.n1424 VGND 0.01165f
C43762 VPWR.n1425 VGND 0.00984f
C43763 VPWR.n1426 VGND 0.0063f
C43764 VPWR.n1427 VGND 0.0073f
C43765 VPWR.n1428 VGND 0.00513f
C43766 VPWR.n1429 VGND 0.0099f
C43767 VPWR.n1430 VGND 0.0143f
C43768 VPWR.n1431 VGND 0.01096f
C43769 VPWR.n1432 VGND 0.0078f
C43770 VPWR.n1433 VGND 0.00919f
C43771 VPWR.n1434 VGND 0.00538f
C43772 VPWR.n1435 VGND 0.01074f
C43773 VPWR.n1436 VGND 0.01174f
C43774 VPWR.n1437 VGND 0.00552f
C43775 VPWR.n1438 VGND 0.00811f
C43776 VPWR.n1439 VGND 0.03918f
C43777 VPWR.n1440 VGND 0.00757f
C43778 VPWR.n1441 VGND 0.00928f
C43779 VPWR.n1442 VGND 0.00325f
C43780 VPWR.n1443 VGND 0.00975f
C43781 VPWR.n1444 VGND 0.00917f
C43782 VPWR.n1445 VGND 0.00935f
C43783 VPWR.n1446 VGND 0.00792f
C43784 VPWR.n1447 VGND 0.01069f
C43785 VPWR.n1448 VGND 0.00917f
C43786 VPWR.n1449 VGND 0.00948f
C43787 VPWR.n1450 VGND 0.00699f
C43788 VPWR.n1451 VGND 0.0099f
C43789 VPWR.n1452 VGND 0.0047f
C43790 VPWR.n1453 VGND 0.00607f
C43791 VPWR.n1454 VGND 0.01059f
C43792 VPWR.n1455 VGND 0.00698f
C43793 VPWR.n1456 VGND 0.00288f
C43794 VPWR.n1457 VGND 0.00996f
C43795 VPWR.n1458 VGND 0.00711f
C43796 VPWR.n1459 VGND 0.00686f
C43797 VPWR.n1460 VGND 0.01165f
C43798 VPWR.n1461 VGND 0.00459f
C43799 VPWR.n1462 VGND 0.00842f
C43800 VPWR.n1463 VGND 0.00664f
C43801 VPWR.n1464 VGND 0.00823f
C43802 VPWR.n1465 VGND 0.00855f
C43803 VPWR.n1466 VGND 0.00368f
C43804 VPWR.n1467 VGND 0.00706f
C43805 VPWR.n1468 VGND 0.01165f
C43806 VPWR.n1469 VGND 0.00677f
C43807 VPWR.n1470 VGND 0.00718f
C43808 VPWR.n1471 VGND 0.20174f
C43809 VPWR.n1472 VGND 0.0272f
C43810 VPWR.n1473 VGND 0.00207f
C43811 VPWR.n1474 VGND 0.01266f
C43812 VPWR.n1475 VGND 0.01093f
C43813 VPWR.n1476 VGND 0.00896f
C43814 VPWR.n1477 VGND 0.01174f
C43815 VPWR.n1478 VGND 0.01501f
C43816 VPWR.n1479 VGND 0.01147f
C43817 VPWR.n1480 VGND 0.01202f
C43818 VPWR.n1481 VGND 0.01115f
C43819 VPWR.n1482 VGND 0.01189f
C43820 VPWR.n1483 VGND 0.01001f
C43821 VPWR.n1484 VGND 0.0268f
C43822 VPWR.n1485 VGND 0.01771f
C43823 VPWR.n1486 VGND 0.00919f
C43824 VPWR.n1487 VGND 0.00452f
C43825 VPWR.n1488 VGND 0.01775f
C43826 VPWR.n1489 VGND 0.01189f
C43827 VPWR.n1490 VGND 0.01371f
C43828 VPWR.n1491 VGND 0.0178f
C43829 VPWR.n1492 VGND 0.0178f
C43830 VPWR.n1493 VGND 0.01679f
C43831 VPWR.n1494 VGND 0.01186f
C43832 VPWR.n1495 VGND 0.0178f
C43833 VPWR.n1496 VGND 0.0178f
C43834 VPWR.n1497 VGND 0.01839f
C43835 VPWR.t7128 VGND 0.00433f
C43836 VPWR.t623 VGND 0.00433f
C43837 VPWR.t4284 VGND 0.00433f
C43838 VPWR.t3282 VGND 0.00433f
C43839 VPWR.t5981 VGND 0.00433f
C43840 VPWR.t5918 VGND 0.00433f
C43841 VPWR.t720 VGND 0.00433f
C43842 VPWR.t5495 VGND 0.00433f
C43843 VPWR.n1498 VGND 0.01634f
C43844 VPWR.n1499 VGND 0.0178f
C43845 VPWR.n1500 VGND 0.0178f
C43846 VPWR.n1501 VGND 0.01186f
C43847 VPWR.n1502 VGND 0.01679f
C43848 VPWR.n1503 VGND 0.0178f
C43849 VPWR.n1504 VGND 0.0178f
C43850 VPWR.n1505 VGND 0.01371f
C43851 VPWR.n1506 VGND 0.01189f
C43852 VPWR.n1507 VGND 0.03832f
C43853 VPWR.t7127 VGND 0.05247f
C43854 VPWR.t622 VGND 0.05996f
C43855 VPWR.t4283 VGND 0.05996f
C43856 VPWR.t3281 VGND 0.05996f
C43857 VPWR.t5980 VGND 0.05996f
C43858 VPWR.t5917 VGND 0.05996f
C43859 VPWR.t719 VGND 0.05996f
C43860 VPWR.t5494 VGND 0.04035f
C43861 VPWR.t6516 VGND 0.02998f
C43862 VPWR.t6524 VGND 0.02998f
C43863 VPWR.t3662 VGND 0.02998f
C43864 VPWR.t3664 VGND 0.02998f
C43865 VPWR.t6514 VGND 0.02998f
C43866 VPWR.t6521 VGND 0.02998f
C43867 VPWR.t3666 VGND 0.02202f
C43868 VPWR.t4314 VGND 0.02255f
C43869 VPWR.t4677 VGND 0.03105f
C43870 VPWR.t6227 VGND 0.03172f
C43871 VPWR.t4679 VGND 0.03403f
C43872 VPWR.t4312 VGND 0.04225f
C43873 VPWR.n1508 VGND 0.0262f
C43874 VPWR.n1509 VGND 0.01165f
C43875 VPWR.n1510 VGND 0.01813f
C43876 VPWR.n1511 VGND 0.02074f
C43877 VPWR.n1512 VGND 0.01007f
C43878 VPWR.n1513 VGND 0.021f
C43879 VPWR.n1514 VGND 0.0171f
C43880 VPWR.n1515 VGND 0.02178f
C43881 VPWR.t5932 VGND 0.00431f
C43882 VPWR.t5928 VGND 0.00431f
C43883 VPWR.t3560 VGND 0.00431f
C43884 VPWR.t2761 VGND 0.00433f
C43885 VPWR.t1164 VGND 0.00433f
C43886 VPWR.n1516 VGND 0.01256f
C43887 VPWR.n1517 VGND 0.01197f
C43888 VPWR.n1518 VGND 0.01015f
C43889 VPWR.n1519 VGND 0.01015f
C43890 VPWR.n1520 VGND 0.01015f
C43891 VPWR.n1521 VGND 0.01165f
C43892 VPWR.n1522 VGND 0.03992f
C43893 VPWR.t2360 VGND 0.03795f
C43894 VPWR.t5931 VGND 0.02269f
C43895 VPWR.t5927 VGND 0.02269f
C43896 VPWR.t6621 VGND 0.03621f
C43897 VPWR.t6771 VGND 0.03795f
C43898 VPWR.t3559 VGND 0.02269f
C43899 VPWR.t2760 VGND 0.04959f
C43900 VPWR.t1163 VGND 0.04035f
C43901 VPWR.n1523 VGND 0.0262f
C43902 VPWR.t1206 VGND 0.03661f
C43903 VPWR.t6785 VGND 0.02998f
C43904 VPWR.t6786 VGND 0.02998f
C43905 VPWR.t1204 VGND 0.02998f
C43906 VPWR.t1202 VGND 0.02998f
C43907 VPWR.t6781 VGND 0.02998f
C43908 VPWR.t6782 VGND 0.02998f
C43909 VPWR.t1200 VGND 0.02202f
C43910 VPWR.t45 VGND 0.02068f
C43911 VPWR.t2356 VGND 0.03025f
C43912 VPWR.t7107 VGND 0.03754f
C43913 VPWR.t2287 VGND 0.02998f
C43914 VPWR.n1524 VGND 0.02794f
C43915 VPWR.t109 VGND 0.00431f
C43916 VPWR.t1233 VGND 0.00433f
C43917 VPWR.t6579 VGND 0.00394f
C43918 VPWR.t6628 VGND 0.00394f
C43919 VPWR.t5832 VGND 0.00431f
C43920 VPWR.t5387 VGND 0.00433f
C43921 VPWR.t2581 VGND 0.00433f
C43922 VPWR.t108 VGND 0.02269f
C43923 VPWR.t6972 VGND 0.03621f
C43924 VPWR.t1232 VGND 0.02998f
C43925 VPWR.t6578 VGND 0.02075f
C43926 VPWR.t6627 VGND 0.04343f
C43927 VPWR.t6622 VGND 0.04544f
C43928 VPWR.t5831 VGND 0.02269f
C43929 VPWR.t5386 VGND 0.02998f
C43930 VPWR.t2580 VGND 0.03286f
C43931 VPWR.n1525 VGND 0.0507f
C43932 VPWR.t779 VGND 0.00433f
C43933 VPWR.t2585 VGND 0.00433f
C43934 VPWR.t4154 VGND 0.00433f
C43935 VPWR.t2307 VGND 0.00433f
C43936 VPWR.t6200 VGND 0.00433f
C43937 VPWR.t1660 VGND 0.00433f
C43938 VPWR.t2149 VGND 0.00433f
C43939 VPWR.t778 VGND 0.03286f
C43940 VPWR.t2584 VGND 0.04959f
C43941 VPWR.t4153 VGND 0.04035f
C43942 VPWR.t2306 VGND 0.02824f
C43943 VPWR.t6199 VGND 0.04959f
C43944 VPWR.t1659 VGND 0.04035f
C43945 VPWR.t2148 VGND 0.02824f
C43946 VPWR.n1526 VGND 0.0262f
C43947 VPWR.t5318 VGND 0.00433f
C43948 VPWR.t546 VGND 0.00433f
C43949 VPWR.t5351 VGND 0.00433f
C43950 VPWR.t848 VGND 0.00433f
C43951 VPWR.t1313 VGND 0.00433f
C43952 VPWR.t6898 VGND 0.00394f
C43953 VPWR.t6904 VGND 0.00394f
C43954 VPWR.t6673 VGND 0.00431f
C43955 VPWR.t5317 VGND 0.02998f
C43956 VPWR.t545 VGND 0.04959f
C43957 VPWR.t5350 VGND 0.05996f
C43958 VPWR.t847 VGND 0.05996f
C43959 VPWR.t1312 VGND 0.04035f
C43960 VPWR.t6897 VGND 0.03038f
C43961 VPWR.t6903 VGND 0.02075f
C43962 VPWR.t6672 VGND 0.02269f
C43963 VPWR.t6899 VGND 0.04082f
C43964 VPWR.t2318 VGND 0.00433f
C43965 VPWR.t2591 VGND 0.00433f
C43966 VPWR.t1904 VGND 0.00433f
C43967 VPWR.t3108 VGND 0.00433f
C43968 VPWR.t2294 VGND 0.00433f
C43969 VPWR.t2082 VGND 0.00433f
C43970 VPWR.t4581 VGND 0.00433f
C43971 VPWR.n1527 VGND 0.00732f
C43972 VPWR.n1528 VGND 0.01544f
C43973 VPWR.n1529 VGND 0.01668f
C43974 VPWR.n1530 VGND 0.01197f
C43975 VPWR.n1531 VGND 0.01811f
C43976 VPWR.n1532 VGND 0.01355f
C43977 VPWR.n1533 VGND 0.00896f
C43978 VPWR.t5304 VGND 0.00433f
C43979 VPWR.t1841 VGND 0.00433f
C43980 VPWR.t544 VGND 0.00433f
C43981 VPWR.t5873 VGND 0.00433f
C43982 VPWR.t2446 VGND 0.00433f
C43983 VPWR.t1408 VGND 0.00433f
C43984 VPWR.t4124 VGND 0.00433f
C43985 VPWR.t5303 VGND 0.02824f
C43986 VPWR.t1840 VGND 0.04959f
C43987 VPWR.t543 VGND 0.04035f
C43988 VPWR.t5872 VGND 0.02824f
C43989 VPWR.t2445 VGND 0.04959f
C43990 VPWR.t1407 VGND 0.04035f
C43991 VPWR.t4123 VGND 0.02824f
C43992 VPWR.n1534 VGND 0.0337f
C43993 VPWR.t2629 VGND 0.00433f
C43994 VPWR.t1382 VGND 0.00435f
C43995 VPWR.t3941 VGND 0.00433f
C43996 VPWR.t1132 VGND 0.00433f
C43997 VPWR.t321 VGND 0.00435f
C43998 VPWR.t2759 VGND 0.00433f
C43999 VPWR.t1221 VGND 0.00435f
C44000 VPWR.t2628 VGND 0.02998f
C44001 VPWR.t1381 VGND 0.02824f
C44002 VPWR.t3940 VGND 0.04959f
C44003 VPWR.t1131 VGND 0.04035f
C44004 VPWR.t320 VGND 0.02824f
C44005 VPWR.t2758 VGND 0.02998f
C44006 VPWR.t1220 VGND 0.03286f
C44007 VPWR.n1535 VGND 0.03985f
C44008 VPWR.t1705 VGND 0.00433f
C44009 VPWR.t1029 VGND 0.00433f
C44010 VPWR.t2292 VGND 0.00435f
C44011 VPWR.t4343 VGND 0.00433f
C44012 VPWR.t3766 VGND 0.00433f
C44013 VPWR.t859 VGND 0.00433f
C44014 VPWR.t5635 VGND 0.00433f
C44015 VPWR.t1704 VGND 0.04959f
C44016 VPWR.t1028 VGND 0.04035f
C44017 VPWR.t2291 VGND 0.02824f
C44018 VPWR.t4342 VGND 0.04959f
C44019 VPWR.t3765 VGND 0.05996f
C44020 VPWR.t858 VGND 0.05996f
C44021 VPWR.t5634 VGND 0.04035f
C44022 VPWR.t4243 VGND 0.00433f
C44023 VPWR.t2835 VGND 0.00433f
C44024 VPWR.t654 VGND 0.00433f
C44025 VPWR.t4893 VGND 0.00433f
C44026 VPWR.t2290 VGND 0.00433f
C44027 VPWR.t351 VGND 0.00433f
C44028 VPWR.n1536 VGND 0.01743f
C44029 VPWR.n1537 VGND 0.01679f
C44030 VPWR.n1538 VGND 0.01186f
C44031 VPWR.n1539 VGND 0.0178f
C44032 VPWR.n1540 VGND 0.0178f
C44033 VPWR.n1541 VGND 0.01842f
C44034 VPWR.t4242 VGND 0.04035f
C44035 VPWR.t2834 VGND 0.05996f
C44036 VPWR.t653 VGND 0.05996f
C44037 VPWR.t4892 VGND 0.05996f
C44038 VPWR.t2289 VGND 0.05996f
C44039 VPWR.t350 VGND 0.05996f
C44040 VPWR.t5400 VGND 0.05996f
C44041 VPWR.t6116 VGND 0.05247f
C44042 VPWR.n1542 VGND 0.03832f
C44043 VPWR.t6117 VGND 0.00433f
C44044 VPWR.t5401 VGND 0.00433f
C44045 VPWR.n1543 VGND 0.01123f
C44046 VPWR.n1544 VGND 0.01371f
C44047 VPWR.n1545 VGND 0.01189f
C44048 VPWR.n1546 VGND 0.01839f
C44049 VPWR.n1547 VGND 0.01197f
C44050 VPWR.n1548 VGND 0.01668f
C44051 VPWR.n1549 VGND 0.01282f
C44052 VPWR.n1550 VGND 0.01349f
C44053 VPWR.n1551 VGND 0.01199f
C44054 VPWR.n1552 VGND 0.01244f
C44055 VPWR.n1553 VGND 0.01165f
C44056 VPWR.n1554 VGND 0.01114f
C44057 VPWR.n1555 VGND 0.00823f
C44058 VPWR.n1556 VGND 0.01349f
C44059 VPWR.n1557 VGND 0.01199f
C44060 VPWR.n1558 VGND 0.01171f
C44061 VPWR.n1559 VGND 0.01114f
C44062 VPWR.n1560 VGND 0.01381f
C44063 VPWR.n1561 VGND 0.008f
C44064 VPWR.n1562 VGND 0.01266f
C44065 VPWR.n1563 VGND 0.01355f
C44066 VPWR.n1564 VGND 0.01228f
C44067 VPWR.n1565 VGND 0.01171f
C44068 VPWR.n1566 VGND 0.01355f
C44069 VPWR.n1567 VGND 0.01228f
C44070 VPWR.n1568 VGND 0.01171f
C44071 VPWR.n1569 VGND 0.00858f
C44072 VPWR.n1570 VGND 0.01165f
C44073 VPWR.n1571 VGND 0.0262f
C44074 VPWR.t2317 VGND 0.02998f
C44075 VPWR.t2590 VGND 0.03574f
C44076 VPWR.t1903 VGND 0.04035f
C44077 VPWR.t3107 VGND 0.05996f
C44078 VPWR.t2293 VGND 0.05996f
C44079 VPWR.t2081 VGND 0.04959f
C44080 VPWR.t4580 VGND 0.02998f
C44081 VPWR.n1572 VGND 0.04675f
C44082 VPWR.n1573 VGND 0.01266f
C44083 VPWR.n1574 VGND 0.01017f
C44084 VPWR.n1575 VGND 0.00925f
C44085 VPWR.n1576 VGND 0.01396f
C44086 VPWR.n1577 VGND 0.01791f
C44087 VPWR.n1578 VGND 0.01197f
C44088 VPWR.n1579 VGND 0.01668f
C44089 VPWR.n1580 VGND 0.01544f
C44090 VPWR.n1581 VGND 0.00823f
C44091 VPWR.n1582 VGND 0.01165f
C44092 VPWR.n1583 VGND 0.01355f
C44093 VPWR.n1584 VGND 0.01228f
C44094 VPWR.n1585 VGND 0.01171f
C44095 VPWR.n1586 VGND 0.01355f
C44096 VPWR.n1587 VGND 0.01228f
C44097 VPWR.n1588 VGND 0.01433f
C44098 VPWR.n1589 VGND 0.0063f
C44099 VPWR.n1590 VGND 0.01431f
C44100 VPWR.n1591 VGND 0.01186f
C44101 VPWR.n1592 VGND 0.00915f
C44102 VPWR.n1593 VGND 0.00915f
C44103 VPWR.n1594 VGND 0.01251f
C44104 VPWR.n1595 VGND 0.01334f
C44105 VPWR.n1596 VGND 0.01161f
C44106 VPWR.n1597 VGND 0.00896f
C44107 VPWR.n1598 VGND 0.01077f
C44108 VPWR.n1599 VGND 0.01189f
C44109 VPWR.n1600 VGND 0.00823f
C44110 VPWR.n1601 VGND 0.01392f
C44111 VPWR.n1602 VGND 0.02379f
C44112 VPWR.n1603 VGND 0.0171f
C44113 VPWR.n1604 VGND 0.02092f
C44114 VPWR.n1605 VGND 0.01407f
C44115 VPWR.n1606 VGND 0.20174f
C44116 VPWR.n1607 VGND 0.00836f
C44117 VPWR.n1608 VGND 0.00941f
C44118 VPWR.n1609 VGND 0.00967f
C44119 VPWR.n1610 VGND 0.00673f
C44120 VPWR.n1611 VGND 0.00728f
C44121 VPWR.n1612 VGND 0.00963f
C44122 VPWR.n1613 VGND 0.01585f
C44123 VPWR.n1614 VGND 0.01628f
C44124 VPWR.n1615 VGND 0.01272f
C44125 VPWR.n1616 VGND 0.016f
C44126 VPWR.n1617 VGND 0.00984f
C44127 VPWR.n1618 VGND 0.00574f
C44128 VPWR.n1619 VGND 0.00944f
C44129 VPWR.n1620 VGND 0.01171f
C44130 VPWR.n1621 VGND 0.01257f
C44131 VPWR.n1622 VGND 0.00486f
C44132 VPWR.n1623 VGND 0.00875f
C44133 VPWR.n1624 VGND 0.01134f
C44134 VPWR.n1625 VGND 0.01125f
C44135 VPWR.n1626 VGND 0.00965f
C44136 VPWR.n1627 VGND 0.00816f
C44137 VPWR.n1628 VGND 0.00713f
C44138 VPWR.n1629 VGND 0.00673f
C44139 VPWR.n1630 VGND 0.01035f
C44140 VPWR.n1631 VGND 0.00827f
C44141 VPWR.n1632 VGND 0.00657f
C44142 VPWR.n1633 VGND 0.00564f
C44143 VPWR.n1634 VGND 0.00796f
C44144 VPWR.n1635 VGND 0.00369f
C44145 VPWR.n1636 VGND 0.00691f
C44146 VPWR.n1637 VGND 0.01189f
C44147 VPWR.n1638 VGND 0.00296f
C44148 VPWR.n1639 VGND 0.0091f
C44149 VPWR.n1640 VGND 0.20174f
C44150 VPWR.n1641 VGND 0.13412f
C44151 VPWR.n1642 VGND 0.01078f
C44152 VPWR.n1643 VGND 0.00704f
C44153 VPWR.n1644 VGND 0.01216f
C44154 VPWR.n1645 VGND 0.00921f
C44155 VPWR.n1646 VGND 0.0093f
C44156 VPWR.n1647 VGND 0.01056f
C44157 VPWR.n1648 VGND 0.01048f
C44158 VPWR.n1649 VGND 0.00494f
C44159 VPWR.n1650 VGND 0.00732f
C44160 VPWR.n1651 VGND 0.0051f
C44161 VPWR.n1652 VGND 0.00284f
C44162 VPWR.n1653 VGND 0.00637f
C44163 VPWR.n1654 VGND 0.01259f
C44164 VPWR.n1655 VGND 0.01189f
C44165 VPWR.n1656 VGND 0.00708f
C44166 VPWR.n1657 VGND 0.00925f
C44167 VPWR.n1658 VGND 0.00853f
C44168 VPWR.n1659 VGND 0.00848f
C44169 VPWR.n1660 VGND 0.01108f
C44170 VPWR.n1661 VGND 0.01146f
C44171 VPWR.n1662 VGND 0.0102f
C44172 VPWR.n1663 VGND 0.00984f
C44173 VPWR.n1664 VGND 0.00829f
C44174 VPWR.n1665 VGND 0.01015f
C44175 VPWR.n1666 VGND 0.00434f
C44176 VPWR.n1667 VGND 0.00655f
C44177 VPWR.n1668 VGND 0.01164f
C44178 VPWR.n1669 VGND 0.00663f
C44179 VPWR.n1670 VGND 0.00769f
C44180 VPWR.n1671 VGND 0.0056f
C44181 VPWR.n1672 VGND 0.00814f
C44182 VPWR.n1673 VGND 0.00594f
C44183 VPWR.n1674 VGND 0.13412f
C44184 VPWR.n1675 VGND 0.13412f
C44185 VPWR.n1676 VGND 0.00631f
C44186 VPWR.n1677 VGND 0.00524f
C44187 VPWR.n1678 VGND 0.01118f
C44188 VPWR.n1679 VGND 0.00883f
C44189 VPWR.n1680 VGND 0.00585f
C44190 VPWR.n1681 VGND 0.00879f
C44191 VPWR.n1682 VGND 0.01008f
C44192 VPWR.n1683 VGND 0.01174f
C44193 VPWR.n1684 VGND 0.00552f
C44194 VPWR.n1685 VGND 0.00884f
C44195 VPWR.n1686 VGND 0.01165f
C44196 VPWR.n1687 VGND 0.01072f
C44197 VPWR.n1688 VGND 0.00992f
C44198 VPWR.n1689 VGND 0.00437f
C44199 VPWR.n1690 VGND 0.00999f
C44200 VPWR.n1691 VGND 0.008f
C44201 VPWR.n1692 VGND 0.00588f
C44202 VPWR.n1693 VGND 0.00855f
C44203 VPWR.n1694 VGND 0.00791f
C44204 VPWR.n1695 VGND 0.00593f
C44205 VPWR.n1696 VGND 0.00655f
C44206 VPWR.n1697 VGND 0.00636f
C44207 VPWR.n1698 VGND 0.01055f
C44208 VPWR.n1699 VGND 0.00946f
C44209 VPWR.n1700 VGND 0.00938f
C44210 VPWR.n1701 VGND 0.0091f
C44211 VPWR.n1702 VGND 0.00544f
C44212 VPWR.n1703 VGND 0.01158f
C44213 VPWR.n1704 VGND 0.00751f
C44214 VPWR.n1705 VGND 0.00792f
C44215 VPWR.n1706 VGND 0.00422f
C44216 VPWR.n1707 VGND 0.00597f
C44217 VPWR.n1708 VGND 0.13412f
C44218 VPWR.n1709 VGND 0.13412f
C44219 VPWR.n1710 VGND 0.00821f
C44220 VPWR.n1711 VGND 0.00422f
C44221 VPWR.n1712 VGND 0.00564f
C44222 VPWR.n1713 VGND 0.00993f
C44223 VPWR.n1714 VGND 0.00642f
C44224 VPWR.n1715 VGND 0.01251f
C44225 VPWR.n1716 VGND 0.0063f
C44226 VPWR.n1717 VGND 0.00584f
C44227 VPWR.n1718 VGND 0.00655f
C44228 VPWR.n1719 VGND 0.00622f
C44229 VPWR.n1720 VGND 0.00443f
C44230 VPWR.n1721 VGND 0.00706f
C44231 VPWR.n1722 VGND 0.01287f
C44232 VPWR.n1723 VGND 0.01588f
C44233 VPWR.n1724 VGND 0.02059f
C44234 VPWR.n1725 VGND 0.01476f
C44235 VPWR.n1726 VGND 0.01588f
C44236 VPWR.n1727 VGND 0.01144f
C44237 VPWR.n1728 VGND 0.01288f
C44238 VPWR.n1729 VGND 0.00983f
C44239 VPWR.n1730 VGND 0.00963f
C44240 VPWR.n1731 VGND 0.00659f
C44241 VPWR.n1732 VGND 0.00805f
C44242 VPWR.n1733 VGND 0.00416f
C44243 VPWR.n1734 VGND 0.00709f
C44244 VPWR.n1735 VGND 0.00693f
C44245 VPWR.n1736 VGND 0.00848f
C44246 VPWR.n1737 VGND 0.01123f
C44247 VPWR.n1738 VGND 0.00392f
C44248 VPWR.n1739 VGND 0.01013f
C44249 VPWR.n1740 VGND 0.01053f
C44250 VPWR.n1741 VGND 0.00402f
C44251 VPWR.n1742 VGND 0.00913f
C44252 VPWR.n1743 VGND 0.00743f
C44253 VPWR.n1744 VGND 0.01189f
C44254 VPWR.n1745 VGND 0.00784f
C44255 VPWR.n1746 VGND 0.00796f
C44256 VPWR.n1747 VGND 0.00827f
C44257 VPWR.n1748 VGND 0.00553f
C44258 VPWR.n1749 VGND 0.00553f
C44259 VPWR.n1750 VGND 0.00827f
C44260 VPWR.n1751 VGND 0.00796f
C44261 VPWR.n1752 VGND 0.00951f
C44262 VPWR.n1753 VGND 0.00907f
C44263 VPWR.n1754 VGND 0.00573f
C44264 VPWR.n1755 VGND 0.00695f
C44265 VPWR.n1756 VGND 0.01077f
C44266 VPWR.n1757 VGND 0.00501f
C44267 VPWR.n1758 VGND 0.00724f
C44268 VPWR.n1759 VGND 0.00775f
C44269 VPWR.n1760 VGND 0.00609f
C44270 VPWR.t30 VGND 0.00379f
C44271 VPWR.t276 VGND 0.00164f
C44272 VPWR.t278 VGND 0.00227f
C44273 VPWR.n1761 VGND 0.00392f
C44274 VPWR.t242 VGND 0.00164f
C44275 VPWR.t236 VGND 0.00227f
C44276 VPWR.n1762 VGND 0.00392f
C44277 VPWR.t32 VGND 0.00147f
C44278 VPWR.t34 VGND 0.00147f
C44279 VPWR.n1763 VGND 0.00295f
C44280 VPWR.t294 VGND 0.00164f
C44281 VPWR.t290 VGND 0.00227f
C44282 VPWR.n1764 VGND 0.00392f
C44283 VPWR.t292 VGND 0.00425f
C44284 VPWR.t6889 VGND 0.00394f
C44285 VPWR.t36 VGND 0.00166f
C44286 VPWR.t5591 VGND 0.00183f
C44287 VPWR.n1765 VGND 0.0043f
C44288 VPWR.t6590 VGND 0.00394f
C44289 VPWR.t2546 VGND 0.00132f
C44290 VPWR.t2538 VGND 0.00132f
C44291 VPWR.n1766 VGND 0.00266f
C44292 VPWR.n1767 VGND 0.01089f
C44293 VPWR.n1768 VGND 0.01031f
C44294 VPWR.n1769 VGND 0.00241f
C44295 VPWR.n1770 VGND 0.009f
C44296 VPWR.n1771 VGND 0.01353f
C44297 VPWR.n1772 VGND 0.00916f
C44298 VPWR.n1773 VGND 0.00811f
C44299 VPWR.n1774 VGND 0.0135f
C44300 VPWR.n1775 VGND 0.00954f
C44301 VPWR.n1776 VGND 0.00862f
C44302 VPWR.n1777 VGND 0.0122f
C44303 VPWR.n1778 VGND 0.02548f
C44304 VPWR.t275 VGND 0.01395f
C44305 VPWR.t29 VGND 0.02581f
C44306 VPWR.t277 VGND 0.02804f
C44307 VPWR.t4694 VGND 0.02428f
C44308 VPWR.t241 VGND 0.02211f
C44309 VPWR.t4681 VGND 0.02428f
C44310 VPWR.t235 VGND 0.02645f
C44311 VPWR.t31 VGND 0.02428f
C44312 VPWR.t293 VGND 0.02211f
C44313 VPWR.t33 VGND 0.02428f
C44314 VPWR.t289 VGND 0.02645f
C44315 VPWR.t4697 VGND 0.02428f
C44316 VPWR.t291 VGND 0.02211f
C44317 VPWR.t4689 VGND 0.03328f
C44318 VPWR.t35 VGND 0.01227f
C44319 VPWR.t6888 VGND 0.02556f
C44320 VPWR.t6589 VGND 0.02445f
C44321 VPWR.t5590 VGND 0.02445f
C44322 VPWR.t2545 VGND 0.04141f
C44323 VPWR.t3623 VGND 0.02277f
C44324 VPWR.t2537 VGND 0.02277f
C44325 VPWR.t3569 VGND 0.02277f
C44326 VPWR.t5594 VGND 0.02322f
C44327 VPWR.t3570 VGND 0.02277f
C44328 VPWR.t5596 VGND 0.025f
C44329 VPWR.t3622 VGND 0.02277f
C44330 VPWR.t2543 VGND 0.02277f
C44331 VPWR.t2457 VGND 0.02277f
C44332 VPWR.t2539 VGND 0.02422f
C44333 VPWR.t5592 VGND 0.02355f
C44334 VPWR.t2455 VGND 0.01395f
C44335 VPWR.n1779 VGND 0.01912f
C44336 VPWR.t6425 VGND 0.00431f
C44337 VPWR.t1786 VGND 0.00433f
C44338 VPWR.t5600 VGND 0.00429f
C44339 VPWR.t974 VGND 0.00425f
C44340 VPWR.t5881 VGND 0.00431f
C44341 VPWR.t6951 VGND 0.00307f
C44342 VPWR.t6289 VGND 0.00114f
C44343 VPWR.t2165 VGND 0.00114f
C44344 VPWR.n1780 VGND 0.00229f
C44345 VPWR.t4822 VGND 0.00307f
C44346 VPWR.t5119 VGND 0.00203f
C44347 VPWR.t2167 VGND 0.00431f
C44348 VPWR.t6858 VGND 0.0018f
C44349 VPWR.t2067 VGND 0.00181f
C44350 VPWR.n1781 VGND 0.00494f
C44351 VPWR.t6424 VGND 0.0298f
C44352 VPWR.t1785 VGND 0.02612f
C44353 VPWR.t4687 VGND 0.0173f
C44354 VPWR.t5599 VGND 0.05034f
C44355 VPWR.t973 VGND 0.025f
C44356 VPWR.t5868 VGND 0.02768f
C44357 VPWR.t3910 VGND 0.025f
C44358 VPWR.t568 VGND 0.02277f
C44359 VPWR.t3568 VGND 0.0221f
C44360 VPWR.t4830 VGND 0.0125f
C44361 VPWR.t5880 VGND 0.02612f
C44362 VPWR.t6950 VGND 0.02277f
C44363 VPWR.t569 VGND 0.02277f
C44364 VPWR.t6288 VGND 0.025f
C44365 VPWR.t201 VGND 0.02277f
C44366 VPWR.t2164 VGND 0.03271f
C44367 VPWR.t4821 VGND 0.02545f
C44368 VPWR.t5118 VGND 0.0125f
C44369 VPWR.t2166 VGND 0.02199f
C44370 VPWR.t6857 VGND 0.02277f
C44371 VPWR.t6381 VGND 0.02992f
C44372 VPWR.t2066 VGND 0.025f
C44373 VPWR.t206 VGND 0.04521f
C44374 VPWR.t2021 VGND 0.0202f
C44375 VPWR.t5913 VGND 0.0173f
C44376 VPWR.t4708 VGND 0.01741f
C44377 VPWR.t3872 VGND 0.03326f
C44378 VPWR.t5914 VGND 0.04443f
C44379 VPWR.t2618 VGND 0.03885f
C44380 VPWR.t3868 VGND 0.03271f
C44381 VPWR.t3870 VGND 0.01395f
C44382 VPWR.t6663 VGND 0.02456f
C44383 VPWR.t6396 VGND 0.03605f
C44384 VPWR.t4876 VGND 0.03494f
C44385 VPWR.t1665 VGND 0.0336f
C44386 VPWR.t1537 VGND 0.02147f
C44387 VPWR.t5641 VGND 0.01772f
C44388 VPWR.n1782 VGND 0.03945f
C44389 VPWR.t6399 VGND 0.02478f
C44390 VPWR.t460 VGND 0.03014f
C44391 VPWR.t6220 VGND 0.02411f
C44392 VPWR.t5642 VGND 0.04387f
C44393 VPWR.t6398 VGND 0.03951f
C44394 VPWR.t3237 VGND 0.03181f
C44395 VPWR.t1667 VGND 0.03271f
C44396 VPWR.t2023 VGND 0.0173f
C44397 VPWR.t1790 VGND 0.02768f
C44398 VPWR.t1668 VGND 0.03271f
C44399 VPWR.n1783 VGND 0.03062f
C44400 VPWR.t2022 VGND 0.00427f
C44401 VPWR.t1791 VGND 0.00433f
C44402 VPWR.t1669 VGND 0.00107f
C44403 VPWR.n1784 VGND 0.00292f
C44404 VPWR.t3238 VGND 0.00433f
C44405 VPWR.t6221 VGND 0.00433f
C44406 VPWR.n1785 VGND 0.00115f
C44407 VPWR.t1538 VGND 0.00433f
C44408 VPWR.t4877 VGND 0.00433f
C44409 VPWR.t1666 VGND 0.00255f
C44410 VPWR.t3871 VGND 0.00603f
C44411 VPWR.t6397 VGND 0.00116f
C44412 VPWR.t6664 VGND 0.00116f
C44413 VPWR.n1786 VGND 0.00236f
C44414 VPWR.t2619 VGND 0.00433f
C44415 VPWR.n1787 VGND 0.01023f
C44416 VPWR.n1788 VGND 0.00319f
C44417 VPWR.n1789 VGND 0.01116f
C44418 VPWR.n1790 VGND 0.01081f
C44419 VPWR.n1791 VGND 0.01302f
C44420 VPWR.n1792 VGND 0.01197f
C44421 VPWR.n1793 VGND 0.00899f
C44422 VPWR.n1794 VGND 0.01333f
C44423 VPWR.n1795 VGND 0.01544f
C44424 VPWR.n1796 VGND 0.00462f
C44425 VPWR.n1797 VGND 0.00693f
C44426 VPWR.n1798 VGND 0.00624f
C44427 VPWR.n1799 VGND 0.00928f
C44428 VPWR.n1800 VGND 0.00417f
C44429 VPWR.n1801 VGND 0.00966f
C44430 VPWR.n1802 VGND 0.00464f
C44431 VPWR.n1803 VGND 0.00456f
C44432 VPWR.n1804 VGND 0.00364f
C44433 VPWR.n1805 VGND 0.00734f
C44434 VPWR.n1806 VGND 0.00955f
C44435 VPWR.n1807 VGND 0.01182f
C44436 VPWR.n1808 VGND 0.01164f
C44437 VPWR.n1809 VGND 0.008f
C44438 VPWR.n1810 VGND 0.00668f
C44439 VPWR.n1811 VGND 0.01015f
C44440 VPWR.n1812 VGND 0.00882f
C44441 VPWR.n1813 VGND 0.00476f
C44442 VPWR.n1814 VGND 0.00745f
C44443 VPWR.n1815 VGND 0.01115f
C44444 VPWR.n1816 VGND 0.13412f
C44445 VPWR.n1817 VGND 0.13412f
C44446 VPWR.n1818 VGND 0.0114f
C44447 VPWR.n1819 VGND 0.00538f
C44448 VPWR.n1820 VGND 0.00849f
C44449 VPWR.n1821 VGND 0.01037f
C44450 VPWR.n1822 VGND 0.01478f
C44451 VPWR.n1823 VGND 0.00811f
C44452 VPWR.n1824 VGND 0.00789f
C44453 VPWR.n1825 VGND 0.01481f
C44454 VPWR.n1826 VGND 0.00938f
C44455 VPWR.n1827 VGND 0.00348f
C44456 VPWR.n1828 VGND 0.00676f
C44457 VPWR.n1829 VGND 0.01165f
C44458 VPWR.n1830 VGND 0.00507f
C44459 VPWR.n1831 VGND 0.01028f
C44460 VPWR.n1832 VGND 0.00592f
C44461 VPWR.n1833 VGND 0.00882f
C44462 VPWR.n1834 VGND 0.00454f
C44463 VPWR.n1835 VGND 0.01068f
C44464 VPWR.n1836 VGND 0.00653f
C44465 VPWR.n1837 VGND 0.00708f
C44466 VPWR.n1838 VGND 0.01172f
C44467 VPWR.n1839 VGND 0.01754f
C44468 VPWR.n1840 VGND 0.021f
C44469 VPWR.n1841 VGND 0.01282f
C44470 VPWR.n1842 VGND 0.00983f
C44471 VPWR.n1843 VGND 0.00793f
C44472 VPWR.n1844 VGND 0.00879f
C44473 VPWR.n1845 VGND 0.13412f
C44474 VPWR.n1846 VGND 0.13412f
C44475 VPWR.n1847 VGND 0.00594f
C44476 VPWR.n1848 VGND 0.00722f
C44477 VPWR.n1849 VGND 0.00952f
C44478 VPWR.n1850 VGND 0.00759f
C44479 VPWR.n1851 VGND 0.00823f
C44480 VPWR.n1852 VGND 0.00552f
C44481 VPWR.n1853 VGND 0.00431f
C44482 VPWR.n1854 VGND 0.00571f
C44483 VPWR.n1855 VGND 0.01006f
C44484 VPWR.n1856 VGND 0.00382f
C44485 VPWR.n1857 VGND 0.00979f
C44486 VPWR.n1858 VGND 0.01136f
C44487 VPWR.n1859 VGND 0.00894f
C44488 VPWR.n1860 VGND 0.0051f
C44489 VPWR.n1861 VGND 0.01165f
C44490 VPWR.n1862 VGND 0.01107f
C44491 VPWR.n1863 VGND 0.01056f
C44492 VPWR.n1864 VGND 0.00713f
C44493 VPWR.n1865 VGND 0.00809f
C44494 VPWR.n1866 VGND 0.01451f
C44495 VPWR.n1867 VGND 0.01544f
C44496 VPWR.n1868 VGND 0.00552f
C44497 VPWR.n1869 VGND 0.00811f
C44498 VPWR.n1870 VGND 0.00855f
C44499 VPWR.n1871 VGND 0.00728f
C44500 VPWR.n1872 VGND 0.00664f
C44501 VPWR.n1873 VGND 0.00881f
C44502 VPWR.n1874 VGND 0.00561f
C44503 VPWR.n1875 VGND 0.00819f
C44504 VPWR.n1876 VGND 0.0063f
C44505 VPWR.n1877 VGND 0.01165f
C44506 VPWR.n1878 VGND 0.00642f
C44507 VPWR.n1879 VGND 0.01353f
C44508 VPWR.n1880 VGND 0.00842f
C44509 VPWR.n1881 VGND 0.00821f
C44510 VPWR.n1882 VGND 0.13412f
C44511 VPWR.n1883 VGND 0.13412f
C44512 VPWR.n1884 VGND 0.00568f
C44513 VPWR.n1885 VGND 0.00743f
C44514 VPWR.n1886 VGND 0.00685f
C44515 VPWR.n1887 VGND 0.00655f
C44516 VPWR.n1888 VGND 0.00655f
C44517 VPWR.n1889 VGND 0.0077f
C44518 VPWR.n1890 VGND 0.0077f
C44519 VPWR.n1891 VGND 0.00655f
C44520 VPWR.n1892 VGND 0.00655f
C44521 VPWR.n1893 VGND 0.0054f
C44522 VPWR.n1894 VGND 0.0054f
C44523 VPWR.n1895 VGND 0.01077f
C44524 VPWR.n1896 VGND 0.00642f
C44525 VPWR.n1897 VGND 0.00584f
C44526 VPWR.n1898 VGND 0.0077f
C44527 VPWR.n1899 VGND 0.0054f
C44528 VPWR.n1900 VGND 0.01055f
C44529 VPWR.n1901 VGND 0.01138f
C44530 VPWR.n1902 VGND 0.00974f
C44531 VPWR.n1903 VGND 0.01085f
C44532 VPWR.n1904 VGND 0.0085f
C44533 VPWR.n1905 VGND 0.008f
C44534 VPWR.n1906 VGND 0.00661f
C44535 VPWR.n1907 VGND 0.00844f
C44536 VPWR.n1908 VGND 0.00675f
C44537 VPWR.n1909 VGND 0.00943f
C44538 VPWR.n1910 VGND 0.0085f
C44539 VPWR.n1911 VGND 0.008f
C44540 VPWR.n1912 VGND 0.00661f
C44541 VPWR.n1913 VGND 0.01266f
C44542 VPWR.n1914 VGND 0.00788f
C44543 VPWR.n1915 VGND 0.00705f
C44544 VPWR.n1916 VGND 0.008f
C44545 VPWR.n1917 VGND 0.00872f
C44546 VPWR.n1918 VGND 0.00767f
C44547 VPWR.n1919 VGND 0.00685f
C44548 VPWR.n1920 VGND 0.00943f
C44549 VPWR.n1921 VGND 0.00729f
C44550 VPWR.n1922 VGND 0.00443f
C44551 VPWR.n1923 VGND 0.00779f
C44552 VPWR.n1924 VGND 0.0083f
C44553 VPWR.n1925 VGND 0.13412f
C44554 VPWR.t4065 VGND 0.00433f
C44555 VPWR.n1926 VGND 0.00899f
C44556 VPWR.t6078 VGND 0.00433f
C44557 VPWR.t3851 VGND 0.00433f
C44558 VPWR.t1673 VGND 0.00433f
C44559 VPWR.t1261 VGND 0.00433f
C44560 VPWR.t1718 VGND 0.00433f
C44561 VPWR.t1675 VGND 0.00433f
C44562 VPWR.t2536 VGND 0.00433f
C44563 VPWR.t632 VGND 0.00433f
C44564 VPWR.t1986 VGND 0.00433f
C44565 VPWR.t2090 VGND 0.00433f
C44566 VPWR.n1927 VGND 0.00676f
C44567 VPWR.n1928 VGND 0.00912f
C44568 VPWR.n1929 VGND 0.00974f
C44569 VPWR.n1930 VGND 0.01085f
C44570 VPWR.n1931 VGND 0.01085f
C44571 VPWR.n1932 VGND 0.01085f
C44572 VPWR.n1933 VGND 0.00676f
C44573 VPWR.n1934 VGND 0.008f
C44574 VPWR.n1935 VGND 0.00661f
C44575 VPWR.t3850 VGND 0.03271f
C44576 VPWR.t1672 VGND 0.0298f
C44577 VPWR.t1260 VGND 0.03271f
C44578 VPWR.t1717 VGND 0.0173f
C44579 VPWR.t1674 VGND 0.04521f
C44580 VPWR.t2535 VGND 0.05001f
C44581 VPWR.t631 VGND 0.05001f
C44582 VPWR.t1985 VGND 0.05001f
C44583 VPWR.t2089 VGND 0.05001f
C44584 VPWR.t4064 VGND 0.0298f
C44585 VPWR.t6077 VGND 0.04122f
C44586 VPWR.t3057 VGND 0.00433f
C44587 VPWR.t5325 VGND 0.00433f
C44588 VPWR.t6161 VGND 0.00433f
C44589 VPWR.t2248 VGND 0.00433f
C44590 VPWR.t3051 VGND 0.00433f
C44591 VPWR.t1722 VGND 0.00433f
C44592 VPWR.t59 VGND 0.00433f
C44593 VPWR.t5106 VGND 0.00433f
C44594 VPWR.t4299 VGND 0.00433f
C44595 VPWR.t1990 VGND 0.00433f
C44596 VPWR.t4863 VGND 0.00433f
C44597 VPWR.t4067 VGND 0.00433f
C44598 VPWR.t5448 VGND 0.00433f
C44599 VPWR.t3860 VGND 0.00433f
C44600 VPWR.t4622 VGND 0.00433f
C44601 VPWR.t6452 VGND 0.00433f
C44602 VPWR.t5966 VGND 0.00433f
C44603 VPWR.t3056 VGND 0.05001f
C44604 VPWR.t2247 VGND 0.08271f
C44605 VPWR.t1721 VGND 0.10001f
C44606 VPWR.t58 VGND 0.10001f
C44607 VPWR.t1989 VGND 0.10001f
C44608 VPWR.t4066 VGND 0.10001f
C44609 VPWR.t3859 VGND 0.10001f
C44610 VPWR.t4621 VGND 0.06731f
C44611 VPWR.n1936 VGND 0.03642f
C44612 VPWR.t1390 VGND 0.00473f
C44613 VPWR.t5884 VGND 0.00473f
C44614 VPWR.t1388 VGND 0.00427f
C44615 VPWR.t5886 VGND 0.00427f
C44616 VPWR.t6132 VGND 0.00427f
C44617 VPWR.t2998 VGND 0.00473f
C44618 VPWR.t6130 VGND 0.00473f
C44619 VPWR.t3000 VGND 0.00427f
C44620 VPWR.t6255 VGND 0.00427f
C44621 VPWR.t2370 VGND 0.00427f
C44622 VPWR.t6253 VGND 0.00473f
C44623 VPWR.t2368 VGND 0.00473f
C44624 VPWR.t5890 VGND 0.00427f
C44625 VPWR.t2767 VGND 0.00433f
C44626 VPWR.t5888 VGND 0.00473f
C44627 VPWR.t1628 VGND 0.00433f
C44628 VPWR.t1193 VGND 0.00433f
C44629 VPWR.t5845 VGND 0.00433f
C44630 VPWR.t5965 VGND 0.0173f
C44631 VPWR.t1389 VGND 0.03538f
C44632 VPWR.t5883 VGND 0.02791f
C44633 VPWR.t1387 VGND 0.02712f
C44634 VPWR.t5885 VGND 0.0125f
C44635 VPWR.t6131 VGND 0.03248f
C44636 VPWR.t2997 VGND 0.02791f
C44637 VPWR.t6129 VGND 0.02791f
C44638 VPWR.t2999 VGND 0.03248f
C44639 VPWR.t6254 VGND 0.0125f
C44640 VPWR.t2369 VGND 0.02712f
C44641 VPWR.t6252 VGND 0.02791f
C44642 VPWR.t2367 VGND 0.03538f
C44643 VPWR.t5889 VGND 0.0221f
C44644 VPWR.t5887 VGND 0.03271f
C44645 VPWR.t2766 VGND 0.03248f
C44646 VPWR.t1627 VGND 0.03271f
C44647 VPWR.t1192 VGND 0.04231f
C44648 VPWR.t5844 VGND 0.0202f
C44649 VPWR.n1937 VGND 0.05372f
C44650 VPWR.t6074 VGND 0.00433f
C44651 VPWR.t4927 VGND 0.00433f
C44652 VPWR.t5324 VGND 0.00433f
C44653 VPWR.t3071 VGND 0.00473f
C44654 VPWR.t6328 VGND 0.00433f
C44655 VPWR.t3073 VGND 0.00427f
C44656 VPWR.t5695 VGND 0.00473f
C44657 VPWR.t5526 VGND 0.00473f
C44658 VPWR.t5693 VGND 0.00427f
C44659 VPWR.t4412 VGND 0.00427f
C44660 VPWR.t5528 VGND 0.00427f
C44661 VPWR.t2122 VGND 0.00473f
C44662 VPWR.t4414 VGND 0.00473f
C44663 VPWR.t2120 VGND 0.00427f
C44664 VPWR.t5421 VGND 0.00433f
C44665 VPWR.t2071 VGND 0.00433f
C44666 VPWR.t4646 VGND 0.00433f
C44667 VPWR.t2852 VGND 0.00433f
C44668 VPWR.t2020 VGND 0.00433f
C44669 VPWR.t4926 VGND 0.05481f
C44670 VPWR.t5323 VGND 0.03538f
C44671 VPWR.t3070 VGND 0.03058f
C44672 VPWR.t3072 VGND 0.03963f
C44673 VPWR.t6327 VGND 0.025f
C44674 VPWR.t5694 VGND 0.03538f
C44675 VPWR.t5525 VGND 0.02791f
C44676 VPWR.t5692 VGND 0.01462f
C44677 VPWR.t5527 VGND 0.0154f
C44678 VPWR.t4411 VGND 0.03003f
C44679 VPWR.t4413 VGND 0.03326f
C44680 VPWR.t2121 VGND 0.03248f
C44681 VPWR.t2119 VGND 0.0125f
C44682 VPWR.t5420 VGND 0.03271f
C44683 VPWR.t2070 VGND 0.0173f
C44684 VPWR.t4645 VGND 0.04521f
C44685 VPWR.t2851 VGND 0.0298f
C44686 VPWR.t2673 VGND 0.01775f
C44687 VPWR.t121 VGND 0.0202f
C44688 VPWR.t786 VGND 0.01931f
C44689 VPWR.t3235 VGND 0.02612f
C44690 VPWR.t1463 VGND 0.04063f
C44691 VPWR.t120 VGND 0.02389f
C44692 VPWR.t2993 VGND 0.02969f
C44693 VPWR.n1938 VGND 0.03208f
C44694 VPWR.t5423 VGND 0.0211f
C44695 VPWR.t4264 VGND 0.04822f
C44696 VPWR.t127 VGND 0.05001f
C44697 VPWR.t5511 VGND 0.02277f
C44698 VPWR.t6756 VGND 0.0298f
C44699 VPWR.t2634 VGND 0.01395f
C44700 VPWR.t2646 VGND 0.03416f
C44701 VPWR.t6619 VGND 0.04085f
C44702 VPWR.t1280 VGND 0.025f
C44703 VPWR.t305 VGND 0.03192f
C44704 VPWR.t193 VGND 0.04085f
C44705 VPWR.t1792 VGND 0.03829f
C44706 VPWR.t4427 VGND 0.0298f
C44707 VPWR.t3624 VGND 0.03271f
C44708 VPWR.t2019 VGND 0.04122f
C44709 VPWR.t3625 VGND 0.00433f
C44710 VPWR.t4428 VGND 0.00433f
C44711 VPWR.t1793 VGND 0.00433f
C44712 VPWR.t194 VGND 0.00473f
C44713 VPWR.t1281 VGND 0.00433f
C44714 VPWR.t2635 VGND 0.00433f
C44715 VPWR.t2647 VGND 0.00498f
C44716 VPWR.t5512 VGND 0.00433f
C44717 VPWR.t6757 VGND 0.00116f
C44718 VPWR.t128 VGND 0.00116f
C44719 VPWR.n1939 VGND 0.00236f
C44720 VPWR.t4265 VGND 0.00433f
C44721 VPWR.t5424 VGND 0.00255f
C44722 VPWR.t2994 VGND 0.00433f
C44723 VPWR.t787 VGND 0.00433f
C44724 VPWR.n1940 VGND 0.01135f
C44725 VPWR.n1941 VGND 0.01699f
C44726 VPWR.n1942 VGND 0.01013f
C44727 VPWR.n1943 VGND 0.00992f
C44728 VPWR.n1944 VGND 0.00784f
C44729 VPWR.n1945 VGND 0.0064f
C44730 VPWR.n1946 VGND 0.01022f
C44731 VPWR.n1947 VGND 0.01147f
C44732 VPWR.n1948 VGND 0.00992f
C44733 VPWR.n1949 VGND 0.00933f
C44734 VPWR.n1950 VGND 0.01005f
C44735 VPWR.n1951 VGND 0.008f
C44736 VPWR.n1952 VGND 0.00661f
C44737 VPWR.n1953 VGND 0.01266f
C44738 VPWR.n1954 VGND 0.00735f
C44739 VPWR.n1955 VGND 0.00912f
C44740 VPWR.n1956 VGND 0.00912f
C44741 VPWR.n1957 VGND 0.00627f
C44742 VPWR.n1958 VGND 0.00661f
C44743 VPWR.n1959 VGND 0.00635f
C44744 VPWR.n1960 VGND 0.0054f
C44745 VPWR.n1961 VGND 0.0054f
C44746 VPWR.n1962 VGND 0.0077f
C44747 VPWR.n1963 VGND 0.00708f
C44748 VPWR.n1964 VGND 0.00646f
C44749 VPWR.n1965 VGND 0.00593f
C44750 VPWR.n1966 VGND 0.00878f
C44751 VPWR.n1967 VGND 0.00822f
C44752 VPWR.n1968 VGND 0.00627f
C44753 VPWR.n1969 VGND 0.00655f
C44754 VPWR.n1970 VGND 0.00964f
C44755 VPWR.n1971 VGND 0.01303f
C44756 VPWR.n1972 VGND 0.01189f
C44757 VPWR.n1973 VGND 0.00909f
C44758 VPWR.n1974 VGND 0.00718f
C44759 VPWR.n1975 VGND 0.00893f
C44760 VPWR.n1976 VGND 0.00665f
C44761 VPWR.n1977 VGND 0.00743f
C44762 VPWR.n1978 VGND 0.00685f
C44763 VPWR.n1979 VGND 0.00776f
C44764 VPWR.n1980 VGND 0.00584f
C44765 VPWR.n1981 VGND 0.0054f
C44766 VPWR.n1982 VGND 0.0077f
C44767 VPWR.n1983 VGND 0.00584f
C44768 VPWR.n1984 VGND 0.00698f
C44769 VPWR.n1985 VGND 0.00655f
C44770 VPWR.n1986 VGND 0.00655f
C44771 VPWR.n1987 VGND 0.00698f
C44772 VPWR.n1988 VGND 0.00584f
C44773 VPWR.n1989 VGND 0.0077f
C44774 VPWR.n1990 VGND 0.0054f
C44775 VPWR.n1991 VGND 0.0063f
C44776 VPWR.n1992 VGND 0.01165f
C44777 VPWR.n1993 VGND 0.01144f
C44778 VPWR.n1994 VGND 0.02171f
C44779 VPWR.n1995 VGND 0.02171f
C44780 VPWR.n1996 VGND 0.01577f
C44781 VPWR.n1997 VGND 0.01476f
C44782 VPWR.n1998 VGND 0.0207f
C44783 VPWR.n1999 VGND 0.02171f
C44784 VPWR.n2000 VGND 0.01935f
C44785 VPWR.n2001 VGND 0.01214f
C44786 VPWR.n2002 VGND 0.01165f
C44787 VPWR.n2003 VGND 0.00809f
C44788 VPWR.n2004 VGND 0.01004f
C44789 VPWR.n2005 VGND 0.13412f
C44790 VPWR.t4017 VGND 0.00433f
C44791 VPWR.n2006 VGND 0.00899f
C44792 VPWR.t3392 VGND 0.00433f
C44793 VPWR.t4934 VGND 0.00433f
C44794 VPWR.t6457 VGND 0.00433f
C44795 VPWR.t2777 VGND 0.00433f
C44796 VPWR.t6436 VGND 0.00433f
C44797 VPWR.t2075 VGND 0.00433f
C44798 VPWR.t1816 VGND 0.00433f
C44799 VPWR.t5027 VGND 0.00433f
C44800 VPWR.t3250 VGND 0.00433f
C44801 VPWR.t661 VGND 0.00433f
C44802 VPWR.n2007 VGND 0.00676f
C44803 VPWR.n2008 VGND 0.00912f
C44804 VPWR.n2009 VGND 0.00974f
C44805 VPWR.n2010 VGND 0.01085f
C44806 VPWR.n2011 VGND 0.01085f
C44807 VPWR.n2012 VGND 0.01085f
C44808 VPWR.n2013 VGND 0.00676f
C44809 VPWR.n2014 VGND 0.008f
C44810 VPWR.n2015 VGND 0.00661f
C44811 VPWR.t4933 VGND 0.03271f
C44812 VPWR.t6456 VGND 0.0298f
C44813 VPWR.t2776 VGND 0.03271f
C44814 VPWR.t6435 VGND 0.0173f
C44815 VPWR.t2074 VGND 0.04521f
C44816 VPWR.t1815 VGND 0.05001f
C44817 VPWR.t5026 VGND 0.05001f
C44818 VPWR.t3249 VGND 0.05001f
C44819 VPWR.t660 VGND 0.05001f
C44820 VPWR.t4016 VGND 0.0298f
C44821 VPWR.t3391 VGND 0.04122f
C44822 VPWR.t1041 VGND 0.00433f
C44823 VPWR.t4122 VGND 0.00433f
C44824 VPWR.t1345 VGND 0.00433f
C44825 VPWR.t1856 VGND 0.00433f
C44826 VPWR.t2412 VGND 0.00433f
C44827 VPWR.t1889 VGND 0.00433f
C44828 VPWR.t2157 VGND 0.00433f
C44829 VPWR.t556 VGND 0.00433f
C44830 VPWR.t2383 VGND 0.00433f
C44831 VPWR.t714 VGND 0.00433f
C44832 VPWR.t870 VGND 0.00433f
C44833 VPWR.t5756 VGND 0.00433f
C44834 VPWR.t313 VGND 0.00433f
C44835 VPWR.t5938 VGND 0.00433f
C44836 VPWR.t4846 VGND 0.00433f
C44837 VPWR.t984 VGND 0.00433f
C44838 VPWR.t5368 VGND 0.00433f
C44839 VPWR.t1040 VGND 0.03271f
C44840 VPWR.t4121 VGND 0.05001f
C44841 VPWR.t1344 VGND 0.05001f
C44842 VPWR.t1855 VGND 0.0173f
C44843 VPWR.t2411 VGND 0.04521f
C44844 VPWR.t1888 VGND 0.05001f
C44845 VPWR.t2156 VGND 0.05001f
C44846 VPWR.t555 VGND 0.05001f
C44847 VPWR.t2382 VGND 0.05001f
C44848 VPWR.t713 VGND 0.05001f
C44849 VPWR.t869 VGND 0.05001f
C44850 VPWR.t5755 VGND 0.05001f
C44851 VPWR.t312 VGND 0.05001f
C44852 VPWR.t5937 VGND 0.05001f
C44853 VPWR.t4845 VGND 0.05001f
C44854 VPWR.t983 VGND 0.0298f
C44855 VPWR.t6311 VGND 0.0202f
C44856 VPWR.t4768 VGND 0.025f
C44857 VPWR.t4056 VGND 0.04231f
C44858 VPWR.t7067 VGND 0.05001f
C44859 VPWR.t3769 VGND 0.03271f
C44860 VPWR.t1601 VGND 0.03248f
C44861 VPWR.t4529 VGND 0.02791f
C44862 VPWR.t1603 VGND 0.02712f
C44863 VPWR.t4531 VGND 0.0125f
C44864 VPWR.t2204 VGND 0.03538f
C44865 VPWR.t1403 VGND 0.02791f
C44866 VPWR.t2202 VGND 0.02712f
C44867 VPWR.t1405 VGND 0.0125f
C44868 VPWR.t2208 VGND 0.0125f
C44869 VPWR.t3172 VGND 0.02712f
C44870 VPWR.t2206 VGND 0.02791f
C44871 VPWR.t3174 VGND 0.03538f
C44872 VPWR.t5293 VGND 0.0173f
C44873 VPWR.t369 VGND 0.05001f
C44874 VPWR.t5367 VGND 0.06143f
C44875 VPWR.t370 VGND 0.00433f
C44876 VPWR.t5294 VGND 0.00433f
C44877 VPWR.t3175 VGND 0.00473f
C44878 VPWR.t2207 VGND 0.00473f
C44879 VPWR.t3173 VGND 0.00427f
C44880 VPWR.t2209 VGND 0.00427f
C44881 VPWR.t1406 VGND 0.00427f
C44882 VPWR.t2203 VGND 0.00427f
C44883 VPWR.t1404 VGND 0.00473f
C44884 VPWR.t2205 VGND 0.00473f
C44885 VPWR.t4532 VGND 0.00427f
C44886 VPWR.t1604 VGND 0.00427f
C44887 VPWR.t4530 VGND 0.00473f
C44888 VPWR.t1602 VGND 0.00473f
C44889 VPWR.t3770 VGND 0.00433f
C44890 VPWR.t7068 VGND 0.00433f
C44891 VPWR.t4057 VGND 0.00433f
C44892 VPWR.n2016 VGND 0.00738f
C44893 VPWR.n2017 VGND 0.00896f
C44894 VPWR.n2018 VGND 0.00665f
C44895 VPWR.n2019 VGND 0.0056f
C44896 VPWR.n2020 VGND 0.0054f
C44897 VPWR.n2021 VGND 0.0077f
C44898 VPWR.n2022 VGND 0.00698f
C44899 VPWR.n2023 VGND 0.00584f
C44900 VPWR.n2024 VGND 0.0054f
C44901 VPWR.n2025 VGND 0.0077f
C44902 VPWR.n2026 VGND 0.00584f
C44903 VPWR.n2027 VGND 0.00584f
C44904 VPWR.n2028 VGND 0.0077f
C44905 VPWR.n2029 VGND 0.0054f
C44906 VPWR.n2030 VGND 0.00993f
C44907 VPWR.n2031 VGND 0.00627f
C44908 VPWR.n2032 VGND 0.0085f
C44909 VPWR.n2033 VGND 0.01189f
C44910 VPWR.n2034 VGND 0.01144f
C44911 VPWR.n2035 VGND 0.01085f
C44912 VPWR.n2036 VGND 0.01085f
C44913 VPWR.n2037 VGND 0.01085f
C44914 VPWR.n2038 VGND 0.00665f
C44915 VPWR.n2039 VGND 0.00985f
C44916 VPWR.n2040 VGND 0.01085f
C44917 VPWR.n2041 VGND 0.01013f
C44918 VPWR.n2042 VGND 0.00985f
C44919 VPWR.n2043 VGND 0.01085f
C44920 VPWR.n2044 VGND 0.01085f
C44921 VPWR.n2045 VGND 0.01085f
C44922 VPWR.n2046 VGND 0.01085f
C44923 VPWR.n2047 VGND 0.01085f
C44924 VPWR.n2048 VGND 0.00676f
C44925 VPWR.n2049 VGND 0.00974f
C44926 VPWR.n2050 VGND 0.0085f
C44927 VPWR.n2051 VGND 0.01189f
C44928 VPWR.n2052 VGND 0.00809f
C44929 VPWR.n2053 VGND 0.01004f
C44930 VPWR.n2054 VGND 0.13412f
C44931 VPWR.t739 VGND 0.00433f
C44932 VPWR.n2055 VGND 0.00899f
C44933 VPWR.t410 VGND 0.00433f
C44934 VPWR.t5689 VGND 0.00433f
C44935 VPWR.t1614 VGND 0.00433f
C44936 VPWR.t5942 VGND 0.00433f
C44937 VPWR.t4626 VGND 0.00433f
C44938 VPWR.t5206 VGND 0.00433f
C44939 VPWR.t4070 VGND 0.00433f
C44940 VPWR.t5900 VGND 0.00433f
C44941 VPWR.t1000 VGND 0.00433f
C44942 VPWR.t619 VGND 0.00433f
C44943 VPWR.t3145 VGND 0.00433f
C44944 VPWR.t3088 VGND 0.00433f
C44945 VPWR.t5940 VGND 0.00433f
C44946 VPWR.t6231 VGND 0.00433f
C44947 VPWR.n2056 VGND 0.0085f
C44948 VPWR.n2057 VGND 0.00974f
C44949 VPWR.n2058 VGND 0.01085f
C44950 VPWR.n2059 VGND 0.0085f
C44951 VPWR.n2060 VGND 0.00974f
C44952 VPWR.n2061 VGND 0.01085f
C44953 VPWR.n2062 VGND 0.0085f
C44954 VPWR.n2063 VGND 0.00896f
C44955 VPWR.n2064 VGND 0.00665f
C44956 VPWR.t5205 VGND 0.03271f
C44957 VPWR.t4069 VGND 0.04231f
C44958 VPWR.t5899 VGND 0.025f
C44959 VPWR.t999 VGND 0.03271f
C44960 VPWR.t618 VGND 0.05001f
C44961 VPWR.t3144 VGND 0.04231f
C44962 VPWR.t3087 VGND 0.03271f
C44963 VPWR.t5939 VGND 0.05001f
C44964 VPWR.t6230 VGND 0.05001f
C44965 VPWR.t738 VGND 0.05001f
C44966 VPWR.t409 VGND 0.04231f
C44967 VPWR.t5688 VGND 0.03271f
C44968 VPWR.t1613 VGND 0.05001f
C44969 VPWR.t5941 VGND 0.04231f
C44970 VPWR.t4625 VGND 0.0202f
C44971 VPWR.n2065 VGND 0.05372f
C44972 VPWR.t4378 VGND 0.00433f
C44973 VPWR.t1872 VGND 0.00433f
C44974 VPWR.t5878 VGND 0.00433f
C44975 VPWR.t5275 VGND 0.00433f
C44976 VPWR.t5259 VGND 0.00433f
C44977 VPWR.t1612 VGND 0.00433f
C44978 VPWR.t2677 VGND 0.00433f
C44979 VPWR.t4405 VGND 0.00433f
C44980 VPWR.t810 VGND 0.00433f
C44981 VPWR.t5684 VGND 0.00433f
C44982 VPWR.t3814 VGND 0.00433f
C44983 VPWR.t941 VGND 0.00433f
C44984 VPWR.t5655 VGND 0.00433f
C44985 VPWR.t1871 VGND 0.08751f
C44986 VPWR.t5274 VGND 0.10001f
C44987 VPWR.t1611 VGND 0.10001f
C44988 VPWR.t2676 VGND 0.10001f
C44989 VPWR.t809 VGND 0.10001f
C44990 VPWR.t940 VGND 0.06731f
C44991 VPWR.n2066 VGND 0.03642f
C44992 VPWR.t2710 VGND 0.00433f
C44993 VPWR.t2811 VGND 0.00433f
C44994 VPWR.t5850 VGND 0.00433f
C44995 VPWR.t5654 VGND 0.0173f
C44996 VPWR.t2709 VGND 0.04521f
C44997 VPWR.t2810 VGND 0.0298f
C44998 VPWR.t1511 VGND 0.04018f
C44999 VPWR.t2365 VGND 0.02791f
C45000 VPWR.t1513 VGND 0.02712f
C45001 VPWR.t2363 VGND 0.0125f
C45002 VPWR.t3571 VGND 0.03248f
C45003 VPWR.t4060 VGND 0.02791f
C45004 VPWR.t3573 VGND 0.02791f
C45005 VPWR.t4062 VGND 0.03248f
C45006 VPWR.t4649 VGND 0.03248f
C45007 VPWR.t5131 VGND 0.02791f
C45008 VPWR.t4651 VGND 0.02791f
C45009 VPWR.t5133 VGND 0.03248f
C45010 VPWR.t966 VGND 0.03248f
C45011 VPWR.t1366 VGND 0.02791f
C45012 VPWR.t968 VGND 0.02791f
C45013 VPWR.t1368 VGND 0.03248f
C45014 VPWR.t5125 VGND 0.01172f
C45015 VPWR.t6004 VGND 0.02791f
C45016 VPWR.t5127 VGND 0.02791f
C45017 VPWR.t6002 VGND 0.01172f
C45018 VPWR.t5849 VGND 0.04122f
C45019 VPWR.t6003 VGND 0.00473f
C45020 VPWR.t5128 VGND 0.00427f
C45021 VPWR.t6005 VGND 0.00427f
C45022 VPWR.t5126 VGND 0.00473f
C45023 VPWR.t1369 VGND 0.00427f
C45024 VPWR.t969 VGND 0.00473f
C45025 VPWR.t1367 VGND 0.00473f
C45026 VPWR.t967 VGND 0.00427f
C45027 VPWR.t5134 VGND 0.00427f
C45028 VPWR.t4652 VGND 0.00473f
C45029 VPWR.t5132 VGND 0.00473f
C45030 VPWR.t4650 VGND 0.00427f
C45031 VPWR.t4063 VGND 0.00427f
C45032 VPWR.n2067 VGND 0.00745f
C45033 VPWR.n2068 VGND 0.00776f
C45034 VPWR.n2069 VGND 0.00655f
C45035 VPWR.n2070 VGND 0.00655f
C45036 VPWR.n2071 VGND 0.00698f
C45037 VPWR.n2072 VGND 0.00698f
C45038 VPWR.n2073 VGND 0.00655f
C45039 VPWR.n2074 VGND 0.00655f
C45040 VPWR.n2075 VGND 0.00813f
C45041 VPWR.n2076 VGND 0.00469f
C45042 VPWR.n2077 VGND 0.00655f
C45043 VPWR.n2078 VGND 0.00655f
C45044 VPWR.n2079 VGND 0.00515f
C45045 VPWR.n2080 VGND 0.01266f
C45046 VPWR.n2081 VGND 0.00735f
C45047 VPWR.n2082 VGND 0.00974f
C45048 VPWR.n2083 VGND 0.00761f
C45049 VPWR.n2084 VGND 0.01165f
C45050 VPWR.n2085 VGND 0.01144f
C45051 VPWR.n2086 VGND 0.02171f
C45052 VPWR.n2087 VGND 0.01577f
C45053 VPWR.n2088 VGND 0.0207f
C45054 VPWR.n2089 VGND 0.01577f
C45055 VPWR.n2090 VGND 0.0207f
C45056 VPWR.n2091 VGND 0.01762f
C45057 VPWR.n2092 VGND 0.01189f
C45058 VPWR.n2093 VGND 0.01144f
C45059 VPWR.n2094 VGND 0.01085f
C45060 VPWR.n2095 VGND 0.01085f
C45061 VPWR.n2096 VGND 0.0085f
C45062 VPWR.n2097 VGND 0.00813f
C45063 VPWR.n2098 VGND 0.0083f
C45064 VPWR.n2099 VGND 0.13412f
C45065 VPWR.n2100 VGND 0.13412f
C45066 VPWR.n2101 VGND 0.00656f
C45067 VPWR.n2102 VGND 0.00924f
C45068 VPWR.n2103 VGND 0.01085f
C45069 VPWR.n2104 VGND 0.01085f
C45070 VPWR.n2105 VGND 0.01085f
C45071 VPWR.n2106 VGND 0.01085f
C45072 VPWR.n2107 VGND 0.01144f
C45073 VPWR.n2108 VGND 0.01189f
C45074 VPWR.n2109 VGND 0.00758f
C45075 VPWR.n2110 VGND 0.00544f
C45076 VPWR.n2111 VGND 0.01023f
C45077 VPWR.n2112 VGND 0.01085f
C45078 VPWR.n2113 VGND 0.01085f
C45079 VPWR.n2114 VGND 0.01085f
C45080 VPWR.n2115 VGND 0.01085f
C45081 VPWR.n2116 VGND 0.01085f
C45082 VPWR.n2117 VGND 0.01085f
C45083 VPWR.n2118 VGND 0.01085f
C45084 VPWR.n2119 VGND 0.01085f
C45085 VPWR.n2120 VGND 0.01085f
C45086 VPWR.n2121 VGND 0.01085f
C45087 VPWR.n2122 VGND 0.01085f
C45088 VPWR.n2123 VGND 0.01085f
C45089 VPWR.n2124 VGND 0.01085f
C45090 VPWR.n2125 VGND 0.01144f
C45091 VPWR.n2126 VGND 0.01165f
C45092 VPWR.n2127 VGND 0.01568f
C45093 VPWR.n2128 VGND 0.02059f
C45094 VPWR.n2129 VGND 0.01588f
C45095 VPWR.n2130 VGND 0.02171f
C45096 VPWR.n2131 VGND 0.01855f
C45097 VPWR.n2132 VGND 0.00768f
C45098 VPWR.n2133 VGND 0.00515f
C45099 VPWR.n2134 VGND 0.0057f
C45100 VPWR.n2135 VGND 0.00761f
C45101 VPWR.n2136 VGND 0.00627f
C45102 VPWR.n2137 VGND 0.01023f
C45103 VPWR.n2138 VGND 0.00974f
C45104 VPWR.n2139 VGND 0.00735f
C45105 VPWR.n2140 VGND 0.01189f
C45106 VPWR.n2141 VGND 0.0085f
C45107 VPWR.n2142 VGND 0.00627f
C45108 VPWR.n2143 VGND 0.01023f
C45109 VPWR.n2144 VGND 0.01085f
C45110 VPWR.n2145 VGND 0.01085f
C45111 VPWR.n2146 VGND 0.01085f
C45112 VPWR.n2147 VGND 0.01085f
C45113 VPWR.n2148 VGND 0.01085f
C45114 VPWR.n2149 VGND 0.00985f
C45115 VPWR.n2150 VGND 0.01013f
C45116 VPWR.n2151 VGND 0.01085f
C45117 VPWR.n2152 VGND 0.01085f
C45118 VPWR.n2153 VGND 0.01085f
C45119 VPWR.n2154 VGND 0.01085f
C45120 VPWR.n2155 VGND 0.01085f
C45121 VPWR.n2156 VGND 0.01085f
C45122 VPWR.n2157 VGND 0.01144f
C45123 VPWR.t495 VGND 0.00433f
C45124 VPWR.t1550 VGND 0.00433f
C45125 VPWR.t3608 VGND 0.00433f
C45126 VPWR.t2662 VGND 0.00433f
C45127 VPWR.t5710 VGND 0.00433f
C45128 VPWR.t6283 VGND 0.00433f
C45129 VPWR.t4239 VGND 0.00433f
C45130 VPWR.t3547 VGND 0.00433f
C45131 VPWR.t3187 VGND 0.00433f
C45132 VPWR.n2158 VGND 0.01085f
C45133 VPWR.n2159 VGND 0.01085f
C45134 VPWR.n2160 VGND 0.01085f
C45135 VPWR.n2161 VGND 0.01085f
C45136 VPWR.n2162 VGND 0.01085f
C45137 VPWR.n2163 VGND 0.01085f
C45138 VPWR.n2164 VGND 0.01023f
C45139 VPWR.n2165 VGND 0.00544f
C45140 VPWR.n2166 VGND 0.00758f
C45141 VPWR.n2167 VGND 0.01189f
C45142 VPWR.t427 VGND 0.06143f
C45143 VPWR.t494 VGND 0.05001f
C45144 VPWR.t1549 VGND 0.0173f
C45145 VPWR.t3607 VGND 0.04521f
C45146 VPWR.t2661 VGND 0.05001f
C45147 VPWR.t5709 VGND 0.05001f
C45148 VPWR.t6282 VGND 0.05001f
C45149 VPWR.t4238 VGND 0.05001f
C45150 VPWR.t3546 VGND 0.05001f
C45151 VPWR.t3186 VGND 0.05001f
C45152 VPWR.t4353 VGND 0.05001f
C45153 VPWR.t4545 VGND 0.05001f
C45154 VPWR.t681 VGND 0.05001f
C45155 VPWR.t5724 VGND 0.05001f
C45156 VPWR.t1474 VGND 0.05001f
C45157 VPWR.t6159 VGND 0.05001f
C45158 VPWR.t4395 VGND 0.0298f
C45159 VPWR.t3617 VGND 0.04122f
C45160 VPWR.t4716 VGND 0.00433f
C45161 VPWR.t1225 VGND 0.00433f
C45162 VPWR.t4033 VGND 0.00433f
C45163 VPWR.t3567 VGND 0.00433f
C45164 VPWR.t1045 VGND 0.00433f
C45165 VPWR.t2713 VGND 0.00433f
C45166 VPWR.t5341 VGND 0.00433f
C45167 VPWR.t976 VGND 0.00433f
C45168 VPWR.t1837 VGND 0.00433f
C45169 VPWR.t349 VGND 0.00433f
C45170 VPWR.t2461 VGND 0.00433f
C45171 VPWR.t394 VGND 0.00433f
C45172 VPWR.t3227 VGND 0.00433f
C45173 VPWR.t3205 VGND 0.00433f
C45174 VPWR.t3038 VGND 0.00433f
C45175 VPWR.t5135 VGND 0.00433f
C45176 VPWR.t1224 VGND 0.08271f
C45177 VPWR.t3566 VGND 0.10001f
C45178 VPWR.t1044 VGND 0.10001f
C45179 VPWR.t975 VGND 0.10001f
C45180 VPWR.t348 VGND 0.10001f
C45181 VPWR.t393 VGND 0.10001f
C45182 VPWR.t3204 VGND 0.10001f
C45183 VPWR.t3037 VGND 0.06731f
C45184 VPWR.n2168 VGND 0.02233f
C45185 VPWR.n2169 VGND 0.02171f
C45186 VPWR.n2170 VGND 0.02171f
C45187 VPWR.n2171 VGND 0.01577f
C45188 VPWR.n2172 VGND 0.0207f
C45189 VPWR.n2173 VGND 0.02171f
C45190 VPWR.n2174 VGND 0.02171f
C45191 VPWR.n2175 VGND 0.01568f
C45192 VPWR.n2176 VGND 0.01165f
C45193 VPWR.n2177 VGND 0.01144f
C45194 VPWR.n2178 VGND 0.01085f
C45195 VPWR.n2179 VGND 0.01085f
C45196 VPWR.n2180 VGND 0.01085f
C45197 VPWR.n2181 VGND 0.01085f
C45198 VPWR.n2182 VGND 0.01085f
C45199 VPWR.n2183 VGND 0.00608f
C45200 VPWR.n2184 VGND 0.01004f
C45201 VPWR.n2185 VGND 0.13412f
C45202 VPWR.t1681 VGND 0.00433f
C45203 VPWR.n2186 VGND 0.01042f
C45204 VPWR.t4505 VGND 0.00433f
C45205 VPWR.t73 VGND 0.00433f
C45206 VPWR.t1287 VGND 0.00433f
C45207 VPWR.t6308 VGND 0.00433f
C45208 VPWR.t1410 VGND 0.00433f
C45209 VPWR.t6445 VGND 0.00433f
C45210 VPWR.t548 VGND 0.00433f
C45211 VPWR.t5556 VGND 0.00433f
C45212 VPWR.t3713 VGND 0.00433f
C45213 VPWR.t3538 VGND 0.00433f
C45214 VPWR.t534 VGND 0.00433f
C45215 VPWR.t2018 VGND 0.00433f
C45216 VPWR.t5944 VGND 0.00433f
C45217 VPWR.t4644 VGND 0.00433f
C45218 VPWR.t2452 VGND 0.00433f
C45219 VPWR.t808 VGND 0.00433f
C45220 VPWR.t680 VGND 0.00433f
C45221 VPWR.t1275 VGND 0.00433f
C45222 VPWR.t4921 VGND 0.00433f
C45223 VPWR.t1679 VGND 0.00433f
C45224 VPWR.t3195 VGND 0.00433f
C45225 VPWR.t1760 VGND 0.00433f
C45226 VPWR.t5995 VGND 0.00433f
C45227 VPWR.t5767 VGND 0.00433f
C45228 VPWR.t1417 VGND 0.05001f
C45229 VPWR.t2797 VGND 0.0173f
C45230 VPWR.t3176 VGND 0.04521f
C45231 VPWR.t7123 VGND 0.05001f
C45232 VPWR.t3466 VGND 0.05001f
C45233 VPWR.t3333 VGND 0.05001f
C45234 VPWR.t4806 VGND 0.05001f
C45235 VPWR.t4458 VGND 0.05001f
C45236 VPWR.t5359 VGND 0.05001f
C45237 VPWR.t4636 VGND 0.05001f
C45238 VPWR.t4594 VGND 0.05001f
C45239 VPWR.t2249 VGND 0.05001f
C45240 VPWR.t3035 VGND 0.05001f
C45241 VPWR.t2425 VGND 0.05001f
C45242 VPWR.t6085 VGND 0.05001f
C45243 VPWR.t2095 VGND 0.0298f
C45244 VPWR.t3712 VGND 0.0298f
C45245 VPWR.t3537 VGND 0.05001f
C45246 VPWR.t533 VGND 0.05001f
C45247 VPWR.t2017 VGND 0.05001f
C45248 VPWR.t5943 VGND 0.05001f
C45249 VPWR.t4643 VGND 0.05001f
C45250 VPWR.t2451 VGND 0.05001f
C45251 VPWR.t807 VGND 0.05001f
C45252 VPWR.t679 VGND 0.05001f
C45253 VPWR.t1274 VGND 0.05001f
C45254 VPWR.t4920 VGND 0.05001f
C45255 VPWR.t1678 VGND 0.05001f
C45256 VPWR.t3194 VGND 0.05001f
C45257 VPWR.t1759 VGND 0.04521f
C45258 VPWR.t5994 VGND 0.0173f
C45259 VPWR.t5766 VGND 0.05001f
C45260 VPWR.t1247 VGND 0.06143f
C45261 VPWR.t1248 VGND 0.00433f
C45262 VPWR.t2096 VGND 0.00433f
C45263 VPWR.t6086 VGND 0.00433f
C45264 VPWR.t2426 VGND 0.00433f
C45265 VPWR.t3036 VGND 0.00433f
C45266 VPWR.n2187 VGND 0.01085f
C45267 VPWR.n2188 VGND 0.01085f
C45268 VPWR.n2189 VGND 0.01085f
C45269 VPWR.n2190 VGND 0.01085f
C45270 VPWR.n2191 VGND 0.01144f
C45271 VPWR.n2192 VGND 0.01189f
C45272 VPWR.n2193 VGND 0.00758f
C45273 VPWR.n2194 VGND 0.00544f
C45274 VPWR.n2195 VGND 0.01023f
C45275 VPWR.n2196 VGND 0.01085f
C45276 VPWR.n2197 VGND 0.01085f
C45277 VPWR.n2198 VGND 0.01085f
C45278 VPWR.n2199 VGND 0.01085f
C45279 VPWR.n2200 VGND 0.01085f
C45280 VPWR.n2201 VGND 0.01085f
C45281 VPWR.n2202 VGND 0.01085f
C45282 VPWR.n2203 VGND 0.01085f
C45283 VPWR.n2204 VGND 0.01085f
C45284 VPWR.n2205 VGND 0.01085f
C45285 VPWR.n2206 VGND 0.01085f
C45286 VPWR.n2207 VGND 0.01085f
C45287 VPWR.n2208 VGND 0.01085f
C45288 VPWR.n2209 VGND 0.01144f
C45289 VPWR.t2474 VGND 0.00433f
C45290 VPWR.t3783 VGND 0.00433f
C45291 VPWR.t2300 VGND 0.00433f
C45292 VPWR.t5450 VGND 0.00433f
C45293 VPWR.t5606 VGND 0.00433f
C45294 VPWR.t5510 VGND 0.00433f
C45295 VPWR.t1184 VGND 0.00433f
C45296 VPWR.t3674 VGND 0.00433f
C45297 VPWR.t3444 VGND 0.00433f
C45298 VPWR.n2210 VGND 0.01085f
C45299 VPWR.n2211 VGND 0.01085f
C45300 VPWR.n2212 VGND 0.01085f
C45301 VPWR.n2213 VGND 0.01085f
C45302 VPWR.n2214 VGND 0.01085f
C45303 VPWR.n2215 VGND 0.01085f
C45304 VPWR.n2216 VGND 0.01023f
C45305 VPWR.n2217 VGND 0.00544f
C45306 VPWR.n2218 VGND 0.00758f
C45307 VPWR.n2219 VGND 0.01189f
C45308 VPWR.t5555 VGND 0.06143f
C45309 VPWR.t2473 VGND 0.05001f
C45310 VPWR.t3782 VGND 0.0173f
C45311 VPWR.t2299 VGND 0.04521f
C45312 VPWR.t5449 VGND 0.05001f
C45313 VPWR.t5605 VGND 0.05001f
C45314 VPWR.t5509 VGND 0.05001f
C45315 VPWR.t1183 VGND 0.05001f
C45316 VPWR.t3673 VGND 0.05001f
C45317 VPWR.t3443 VGND 0.05001f
C45318 VPWR.t1680 VGND 0.05001f
C45319 VPWR.t4504 VGND 0.05001f
C45320 VPWR.t72 VGND 0.05001f
C45321 VPWR.t1286 VGND 0.05001f
C45322 VPWR.t6307 VGND 0.05001f
C45323 VPWR.t1409 VGND 0.05001f
C45324 VPWR.t6444 VGND 0.0298f
C45325 VPWR.t547 VGND 0.04122f
C45326 VPWR.t4726 VGND 0.00433f
C45327 VPWR.t6127 VGND 0.00433f
C45328 VPWR.t5195 VGND 0.00433f
C45329 VPWR.t4170 VGND 0.00433f
C45330 VPWR.t1053 VGND 0.00433f
C45331 VPWR.t4878 VGND 0.00433f
C45332 VPWR.t4051 VGND 0.00433f
C45333 VPWR.t3382 VGND 0.00433f
C45334 VPWR.t1420 VGND 0.00433f
C45335 VPWR.t4129 VGND 0.00433f
C45336 VPWR.t2465 VGND 0.00433f
C45337 VPWR.t6450 VGND 0.00433f
C45338 VPWR.t3196 VGND 0.00433f
C45339 VPWR.t1227 VGND 0.00433f
C45340 VPWR.t3363 VGND 0.00433f
C45341 VPWR.t347 VGND 0.00433f
C45342 VPWR.t4725 VGND 0.08271f
C45343 VPWR.t4169 VGND 0.10001f
C45344 VPWR.t1052 VGND 0.10001f
C45345 VPWR.t3381 VGND 0.10001f
C45346 VPWR.t1419 VGND 0.10001f
C45347 VPWR.t2464 VGND 0.10001f
C45348 VPWR.t1226 VGND 0.10001f
C45349 VPWR.t346 VGND 0.06731f
C45350 VPWR.n2220 VGND 0.02233f
C45351 VPWR.n2221 VGND 0.02171f
C45352 VPWR.n2222 VGND 0.02171f
C45353 VPWR.n2223 VGND 0.01577f
C45354 VPWR.n2224 VGND 0.0207f
C45355 VPWR.n2225 VGND 0.02171f
C45356 VPWR.n2226 VGND 0.02171f
C45357 VPWR.n2227 VGND 0.01568f
C45358 VPWR.n2228 VGND 0.01165f
C45359 VPWR.n2229 VGND 0.01144f
C45360 VPWR.n2230 VGND 0.01085f
C45361 VPWR.n2231 VGND 0.01085f
C45362 VPWR.n2232 VGND 0.01085f
C45363 VPWR.n2233 VGND 0.01085f
C45364 VPWR.n2234 VGND 0.01085f
C45365 VPWR.n2235 VGND 0.00608f
C45366 VPWR.n2236 VGND 0.01004f
C45367 VPWR.n2237 VGND 0.13412f
C45368 VPWR.n2238 VGND 0.13412f
C45369 VPWR.n2239 VGND 0.01004f
C45370 VPWR.n2240 VGND 0.01042f
C45371 VPWR.n2241 VGND 0.01085f
C45372 VPWR.n2242 VGND 0.01085f
C45373 VPWR.n2243 VGND 0.01085f
C45374 VPWR.n2244 VGND 0.01085f
C45375 VPWR.n2245 VGND 0.01085f
C45376 VPWR.n2246 VGND 0.01085f
C45377 VPWR.n2247 VGND 0.01023f
C45378 VPWR.n2248 VGND 0.00544f
C45379 VPWR.n2249 VGND 0.00758f
C45380 VPWR.n2250 VGND 0.01189f
C45381 VPWR.n2251 VGND 0.01144f
C45382 VPWR.n2252 VGND 0.01085f
C45383 VPWR.n2253 VGND 0.01085f
C45384 VPWR.n2254 VGND 0.01085f
C45385 VPWR.n2255 VGND 0.01085f
C45386 VPWR.n2256 VGND 0.01085f
C45387 VPWR.n2257 VGND 0.01085f
C45388 VPWR.n2258 VGND 0.01085f
C45389 VPWR.n2259 VGND 0.01085f
C45390 VPWR.n2260 VGND 0.01085f
C45391 VPWR.n2261 VGND 0.01085f
C45392 VPWR.n2262 VGND 0.01085f
C45393 VPWR.n2263 VGND 0.01085f
C45394 VPWR.n2264 VGND 0.01085f
C45395 VPWR.n2265 VGND 0.01023f
C45396 VPWR.n2266 VGND 0.00544f
C45397 VPWR.n2267 VGND 0.00758f
C45398 VPWR.n2268 VGND 0.01189f
C45399 VPWR.n2269 VGND 0.01144f
C45400 VPWR.n2270 VGND 0.01085f
C45401 VPWR.n2271 VGND 0.01085f
C45402 VPWR.n2272 VGND 0.01085f
C45403 VPWR.n2273 VGND 0.01085f
C45404 VPWR.n2274 VGND 0.01027f
C45405 VPWR.n2275 VGND 0.00656f
C45406 VPWR.n2276 VGND 0.13412f
C45407 VPWR.n2277 VGND 0.13412f
C45408 VPWR.n2278 VGND 0.00656f
C45409 VPWR.n2279 VGND 0.00971f
C45410 VPWR.n2280 VGND 0.01085f
C45411 VPWR.n2281 VGND 0.01085f
C45412 VPWR.n2282 VGND 0.01085f
C45413 VPWR.n2283 VGND 0.01085f
C45414 VPWR.n2284 VGND 0.01085f
C45415 VPWR.n2285 VGND 0.01085f
C45416 VPWR.n2286 VGND 0.01085f
C45417 VPWR.n2287 VGND 0.01023f
C45418 VPWR.n2288 VGND 0.00544f
C45419 VPWR.n2289 VGND 0.00758f
C45420 VPWR.n2290 VGND 0.01189f
C45421 VPWR.n2291 VGND 0.01144f
C45422 VPWR.n2292 VGND 0.01085f
C45423 VPWR.n2293 VGND 0.01085f
C45424 VPWR.n2294 VGND 0.01085f
C45425 VPWR.n2295 VGND 0.01085f
C45426 VPWR.n2296 VGND 0.01085f
C45427 VPWR.n2297 VGND 0.01085f
C45428 VPWR.n2298 VGND 0.01085f
C45429 VPWR.n2299 VGND 0.01085f
C45430 VPWR.n2300 VGND 0.01085f
C45431 VPWR.n2301 VGND 0.01085f
C45432 VPWR.n2302 VGND 0.01085f
C45433 VPWR.n2303 VGND 0.01085f
C45434 VPWR.n2304 VGND 0.01085f
C45435 VPWR.n2305 VGND 0.01023f
C45436 VPWR.n2306 VGND 0.00544f
C45437 VPWR.n2307 VGND 0.00758f
C45438 VPWR.n2308 VGND 0.01189f
C45439 VPWR.n2309 VGND 0.01144f
C45440 VPWR.n2310 VGND 0.01085f
C45441 VPWR.n2311 VGND 0.01085f
C45442 VPWR.n2312 VGND 0.01085f
C45443 VPWR.n2313 VGND 0.01085f
C45444 VPWR.n2314 VGND 0.00924f
C45445 VPWR.n2315 VGND 0.00656f
C45446 VPWR.n2316 VGND 0.13412f
C45447 VPWR.t5987 VGND 0.00433f
C45448 VPWR.t884 VGND 0.00433f
C45449 VPWR.n2317 VGND 0.01985f
C45450 VPWR.t990 VGND 0.00433f
C45451 VPWR.t5181 VGND 0.00433f
C45452 VPWR.t1343 VGND 0.00433f
C45453 VPWR.t4266 VGND 0.00433f
C45454 VPWR.t3968 VGND 0.00433f
C45455 VPWR.t4754 VGND 0.00433f
C45456 VPWR.t5646 VGND 0.00433f
C45457 VPWR.t5078 VGND 0.00433f
C45458 VPWR.n2318 VGND 0.02392f
C45459 VPWR.n2319 VGND 0.01074f
C45460 VPWR.t4011 VGND 0.00433f
C45461 VPWR.t4304 VGND 0.00433f
C45462 VPWR.t1580 VGND 0.00433f
C45463 VPWR.t5098 VGND 0.00433f
C45464 VPWR.t1896 VGND 0.00433f
C45465 VPWR.t579 VGND 0.00433f
C45466 VPWR.n2320 VGND 0.02171f
C45467 VPWR.n2321 VGND 0.02171f
C45468 VPWR.n2322 VGND 0.01673f
C45469 VPWR.n2323 VGND 0.00992f
C45470 VPWR.n2324 VGND 0.02102f
C45471 VPWR.t4010 VGND 0.08271f
C45472 VPWR.t1579 VGND 0.10001f
C45473 VPWR.t578 VGND 0.10001f
C45474 VPWR.t883 VGND 0.10001f
C45475 VPWR.t989 VGND 0.10001f
C45476 VPWR.t1342 VGND 0.10001f
C45477 VPWR.t3967 VGND 0.10001f
C45478 VPWR.t5077 VGND 0.06731f
C45479 VPWR.n2325 VGND 0.02437f
C45480 VPWR.n2326 VGND 0.04223f
C45481 VPWR.t692 VGND 0.00433f
C45482 VPWR.t2856 VGND 0.00433f
C45483 VPWR.t4407 VGND 0.00433f
C45484 VPWR.t1578 VGND 0.00433f
C45485 VPWR.t3794 VGND 0.00433f
C45486 VPWR.t5083 VGND 0.00433f
C45487 VPWR.t5581 VGND 0.00433f
C45488 VPWR.t5812 VGND 0.00433f
C45489 VPWR.t691 VGND 0.05334f
C45490 VPWR.t2855 VGND 0.05996f
C45491 VPWR.t4406 VGND 0.05996f
C45492 VPWR.t1577 VGND 0.05996f
C45493 VPWR.t3793 VGND 0.05996f
C45494 VPWR.t5082 VGND 0.05996f
C45495 VPWR.t5580 VGND 0.05996f
C45496 VPWR.t5811 VGND 0.04035f
C45497 VPWR.n2327 VGND 0.03832f
C45498 VPWR.t4377 VGND 0.00433f
C45499 VPWR.t552 VGND 0.00433f
C45500 VPWR.t1349 VGND 0.00433f
C45501 VPWR.t2088 VGND 0.00433f
C45502 VPWR.t4860 VGND 0.00433f
C45503 VPWR.t1546 VGND 0.00433f
C45504 VPWR.t447 VGND 0.00433f
C45505 VPWR.t3522 VGND 0.00433f
C45506 VPWR.t4376 VGND 0.05247f
C45507 VPWR.t551 VGND 0.05996f
C45508 VPWR.t1348 VGND 0.05996f
C45509 VPWR.t2087 VGND 0.05996f
C45510 VPWR.t4859 VGND 0.05996f
C45511 VPWR.t1545 VGND 0.05996f
C45512 VPWR.t446 VGND 0.05996f
C45513 VPWR.t3521 VGND 0.04035f
C45514 VPWR.n2328 VGND 0.03832f
C45515 VPWR.t1094 VGND 0.00433f
C45516 VPWR.t4078 VGND 0.00433f
C45517 VPWR.t4976 VGND 0.00433f
C45518 VPWR.t5375 VGND 0.00433f
C45519 VPWR.t5787 VGND 0.00433f
C45520 VPWR.t6122 VGND 0.00433f
C45521 VPWR.t1498 VGND 0.00433f
C45522 VPWR.t3939 VGND 0.00433f
C45523 VPWR.t1093 VGND 0.05247f
C45524 VPWR.t4077 VGND 0.05996f
C45525 VPWR.t4975 VGND 0.05996f
C45526 VPWR.t5374 VGND 0.05996f
C45527 VPWR.t5786 VGND 0.05996f
C45528 VPWR.t6121 VGND 0.05996f
C45529 VPWR.t1497 VGND 0.05996f
C45530 VPWR.t3938 VGND 0.04035f
C45531 VPWR.n2329 VGND 0.03832f
C45532 VPWR.t1939 VGND 0.00433f
C45533 VPWR.t5066 VGND 0.00433f
C45534 VPWR.t5649 VGND 0.00433f
C45535 VPWR.t1803 VGND 0.00433f
C45536 VPWR.t3294 VGND 0.00433f
C45537 VPWR.t6237 VGND 0.00433f
C45538 VPWR.t6273 VGND 0.00433f
C45539 VPWR.t4364 VGND 0.00433f
C45540 VPWR.t1938 VGND 0.05247f
C45541 VPWR.t5065 VGND 0.05996f
C45542 VPWR.t5648 VGND 0.05996f
C45543 VPWR.t1802 VGND 0.05996f
C45544 VPWR.t3293 VGND 0.05996f
C45545 VPWR.t6236 VGND 0.05996f
C45546 VPWR.t6272 VGND 0.05996f
C45547 VPWR.t4363 VGND 0.04035f
C45548 VPWR.n2330 VGND 0.03832f
C45549 VPWR.t5715 VGND 0.00433f
C45550 VPWR.t2460 VGND 0.00433f
C45551 VPWR.t5839 VGND 0.00433f
C45552 VPWR.t5280 VGND 0.00433f
C45553 VPWR.t2693 VGND 0.00433f
C45554 VPWR.t6051 VGND 0.00433f
C45555 VPWR.t5286 VGND 0.00433f
C45556 VPWR.t1830 VGND 0.00433f
C45557 VPWR.t5714 VGND 0.05247f
C45558 VPWR.t2459 VGND 0.05996f
C45559 VPWR.t5838 VGND 0.05996f
C45560 VPWR.t5279 VGND 0.05996f
C45561 VPWR.t2692 VGND 0.05996f
C45562 VPWR.t6050 VGND 0.05996f
C45563 VPWR.t5285 VGND 0.05996f
C45564 VPWR.t1829 VGND 0.04035f
C45565 VPWR.n2331 VGND 0.01842f
C45566 VPWR.n2332 VGND 0.0178f
C45567 VPWR.n2333 VGND 0.0178f
C45568 VPWR.n2334 VGND 0.01186f
C45569 VPWR.n2335 VGND 0.01679f
C45570 VPWR.n2336 VGND 0.0178f
C45571 VPWR.n2337 VGND 0.0178f
C45572 VPWR.n2338 VGND 0.01371f
C45573 VPWR.n2339 VGND 0.01189f
C45574 VPWR.n2340 VGND 0.01839f
C45575 VPWR.n2341 VGND 0.0178f
C45576 VPWR.n2342 VGND 0.01476f
C45577 VPWR.n2343 VGND 0.01177f
C45578 VPWR.n2344 VGND 0.00795f
C45579 VPWR.n2345 VGND 0.01679f
C45580 VPWR.n2346 VGND 0.0178f
C45581 VPWR.n2347 VGND 0.0178f
C45582 VPWR.n2348 VGND 0.01371f
C45583 VPWR.n2349 VGND 0.01189f
C45584 VPWR.n2350 VGND 0.01839f
C45585 VPWR.n2351 VGND 0.0178f
C45586 VPWR.n2352 VGND 0.0178f
C45587 VPWR.n2353 VGND 0.01186f
C45588 VPWR.n2354 VGND 0.01679f
C45589 VPWR.n2355 VGND 0.0178f
C45590 VPWR.n2356 VGND 0.0178f
C45591 VPWR.n2357 VGND 0.01371f
C45592 VPWR.n2358 VGND 0.01189f
C45593 VPWR.n2359 VGND 0.01839f
C45594 VPWR.n2360 VGND 0.0178f
C45595 VPWR.n2361 VGND 0.01721f
C45596 VPWR.n2362 VGND 0.01177f
C45597 VPWR.n2363 VGND 0.00551f
C45598 VPWR.n2364 VGND 0.01679f
C45599 VPWR.n2365 VGND 0.0178f
C45600 VPWR.n2366 VGND 0.0178f
C45601 VPWR.n2367 VGND 0.01371f
C45602 VPWR.n2368 VGND 0.01189f
C45603 VPWR.n2369 VGND 0.01839f
C45604 VPWR.n2370 VGND 0.0178f
C45605 VPWR.n2371 VGND 0.0178f
C45606 VPWR.n2372 VGND 0.01186f
C45607 VPWR.n2373 VGND 0.01679f
C45608 VPWR.n2374 VGND 0.0178f
C45609 VPWR.n2375 VGND 0.0178f
C45610 VPWR.n2376 VGND 0.01364f
C45611 VPWR.n2377 VGND 0.01156f
C45612 VPWR.n2378 VGND 0.0223f
C45613 VPWR.n2379 VGND 0.02171f
C45614 VPWR.n2380 VGND 0.02171f
C45615 VPWR.n2381 VGND 0.01577f
C45616 VPWR.n2382 VGND 0.01076f
C45617 VPWR.n2383 VGND 0.13412f
C45618 VPWR.t4371 VGND 0.00433f
C45619 VPWR.t1616 VGND 0.00433f
C45620 VPWR.n2384 VGND 0.01985f
C45621 VPWR.t5820 VGND 0.00433f
C45622 VPWR.t6441 VGND 0.00433f
C45623 VPWR.t3455 VGND 0.00433f
C45624 VPWR.t7114 VGND 0.00433f
C45625 VPWR.t3433 VGND 0.00433f
C45626 VPWR.t6238 VGND 0.00433f
C45627 VPWR.t2341 VGND 0.00433f
C45628 VPWR.t5837 VGND 0.00433f
C45629 VPWR.t6202 VGND 0.00433f
C45630 VPWR.n2385 VGND 0.0072f
C45631 VPWR.t3234 VGND 0.00433f
C45632 VPWR.t1402 VGND 0.00433f
C45633 VPWR.t5035 VGND 0.00433f
C45634 VPWR.t5677 VGND 0.00433f
C45635 VPWR.t4827 VGND 0.00433f
C45636 VPWR.t2732 VGND 0.00433f
C45637 VPWR.n2386 VGND 0.02171f
C45638 VPWR.n2387 VGND 0.02171f
C45639 VPWR.n2388 VGND 0.01673f
C45640 VPWR.t6201 VGND 0.04122f
C45641 VPWR.t1401 VGND 0.08271f
C45642 VPWR.t5034 VGND 0.10001f
C45643 VPWR.t2731 VGND 0.10001f
C45644 VPWR.t1615 VGND 0.10001f
C45645 VPWR.t5819 VGND 0.10001f
C45646 VPWR.t3454 VGND 0.10001f
C45647 VPWR.t3432 VGND 0.10001f
C45648 VPWR.t2340 VGND 0.06731f
C45649 VPWR.n2389 VGND 0.02233f
C45650 VPWR.n2390 VGND 0.02171f
C45651 VPWR.n2391 VGND 0.02171f
C45652 VPWR.n2392 VGND 0.01577f
C45653 VPWR.n2393 VGND 0.01076f
C45654 VPWR.n2394 VGND 0.13412f
C45655 VPWR.t6186 VGND 0.00433f
C45656 VPWR.t1209 VGND 0.00433f
C45657 VPWR.n2395 VGND 0.01985f
C45658 VPWR.t3690 VGND 0.00433f
C45659 VPWR.t5182 VGND 0.00433f
C45660 VPWR.t3103 VGND 0.00433f
C45661 VPWR.t3513 VGND 0.00433f
C45662 VPWR.t2840 VGND 0.00433f
C45663 VPWR.t4757 VGND 0.00433f
C45664 VPWR.t6113 VGND 0.00433f
C45665 VPWR.t5307 VGND 0.00433f
C45666 VPWR.t3524 VGND 0.00433f
C45667 VPWR.n2396 VGND 0.0072f
C45668 VPWR.t4214 VGND 0.00433f
C45669 VPWR.t4445 VGND 0.00433f
C45670 VPWR.t996 VGND 0.00433f
C45671 VPWR.t3539 VGND 0.00433f
C45672 VPWR.t5506 VGND 0.00433f
C45673 VPWR.t6020 VGND 0.00433f
C45674 VPWR.n2397 VGND 0.02171f
C45675 VPWR.n2398 VGND 0.02171f
C45676 VPWR.n2399 VGND 0.01673f
C45677 VPWR.t3523 VGND 0.04122f
C45678 VPWR.t4213 VGND 0.08271f
C45679 VPWR.t995 VGND 0.10001f
C45680 VPWR.t5505 VGND 0.10001f
C45681 VPWR.t1208 VGND 0.10001f
C45682 VPWR.t3689 VGND 0.10001f
C45683 VPWR.t3102 VGND 0.10001f
C45684 VPWR.t2839 VGND 0.10001f
C45685 VPWR.t5306 VGND 0.06731f
C45686 VPWR.n2400 VGND 0.02233f
C45687 VPWR.n2401 VGND 0.02171f
C45688 VPWR.n2402 VGND 0.02171f
C45689 VPWR.n2403 VGND 0.01577f
C45690 VPWR.n2404 VGND 0.01076f
C45691 VPWR.n2405 VGND 0.13412f
C45692 VPWR.t892 VGND 0.00433f
C45693 VPWR.t2780 VGND 0.00433f
C45694 VPWR.n2406 VGND 0.01985f
C45695 VPWR.t998 VGND 0.00433f
C45696 VPWR.t5993 VGND 0.00433f
C45697 VPWR.t3248 VGND 0.00433f
C45698 VPWR.t678 VGND 0.00433f
C45699 VPWR.t6181 VGND 0.00433f
C45700 VPWR.t3117 VGND 0.00433f
C45701 VPWR.t2929 VGND 0.00433f
C45702 VPWR.t2496 VGND 0.00433f
C45703 VPWR.t3643 VGND 0.00433f
C45704 VPWR.n2407 VGND 0.0072f
C45705 VPWR.t4741 VGND 0.00433f
C45706 VPWR.t3378 VGND 0.00433f
C45707 VPWR.t4055 VGND 0.00433f
C45708 VPWR.t6136 VGND 0.00433f
C45709 VPWR.t3437 VGND 0.00433f
C45710 VPWR.t3858 VGND 0.00433f
C45711 VPWR.n2408 VGND 0.02171f
C45712 VPWR.n2409 VGND 0.02171f
C45713 VPWR.n2410 VGND 0.01673f
C45714 VPWR.t3642 VGND 0.04122f
C45715 VPWR.t3377 VGND 0.08271f
C45716 VPWR.t4054 VGND 0.10001f
C45717 VPWR.t3436 VGND 0.10001f
C45718 VPWR.t891 VGND 0.10001f
C45719 VPWR.t997 VGND 0.10001f
C45720 VPWR.t677 VGND 0.10001f
C45721 VPWR.t3116 VGND 0.10001f
C45722 VPWR.t2495 VGND 0.06731f
C45723 VPWR.n2411 VGND 0.02233f
C45724 VPWR.n2412 VGND 0.02171f
C45725 VPWR.n2413 VGND 0.02171f
C45726 VPWR.n2414 VGND 0.01577f
C45727 VPWR.n2415 VGND 0.01076f
C45728 VPWR.n2416 VGND 0.13412f
C45729 VPWR.t5968 VGND 0.00433f
C45730 VPWR.n2417 VGND 0.00899f
C45731 VPWR.t5762 VGND 0.00433f
C45732 VPWR.t840 VGND 0.00433f
C45733 VPWR.t4489 VGND 0.00433f
C45734 VPWR.t2199 VGND 0.00433f
C45735 VPWR.t2116 VGND 0.00433f
C45736 VPWR.t1754 VGND 0.00433f
C45737 VPWR.t2813 VGND 0.00433f
C45738 VPWR.t834 VGND 0.00433f
C45739 VPWR.t712 VGND 0.00433f
C45740 VPWR.t378 VGND 0.00433f
C45741 VPWR.t4553 VGND 0.00433f
C45742 VPWR.n2418 VGND 0.0085f
C45743 VPWR.n2419 VGND 0.00974f
C45744 VPWR.n2420 VGND 0.01085f
C45745 VPWR.n2421 VGND 0.01085f
C45746 VPWR.n2422 VGND 0.01085f
C45747 VPWR.n2423 VGND 0.0085f
C45748 VPWR.n2424 VGND 0.00738f
C45749 VPWR.n2425 VGND 0.00896f
C45750 VPWR.n2426 VGND 0.00665f
C45751 VPWR.t4488 VGND 0.03271f
C45752 VPWR.t2198 VGND 0.05001f
C45753 VPWR.t2115 VGND 0.04231f
C45754 VPWR.t1753 VGND 0.025f
C45755 VPWR.t2812 VGND 0.03271f
C45756 VPWR.t833 VGND 0.05001f
C45757 VPWR.t711 VGND 0.05001f
C45758 VPWR.t377 VGND 0.05001f
C45759 VPWR.t4552 VGND 0.05001f
C45760 VPWR.t5967 VGND 0.05001f
C45761 VPWR.t5761 VGND 0.04231f
C45762 VPWR.t839 VGND 0.0202f
C45763 VPWR.n2427 VGND 0.05372f
C45764 VPWR.t5362 VGND 0.00433f
C45765 VPWR.t6120 VGND 0.00433f
C45766 VPWR.t1098 VGND 0.00433f
C45767 VPWR.t4102 VGND 0.00433f
C45768 VPWR.t1010 VGND 0.00433f
C45769 VPWR.t1341 VGND 0.00433f
C45770 VPWR.t1283 VGND 0.00433f
C45771 VPWR.t4945 VGND 0.00433f
C45772 VPWR.t4772 VGND 0.00433f
C45773 VPWR.t5361 VGND 0.08751f
C45774 VPWR.t1097 VGND 0.10001f
C45775 VPWR.t1009 VGND 0.10001f
C45776 VPWR.t1282 VGND 0.06731f
C45777 VPWR.n2428 VGND 0.03642f
C45778 VPWR.t855 VGND 0.00433f
C45779 VPWR.t4176 VGND 0.00433f
C45780 VPWR.t769 VGND 0.00433f
C45781 VPWR.t2063 VGND 0.00433f
C45782 VPWR.t3655 VGND 0.00433f
C45783 VPWR.t3084 VGND 0.00433f
C45784 VPWR.t4784 VGND 0.00433f
C45785 VPWR.t4771 VGND 0.03751f
C45786 VPWR.t854 VGND 0.04231f
C45787 VPWR.t4175 VGND 0.03271f
C45788 VPWR.t768 VGND 0.05001f
C45789 VPWR.t2062 VGND 0.05001f
C45790 VPWR.t3654 VGND 0.05001f
C45791 VPWR.t3083 VGND 0.04231f
C45792 VPWR.t4783 VGND 0.0202f
C45793 VPWR.t914 VGND 0.06731f
C45794 VPWR.t456 VGND 0.10001f
C45795 VPWR.t762 VGND 0.10001f
C45796 VPWR.t1065 VGND 0.10001f
C45797 VPWR.t2551 VGND 0.10001f
C45798 VPWR.t821 VGND 0.10001f
C45799 VPWR.t1771 VGND 0.10001f
C45800 VPWR.t2099 VGND 0.08751f
C45801 VPWR.n2429 VGND 0.05372f
C45802 VPWR.t2100 VGND 0.00433f
C45803 VPWR.t6012 VGND 0.00433f
C45804 VPWR.t1772 VGND 0.00433f
C45805 VPWR.t2566 VGND 0.00433f
C45806 VPWR.t822 VGND 0.00433f
C45807 VPWR.t5081 VGND 0.00433f
C45808 VPWR.t4475 VGND 0.00433f
C45809 VPWR.t2552 VGND 0.00433f
C45810 VPWR.t1066 VGND 0.00433f
C45811 VPWR.t4487 VGND 0.00433f
C45812 VPWR.t763 VGND 0.00433f
C45813 VPWR.t5500 VGND 0.00433f
C45814 VPWR.t457 VGND 0.00433f
C45815 VPWR.t5200 VGND 0.00433f
C45816 VPWR.n2430 VGND 0.02171f
C45817 VPWR.n2431 VGND 0.01568f
C45818 VPWR.n2432 VGND 0.01486f
C45819 VPWR.n2433 VGND 0.0207f
C45820 VPWR.n2434 VGND 0.02171f
C45821 VPWR.n2435 VGND 0.02171f
C45822 VPWR.n2436 VGND 0.01762f
C45823 VPWR.n2437 VGND 0.01189f
C45824 VPWR.n2438 VGND 0.01144f
C45825 VPWR.n2439 VGND 0.01085f
C45826 VPWR.n2440 VGND 0.01085f
C45827 VPWR.n2441 VGND 0.01085f
C45828 VPWR.n2442 VGND 0.01085f
C45829 VPWR.n2443 VGND 0.0085f
C45830 VPWR.n2444 VGND 0.00912f
C45831 VPWR.n2445 VGND 0.01189f
C45832 VPWR.n2446 VGND 0.00551f
C45833 VPWR.n2447 VGND 0.0207f
C45834 VPWR.n2448 VGND 0.02171f
C45835 VPWR.n2449 VGND 0.02171f
C45836 VPWR.n2450 VGND 0.01577f
C45837 VPWR.n2451 VGND 0.01088f
C45838 VPWR.n2452 VGND 0.01144f
C45839 VPWR.n2453 VGND 0.00924f
C45840 VPWR.n2454 VGND 0.0083f
C45841 VPWR.n2455 VGND 0.10419f
C45842 VPWR.n2456 VGND 0.13412f
C45843 VPWR.n2457 VGND 0.01076f
C45844 VPWR.n2458 VGND 0.01577f
C45845 VPWR.n2459 VGND 0.01144f
C45846 VPWR.n2460 VGND 0.01189f
C45847 VPWR.n2461 VGND 0.01023f
C45848 VPWR.n2462 VGND 0.01085f
C45849 VPWR.n2463 VGND 0.01085f
C45850 VPWR.n2464 VGND 0.01085f
C45851 VPWR.n2465 VGND 0.01147f
C45852 VPWR.n2466 VGND 0.01156f
C45853 VPWR.n2467 VGND 0.01264f
C45854 VPWR.n2468 VGND 0.01186f
C45855 VPWR.n2469 VGND 0.0178f
C45856 VPWR.n2470 VGND 0.0178f
C45857 VPWR.n2471 VGND 0.01839f
C45858 VPWR.t988 VGND 0.00433f
C45859 VPWR.t4953 VGND 0.00433f
C45860 VPWR.t7120 VGND 0.00433f
C45861 VPWR.t4624 VGND 0.00433f
C45862 VPWR.t5860 VGND 0.00433f
C45863 VPWR.t1440 VGND 0.00433f
C45864 VPWR.t626 VGND 0.00433f
C45865 VPWR.n2472 VGND 0.0178f
C45866 VPWR.n2473 VGND 0.0178f
C45867 VPWR.n2474 VGND 0.01186f
C45868 VPWR.n2475 VGND 0.01679f
C45869 VPWR.n2476 VGND 0.0178f
C45870 VPWR.n2477 VGND 0.0178f
C45871 VPWR.n2478 VGND 0.01371f
C45872 VPWR.n2479 VGND 0.01189f
C45873 VPWR.n2480 VGND 0.03832f
C45874 VPWR.t987 VGND 0.05247f
C45875 VPWR.t4952 VGND 0.05996f
C45876 VPWR.t7119 VGND 0.05996f
C45877 VPWR.t4623 VGND 0.05996f
C45878 VPWR.t5859 VGND 0.05996f
C45879 VPWR.t1439 VGND 0.05996f
C45880 VPWR.t625 VGND 0.05996f
C45881 VPWR.t867 VGND 0.04035f
C45882 VPWR.n2481 VGND 0.03832f
C45883 VPWR.t4373 VGND 0.00433f
C45884 VPWR.t1309 VGND 0.00433f
C45885 VPWR.t1240 VGND 0.00433f
C45886 VPWR.t4453 VGND 0.00433f
C45887 VPWR.t2928 VGND 0.00433f
C45888 VPWR.t5199 VGND 0.00433f
C45889 VPWR.t453 VGND 0.00433f
C45890 VPWR.t5171 VGND 0.00433f
C45891 VPWR.t4372 VGND 0.05247f
C45892 VPWR.t1308 VGND 0.05996f
C45893 VPWR.t1239 VGND 0.05996f
C45894 VPWR.t4452 VGND 0.05996f
C45895 VPWR.t2927 VGND 0.05996f
C45896 VPWR.t5198 VGND 0.05996f
C45897 VPWR.t452 VGND 0.05996f
C45898 VPWR.t5170 VGND 0.04035f
C45899 VPWR.t6322 VGND 0.04035f
C45900 VPWR.t2748 VGND 0.05996f
C45901 VPWR.t2934 VGND 0.05996f
C45902 VPWR.t1038 VGND 0.05996f
C45903 VPWR.t2696 VGND 0.05996f
C45904 VPWR.t5893 VGND 0.05996f
C45905 VPWR.t3738 VGND 0.05996f
C45906 VPWR.t4657 VGND 0.05247f
C45907 VPWR.n2482 VGND 0.03832f
C45908 VPWR.t4658 VGND 0.00433f
C45909 VPWR.t3739 VGND 0.00433f
C45910 VPWR.t5894 VGND 0.00433f
C45911 VPWR.t2697 VGND 0.00433f
C45912 VPWR.t1039 VGND 0.00433f
C45913 VPWR.t2935 VGND 0.00433f
C45914 VPWR.t2749 VGND 0.00433f
C45915 VPWR.n2483 VGND 0.0178f
C45916 VPWR.n2484 VGND 0.0178f
C45917 VPWR.n2485 VGND 0.01186f
C45918 VPWR.n2486 VGND 0.01679f
C45919 VPWR.n2487 VGND 0.0178f
C45920 VPWR.n2488 VGND 0.0178f
C45921 VPWR.n2489 VGND 0.01371f
C45922 VPWR.n2490 VGND 0.01189f
C45923 VPWR.n2491 VGND 0.01839f
C45924 VPWR.n2492 VGND 0.0178f
C45925 VPWR.n2493 VGND 0.0178f
C45926 VPWR.n2494 VGND 0.01186f
C45927 VPWR.n2495 VGND 0.01679f
C45928 VPWR.n2496 VGND 0.0178f
C45929 VPWR.n2497 VGND 0.0178f
C45930 VPWR.n2498 VGND 0.01371f
C45931 VPWR.n2499 VGND 0.01189f
C45932 VPWR.n2500 VGND 0.01236f
C45933 VPWR.n2501 VGND 0.32859f
C45934 VPWR.n2502 VGND 0.10419f
C45935 VPWR.n2503 VGND 0.01177f
C45936 VPWR.n2504 VGND 0.01085f
C45937 VPWR.n2505 VGND 0.01189f
C45938 VPWR.n2506 VGND 0.01023f
C45939 VPWR.n2507 VGND 0.01085f
C45940 VPWR.n2508 VGND 0.01085f
C45941 VPWR.n2509 VGND 0.01085f
C45942 VPWR.n2510 VGND 0.01085f
C45943 VPWR.n2511 VGND 0.01085f
C45944 VPWR.n2512 VGND 0.01085f
C45945 VPWR.n2513 VGND 0.00985f
C45946 VPWR.n2514 VGND 0.00898f
C45947 VPWR.n2515 VGND 0.01189f
C45948 VPWR.n2516 VGND 0.01303f
C45949 VPWR.n2517 VGND 0.01935f
C45950 VPWR.n2518 VGND 0.02171f
C45951 VPWR.n2519 VGND 0.01144f
C45952 VPWR.t6204 VGND 0.00433f
C45953 VPWR.t2055 VGND 0.00433f
C45954 VPWR.t4763 VGND 0.00433f
C45955 VPWR.t6251 VGND 0.00433f
C45956 VPWR.t5830 VGND 0.00433f
C45957 VPWR.t3165 VGND 0.00433f
C45958 VPWR.t6093 VGND 0.00433f
C45959 VPWR.t4913 VGND 0.00433f
C45960 VPWR.t2613 VGND 0.00433f
C45961 VPWR.t3877 VGND 0.00433f
C45962 VPWR.t3875 VGND 0.00433f
C45963 VPWR.t4021 VGND 0.00433f
C45964 VPWR.t5867 VGND 0.00433f
C45965 VPWR.t4639 VGND 0.00433f
C45966 VPWR.n2520 VGND 0.01085f
C45967 VPWR.n2521 VGND 0.01085f
C45968 VPWR.n2522 VGND 0.0083f
C45969 VPWR.n2523 VGND 0.00994f
C45970 VPWR.n2524 VGND 0.01085f
C45971 VPWR.n2525 VGND 0.00839f
C45972 VPWR.n2526 VGND 0.00985f
C45973 VPWR.n2527 VGND 0.01085f
C45974 VPWR.n2528 VGND 0.01085f
C45975 VPWR.n2529 VGND 0.01085f
C45976 VPWR.n2530 VGND 0.01085f
C45977 VPWR.n2531 VGND 0.01085f
C45978 VPWR.n2532 VGND 0.01085f
C45979 VPWR.n2533 VGND 0.01023f
C45980 VPWR.n2534 VGND 0.01189f
C45981 VPWR.n2535 VGND 0.03642f
C45982 VPWR.t1779 VGND 0.03751f
C45983 VPWR.t6203 VGND 0.05001f
C45984 VPWR.t2054 VGND 0.05001f
C45985 VPWR.t4762 VGND 0.05001f
C45986 VPWR.t6250 VGND 0.05001f
C45987 VPWR.t5829 VGND 0.05001f
C45988 VPWR.t3164 VGND 0.05001f
C45989 VPWR.t6092 VGND 0.05001f
C45990 VPWR.t4912 VGND 0.05001f
C45991 VPWR.t2612 VGND 0.05001f
C45992 VPWR.t3876 VGND 0.05001f
C45993 VPWR.t3874 VGND 0.05001f
C45994 VPWR.t4020 VGND 0.05001f
C45995 VPWR.t5866 VGND 0.05001f
C45996 VPWR.t4638 VGND 0.05001f
C45997 VPWR.t4415 VGND 0.04231f
C45998 VPWR.t1723 VGND 0.0202f
C45999 VPWR.n2536 VGND 0.05372f
C46000 VPWR.t4147 VGND 0.00433f
C46001 VPWR.t4746 VGND 0.00433f
C46002 VPWR.t3494 VGND 0.00433f
C46003 VPWR.t2911 VGND 0.00433f
C46004 VPWR.t3086 VGND 0.00433f
C46005 VPWR.t3312 VGND 0.00433f
C46006 VPWR.t2195 VGND 0.00433f
C46007 VPWR.t2807 VGND 0.00433f
C46008 VPWR.t3128 VGND 0.00433f
C46009 VPWR.t5754 VGND 0.00433f
C46010 VPWR.t630 VGND 0.00433f
C46011 VPWR.t4146 VGND 0.08751f
C46012 VPWR.t2910 VGND 0.10001f
C46013 VPWR.t3085 VGND 0.10001f
C46014 VPWR.t2194 VGND 0.10001f
C46015 VPWR.t3127 VGND 0.06731f
C46016 VPWR.n2537 VGND 0.03642f
C46017 VPWR.t3243 VGND 0.00433f
C46018 VPWR.t4753 VGND 0.00433f
C46019 VPWR.t3593 VGND 0.00433f
C46020 VPWR.t2069 VGND 0.00433f
C46021 VPWR.t2717 VGND 0.00433f
C46022 VPWR.t629 VGND 0.03751f
C46023 VPWR.t3242 VGND 0.04231f
C46024 VPWR.t4752 VGND 0.03271f
C46025 VPWR.t3592 VGND 0.05001f
C46026 VPWR.t2068 VGND 0.04231f
C46027 VPWR.t2716 VGND 0.0202f
C46028 VPWR.n2538 VGND 0.05372f
C46029 VPWR.t5473 VGND 0.00433f
C46030 VPWR.t2236 VGND 0.00433f
C46031 VPWR.t5875 VGND 0.00433f
C46032 VPWR.t7072 VGND 0.00433f
C46033 VPWR.t4932 VGND 0.00433f
C46034 VPWR.t6356 VGND 0.00433f
C46035 VPWR.t3408 VGND 0.00433f
C46036 VPWR.t925 VGND 0.00433f
C46037 VPWR.t1252 VGND 0.00433f
C46038 VPWR.t5148 VGND 0.00433f
C46039 VPWR.t2410 VGND 0.00433f
C46040 VPWR.t4547 VGND 0.00433f
C46041 VPWR.t2073 VGND 0.00433f
C46042 VPWR.t5399 VGND 0.00433f
C46043 VPWR.t5309 VGND 0.00433f
C46044 VPWR.t5897 VGND 0.00433f
C46045 VPWR.t1843 VGND 0.00433f
C46046 VPWR.t2235 VGND 0.08751f
C46047 VPWR.t5874 VGND 0.10001f
C46048 VPWR.t4931 VGND 0.10001f
C46049 VPWR.t924 VGND 0.10001f
C46050 VPWR.t1251 VGND 0.10001f
C46051 VPWR.t2409 VGND 0.10001f
C46052 VPWR.t2072 VGND 0.10001f
C46053 VPWR.t5308 VGND 0.06731f
C46054 VPWR.n2539 VGND 0.03642f
C46055 VPWR.t2243 VGND 0.00433f
C46056 VPWR.t2268 VGND 0.00433f
C46057 VPWR.t4738 VGND 0.00433f
C46058 VPWR.t1018 VGND 0.00433f
C46059 VPWR.t420 VGND 0.00433f
C46060 VPWR.t1992 VGND 0.00433f
C46061 VPWR.t1634 VGND 0.00433f
C46062 VPWR.t1096 VGND 0.00433f
C46063 VPWR.t3520 VGND 0.00433f
C46064 VPWR.t3025 VGND 0.00433f
C46065 VPWR.t4899 VGND 0.00433f
C46066 VPWR.t1842 VGND 0.03751f
C46067 VPWR.t2242 VGND 0.05001f
C46068 VPWR.t2267 VGND 0.05001f
C46069 VPWR.t4737 VGND 0.05001f
C46070 VPWR.t1017 VGND 0.05001f
C46071 VPWR.t419 VGND 0.05001f
C46072 VPWR.t1991 VGND 0.05001f
C46073 VPWR.t1633 VGND 0.05001f
C46074 VPWR.t1095 VGND 0.05001f
C46075 VPWR.t3519 VGND 0.05001f
C46076 VPWR.t3024 VGND 0.04231f
C46077 VPWR.t4898 VGND 0.0202f
C46078 VPWR.n2540 VGND 0.05372f
C46079 VPWR.t2104 VGND 0.00433f
C46080 VPWR.t4534 VGND 0.00433f
C46081 VPWR.t5557 VGND 0.00433f
C46082 VPWR.t628 VGND 0.00433f
C46083 VPWR.t1984 VGND 0.00433f
C46084 VPWR.t2103 VGND 0.05481f
C46085 VPWR.t627 VGND 0.05001f
C46086 VPWR.t758 VGND 0.0202f
C46087 VPWR.t6079 VGND 0.04231f
C46088 VPWR.t5227 VGND 0.05001f
C46089 VPWR.t4781 VGND 0.05001f
C46090 VPWR.t4750 VGND 0.05001f
C46091 VPWR.t616 VGND 0.05001f
C46092 VPWR.t1811 VGND 0.05001f
C46093 VPWR.t5233 VGND 0.05001f
C46094 VPWR.t1557 VGND 0.05001f
C46095 VPWR.t852 VGND 0.05001f
C46096 VPWR.t4774 VGND 0.05001f
C46097 VPWR.t5440 VGND 0.05001f
C46098 VPWR.t395 VGND 0.05001f
C46099 VPWR.t4812 VGND 0.05001f
C46100 VPWR.t635 VGND 0.05001f
C46101 VPWR.t3329 VGND 0.05001f
C46102 VPWR.t1983 VGND 0.03751f
C46103 VPWR.n2541 VGND 0.03642f
C46104 VPWR.t3330 VGND 0.00433f
C46105 VPWR.t636 VGND 0.00433f
C46106 VPWR.t4813 VGND 0.00433f
C46107 VPWR.t396 VGND 0.00433f
C46108 VPWR.t5441 VGND 0.00433f
C46109 VPWR.t4775 VGND 0.00433f
C46110 VPWR.t853 VGND 0.00433f
C46111 VPWR.t1558 VGND 0.00433f
C46112 VPWR.t5234 VGND 0.00433f
C46113 VPWR.t1812 VGND 0.00433f
C46114 VPWR.t617 VGND 0.00433f
C46115 VPWR.t4751 VGND 0.00433f
C46116 VPWR.t4782 VGND 0.00433f
C46117 VPWR.t5228 VGND 0.00433f
C46118 VPWR.t6080 VGND 0.00433f
C46119 VPWR.n2542 VGND 0.01085f
C46120 VPWR.n2543 VGND 0.0083f
C46121 VPWR.n2544 VGND 0.00994f
C46122 VPWR.n2545 VGND 0.01085f
C46123 VPWR.n2546 VGND 0.01085f
C46124 VPWR.n2547 VGND 0.01085f
C46125 VPWR.n2548 VGND 0.00839f
C46126 VPWR.n2549 VGND 0.00985f
C46127 VPWR.n2550 VGND 0.01085f
C46128 VPWR.n2551 VGND 0.01085f
C46129 VPWR.n2552 VGND 0.01085f
C46130 VPWR.n2553 VGND 0.01085f
C46131 VPWR.n2554 VGND 0.01085f
C46132 VPWR.n2555 VGND 0.01085f
C46133 VPWR.n2556 VGND 0.01023f
C46134 VPWR.n2557 VGND 0.01189f
C46135 VPWR.n2558 VGND 0.01144f
C46136 VPWR.n2559 VGND 0.01935f
C46137 VPWR.n2560 VGND 0.01303f
C46138 VPWR.n2561 VGND 0.01189f
C46139 VPWR.n2562 VGND 0.01144f
C46140 VPWR.n2563 VGND 0.01085f
C46141 VPWR.n2564 VGND 0.00839f
C46142 VPWR.n2565 VGND 0.00985f
C46143 VPWR.n2566 VGND 0.01085f
C46144 VPWR.n2567 VGND 0.01085f
C46145 VPWR.n2568 VGND 0.01085f
C46146 VPWR.n2569 VGND 0.01085f
C46147 VPWR.n2570 VGND 0.01085f
C46148 VPWR.n2571 VGND 0.01085f
C46149 VPWR.n2572 VGND 0.01023f
C46150 VPWR.n2573 VGND 0.01189f
C46151 VPWR.n2574 VGND 0.00596f
C46152 VPWR.n2575 VGND 0.01177f
C46153 VPWR.n2576 VGND 0.02025f
C46154 VPWR.n2577 VGND 0.01568f
C46155 VPWR.n2578 VGND 0.02079f
C46156 VPWR.n2579 VGND 0.01577f
C46157 VPWR.n2580 VGND 0.0207f
C46158 VPWR.n2581 VGND 0.02171f
C46159 VPWR.n2582 VGND 0.02171f
C46160 VPWR.n2583 VGND 0.01762f
C46161 VPWR.n2584 VGND 0.01189f
C46162 VPWR.n2585 VGND 0.01144f
C46163 VPWR.n2586 VGND 0.01085f
C46164 VPWR.n2587 VGND 0.01085f
C46165 VPWR.n2588 VGND 0.0085f
C46166 VPWR.n2589 VGND 0.00912f
C46167 VPWR.n2590 VGND 0.01189f
C46168 VPWR.n2591 VGND 0.01144f
C46169 VPWR.n2592 VGND 0.01577f
C46170 VPWR.n2593 VGND 0.0207f
C46171 VPWR.n2594 VGND 0.02171f
C46172 VPWR.n2595 VGND 0.02171f
C46173 VPWR.n2596 VGND 0.01762f
C46174 VPWR.n2597 VGND 0.01189f
C46175 VPWR.n2598 VGND 0.0084f
C46176 VPWR.n2599 VGND 0.0083f
C46177 VPWR.n2600 VGND 0.10419f
C46178 VPWR.n2601 VGND 0.32859f
C46179 VPWR.n2602 VGND 0.01236f
C46180 VPWR.n2603 VGND 0.01189f
C46181 VPWR.n2604 VGND 0.01371f
C46182 VPWR.n2605 VGND 0.0178f
C46183 VPWR.n2606 VGND 0.0178f
C46184 VPWR.n2607 VGND 0.01679f
C46185 VPWR.n2608 VGND 0.01186f
C46186 VPWR.n2609 VGND 0.0178f
C46187 VPWR.n2610 VGND 0.0178f
C46188 VPWR.n2611 VGND 0.01839f
C46189 VPWR.t640 VGND 0.00433f
C46190 VPWR.t1117 VGND 0.00433f
C46191 VPWR.t1016 VGND 0.00433f
C46192 VPWR.t501 VGND 0.00433f
C46193 VPWR.t3133 VGND 0.00433f
C46194 VPWR.t826 VGND 0.00433f
C46195 VPWR.t5578 VGND 0.00433f
C46196 VPWR.n2612 VGND 0.0178f
C46197 VPWR.n2613 VGND 0.0178f
C46198 VPWR.n2614 VGND 0.01186f
C46199 VPWR.n2615 VGND 0.01679f
C46200 VPWR.n2616 VGND 0.0178f
C46201 VPWR.n2617 VGND 0.0178f
C46202 VPWR.n2618 VGND 0.01371f
C46203 VPWR.n2619 VGND 0.01189f
C46204 VPWR.n2620 VGND 0.03832f
C46205 VPWR.t639 VGND 0.05247f
C46206 VPWR.t1116 VGND 0.05996f
C46207 VPWR.t1015 VGND 0.05996f
C46208 VPWR.t500 VGND 0.05996f
C46209 VPWR.t3132 VGND 0.05996f
C46210 VPWR.t825 VGND 0.05996f
C46211 VPWR.t5577 VGND 0.05996f
C46212 VPWR.t4788 VGND 0.04035f
C46213 VPWR.n2621 VGND 0.03832f
C46214 VPWR.t319 VGND 0.00433f
C46215 VPWR.t861 VGND 0.00433f
C46216 VPWR.t3161 VGND 0.00433f
C46217 VPWR.t6353 VGND 0.00433f
C46218 VPWR.t2809 VGND 0.00433f
C46219 VPWR.t3555 VGND 0.00433f
C46220 VPWR.t1138 VGND 0.00433f
C46221 VPWR.t1776 VGND 0.00433f
C46222 VPWR.t318 VGND 0.05247f
C46223 VPWR.t860 VGND 0.05996f
C46224 VPWR.t3160 VGND 0.05996f
C46225 VPWR.t6352 VGND 0.05996f
C46226 VPWR.t2808 VGND 0.05996f
C46227 VPWR.t3554 VGND 0.05996f
C46228 VPWR.t1137 VGND 0.05996f
C46229 VPWR.t1775 VGND 0.04035f
C46230 VPWR.t4535 VGND 0.04035f
C46231 VPWR.t3486 VGND 0.05996f
C46232 VPWR.t379 VGND 0.05996f
C46233 VPWR.t2005 VGND 0.05996f
C46234 VPWR.t748 VGND 0.05996f
C46235 VPWR.t3811 VGND 0.05996f
C46236 VPWR.t2816 VGND 0.05996f
C46237 VPWR.t4810 VGND 0.05247f
C46238 VPWR.n2622 VGND 0.03832f
C46239 VPWR.t6448 VGND 0.04035f
C46240 VPWR.t2101 VGND 0.05996f
C46241 VPWR.t725 VGND 0.05996f
C46242 VPWR.t4896 VGND 0.05996f
C46243 VPWR.t4028 VGND 0.05996f
C46244 VPWR.t831 VGND 0.05996f
C46245 VPWR.t2803 VGND 0.05996f
C46246 VPWR.t2083 VGND 0.05247f
C46247 VPWR.n2623 VGND 0.03832f
C46248 VPWR.t2084 VGND 0.00433f
C46249 VPWR.t2804 VGND 0.00433f
C46250 VPWR.t832 VGND 0.00433f
C46251 VPWR.t4029 VGND 0.00433f
C46252 VPWR.t4897 VGND 0.00433f
C46253 VPWR.t726 VGND 0.00433f
C46254 VPWR.t2102 VGND 0.00433f
C46255 VPWR.t6449 VGND 0.00433f
C46256 VPWR.n2624 VGND 0.01839f
C46257 VPWR.n2625 VGND 0.0178f
C46258 VPWR.n2626 VGND 0.0178f
C46259 VPWR.n2627 VGND 0.01186f
C46260 VPWR.n2628 VGND 0.01679f
C46261 VPWR.n2629 VGND 0.0178f
C46262 VPWR.n2630 VGND 0.0178f
C46263 VPWR.n2631 VGND 0.01371f
C46264 VPWR.n2632 VGND 0.01189f
C46265 VPWR.n2633 VGND 0.01839f
C46266 VPWR.n2634 VGND 0.0178f
C46267 VPWR.n2635 VGND 0.0178f
C46268 VPWR.n2636 VGND 0.01186f
C46269 VPWR.n2637 VGND 0.01679f
C46270 VPWR.n2638 VGND 0.0178f
C46271 VPWR.n2639 VGND 0.0178f
C46272 VPWR.n2640 VGND 0.01371f
C46273 VPWR.n2641 VGND 0.01189f
C46274 VPWR.n2642 VGND 0.01236f
C46275 VPWR.n2643 VGND 0.58789f
C46276 VPWR.n2644 VGND 0.58789f
C46277 VPWR.n2645 VGND 0.01177f
C46278 VPWR.n2646 VGND 0.01678f
C46279 VPWR.n2647 VGND 0.02171f
C46280 VPWR.n2648 VGND 0.01577f
C46281 VPWR.n2649 VGND 0.0207f
C46282 VPWR.n2650 VGND 0.02171f
C46283 VPWR.n2651 VGND 0.02171f
C46284 VPWR.n2652 VGND 0.01762f
C46285 VPWR.n2653 VGND 0.01189f
C46286 VPWR.n2654 VGND 0.00912f
C46287 VPWR.n2655 VGND 0.01189f
C46288 VPWR.n2656 VGND 0.01144f
C46289 VPWR.n2657 VGND 0.02171f
C46290 VPWR.n2658 VGND 0.02171f
C46291 VPWR.n2659 VGND 0.01577f
C46292 VPWR.n2660 VGND 0.0207f
C46293 VPWR.n2661 VGND 0.02171f
C46294 VPWR.n2662 VGND 0.02171f
C46295 VPWR.n2663 VGND 0.01762f
C46296 VPWR.n2664 VGND 0.01189f
C46297 VPWR.n2665 VGND 0.00889f
C46298 VPWR.n2666 VGND 0.00994f
C46299 VPWR.n2667 VGND 0.01085f
C46300 VPWR.n2668 VGND 0.00782f
C46301 VPWR.n2669 VGND 0.0083f
C46302 VPWR.n2670 VGND 0.01042f
C46303 VPWR.n2671 VGND 0.01085f
C46304 VPWR.n2672 VGND 0.01085f
C46305 VPWR.n2673 VGND 0.00839f
C46306 VPWR.n2674 VGND 0.00985f
C46307 VPWR.n2675 VGND 0.01085f
C46308 VPWR.n2676 VGND 0.01085f
C46309 VPWR.n2677 VGND 0.01085f
C46310 VPWR.n2678 VGND 0.01085f
C46311 VPWR.n2679 VGND 0.01085f
C46312 VPWR.n2680 VGND 0.01085f
C46313 VPWR.n2681 VGND 0.01023f
C46314 VPWR.n2682 VGND 0.01189f
C46315 VPWR.n2683 VGND 0.00909f
C46316 VPWR.n2684 VGND 0.01303f
C46317 VPWR.n2685 VGND 0.01189f
C46318 VPWR.n2686 VGND 0.01144f
C46319 VPWR.n2687 VGND 0.0085f
C46320 VPWR.n2688 VGND 0.00974f
C46321 VPWR.n2689 VGND 0.01085f
C46322 VPWR.n2690 VGND 0.00839f
C46323 VPWR.n2691 VGND 0.00896f
C46324 VPWR.n2692 VGND 0.00665f
C46325 VPWR.n2693 VGND 0.00743f
C46326 VPWR.n2694 VGND 0.00685f
C46327 VPWR.n2695 VGND 0.00943f
C46328 VPWR.n2696 VGND 0.00729f
C46329 VPWR.n2697 VGND 0.00705f
C46330 VPWR.n2698 VGND 0.008f
C46331 VPWR.n2699 VGND 0.00646f
C46332 VPWR.n2700 VGND 0.01015f
C46333 VPWR.n2701 VGND 0.00643f
C46334 VPWR.n2702 VGND 0.0054f
C46335 VPWR.n2703 VGND 0.0077f
C46336 VPWR.n2704 VGND 0.00584f
C46337 VPWR.n2705 VGND 0.00698f
C46338 VPWR.n2706 VGND 0.00655f
C46339 VPWR.n2707 VGND 0.00604f
C46340 VPWR.n2708 VGND 0.13412f
C46341 VPWR.n2709 VGND 0.13412f
C46342 VPWR.n2710 VGND 0.0083f
C46343 VPWR.n2711 VGND 0.00912f
C46344 VPWR.n2712 VGND 0.01165f
C46345 VPWR.n2713 VGND 0.00588f
C46346 VPWR.n2714 VGND 0.008f
C46347 VPWR.n2715 VGND 0.00791f
C46348 VPWR.n2716 VGND 0.00829f
C46349 VPWR.n2717 VGND 0.008f
C46350 VPWR.n2718 VGND 0.00881f
C46351 VPWR.n2719 VGND 0.00872f
C46352 VPWR.n2720 VGND 0.00655f
C46353 VPWR.n2721 VGND 0.00655f
C46354 VPWR.n2722 VGND 0.00698f
C46355 VPWR.n2723 VGND 0.00584f
C46356 VPWR.n2724 VGND 0.0077f
C46357 VPWR.n2725 VGND 0.0054f
C46358 VPWR.n2726 VGND 0.0056f
C46359 VPWR.n2727 VGND 0.01184f
C46360 VPWR.n2728 VGND 0.00685f
C46361 VPWR.n2729 VGND 0.0057f
C46362 VPWR.n2730 VGND 0.0072f
C46363 VPWR.t2719 VGND 0.00433f
C46364 VPWR.t7084 VGND 0.00433f
C46365 VPWR.t2173 VGND 0.00433f
C46366 VPWR.t4664 VGND 0.00433f
C46367 VPWR.t565 VGND 0.00433f
C46368 VPWR.t3419 VGND 0.00433f
C46369 VPWR.t741 VGND 0.00433f
C46370 VPWR.t5904 VGND 0.00433f
C46371 VPWR.t6106 VGND 0.00433f
C46372 VPWR.t2701 VGND 0.00433f
C46373 VPWR.t6018 VGND 0.00433f
C46374 VPWR.t1885 VGND 0.00433f
C46375 VPWR.t1502 VGND 0.00433f
C46376 VPWR.t5504 VGND 0.00433f
C46377 VPWR.t6325 VGND 0.00433f
C46378 VPWR.n2731 VGND 0.01085f
C46379 VPWR.n2732 VGND 0.01085f
C46380 VPWR.n2733 VGND 0.01085f
C46381 VPWR.n2734 VGND 0.01085f
C46382 VPWR.n2735 VGND 0.01085f
C46383 VPWR.n2736 VGND 0.01013f
C46384 VPWR.n2737 VGND 0.00985f
C46385 VPWR.n2738 VGND 0.01085f
C46386 VPWR.n2739 VGND 0.01085f
C46387 VPWR.n2740 VGND 0.01085f
C46388 VPWR.n2741 VGND 0.01085f
C46389 VPWR.n2742 VGND 0.01085f
C46390 VPWR.n2743 VGND 0.01023f
C46391 VPWR.n2744 VGND 0.00627f
C46392 VPWR.n2745 VGND 0.0085f
C46393 VPWR.n2746 VGND 0.01189f
C46394 VPWR.t7131 VGND 0.04122f
C46395 VPWR.t2718 VGND 0.03271f
C46396 VPWR.t7083 VGND 0.0173f
C46397 VPWR.t2172 VGND 0.04521f
C46398 VPWR.t4663 VGND 0.05001f
C46399 VPWR.t564 VGND 0.05001f
C46400 VPWR.t3418 VGND 0.05001f
C46401 VPWR.t740 VGND 0.05001f
C46402 VPWR.t5903 VGND 0.05001f
C46403 VPWR.t6105 VGND 0.05001f
C46404 VPWR.t2700 VGND 0.05001f
C46405 VPWR.t6017 VGND 0.05001f
C46406 VPWR.t1884 VGND 0.05001f
C46407 VPWR.t1501 VGND 0.05001f
C46408 VPWR.t5503 VGND 0.05001f
C46409 VPWR.t6324 VGND 0.05001f
C46410 VPWR.t4573 VGND 0.0298f
C46411 VPWR.t4336 VGND 0.06143f
C46412 VPWR.t1060 VGND 0.00433f
C46413 VPWR.t5960 VGND 0.00433f
C46414 VPWR.t3761 VGND 0.00433f
C46415 VPWR.t5334 VGND 0.00433f
C46416 VPWR.t3954 VGND 0.00433f
C46417 VPWR.t771 VGND 0.00433f
C46418 VPWR.t1123 VGND 0.00433f
C46419 VPWR.t5538 VGND 0.00433f
C46420 VPWR.t1642 VGND 0.00433f
C46421 VPWR.t3063 VGND 0.00433f
C46422 VPWR.t7070 VGND 0.00433f
C46423 VPWR.t2833 VGND 0.00433f
C46424 VPWR.t4519 VGND 0.00433f
C46425 VPWR.t6104 VGND 0.00433f
C46426 VPWR.t603 VGND 0.00433f
C46427 VPWR.t5428 VGND 0.00433f
C46428 VPWR.t2313 VGND 0.00433f
C46429 VPWR.t1059 VGND 0.05001f
C46430 VPWR.t5959 VGND 0.0173f
C46431 VPWR.t3760 VGND 0.04521f
C46432 VPWR.t5333 VGND 0.05001f
C46433 VPWR.t3953 VGND 0.05001f
C46434 VPWR.t770 VGND 0.05001f
C46435 VPWR.t1122 VGND 0.05001f
C46436 VPWR.t5537 VGND 0.05001f
C46437 VPWR.t1641 VGND 0.05001f
C46438 VPWR.t3062 VGND 0.05001f
C46439 VPWR.t7069 VGND 0.05001f
C46440 VPWR.t2832 VGND 0.05001f
C46441 VPWR.t4518 VGND 0.05001f
C46442 VPWR.t6103 VGND 0.05001f
C46443 VPWR.t602 VGND 0.05001f
C46444 VPWR.t5427 VGND 0.0298f
C46445 VPWR.t2312 VGND 0.04122f
C46446 VPWR.t577 VGND 0.00433f
C46447 VPWR.t1180 VGND 0.00433f
C46448 VPWR.t5347 VGND 0.00433f
C46449 VPWR.t1979 VGND 0.00433f
C46450 VPWR.t3977 VGND 0.00433f
C46451 VPWR.t6348 VGND 0.00433f
C46452 VPWR.t327 VGND 0.00433f
C46453 VPWR.t4476 VGND 0.00433f
C46454 VPWR.t4577 VGND 0.00433f
C46455 VPWR.t2256 VGND 0.00433f
C46456 VPWR.t2765 VGND 0.00425f
C46457 VPWR.t3012 VGND 0.00433f
C46458 VPWR.t6644 VGND 0.00116f
C46459 VPWR.t164 VGND 0.00116f
C46460 VPWR.n2747 VGND 0.00236f
C46461 VPWR.t1351 VGND 0.00433f
C46462 VPWR.t5013 VGND 0.00255f
C46463 VPWR.t576 VGND 0.08271f
C46464 VPWR.t1978 VGND 0.10001f
C46465 VPWR.t3976 VGND 0.10001f
C46466 VPWR.t326 VGND 0.06731f
C46467 VPWR.t6391 VGND 0.0173f
C46468 VPWR.t4576 VGND 0.02277f
C46469 VPWR.t6828 VGND 0.04487f
C46470 VPWR.t2764 VGND 0.03282f
C46471 VPWR.t2255 VGND 0.03784f
C46472 VPWR.t6643 VGND 0.0173f
C46473 VPWR.t3011 VGND 0.02277f
C46474 VPWR.t163 VGND 0.05001f
C46475 VPWR.t1350 VGND 0.04789f
C46476 VPWR.t5012 VGND 0.0163f
C46477 VPWR.t2636 VGND 0.01775f
C46478 VPWR.n2748 VGND 0.03707f
C46479 VPWR.t1564 VGND 0.00433f
C46480 VPWR.n2749 VGND 0.00115f
C46481 VPWR.t3822 VGND 0.00433f
C46482 VPWR.t5748 VGND 0.00433f
C46483 VPWR.t2065 VGND 0.00433f
C46484 VPWR.t1456 VGND 0.00107f
C46485 VPWR.n2750 VGND 0.00292f
C46486 VPWR.t5249 VGND 0.00427f
C46487 VPWR.t1504 VGND 0.00433f
C46488 VPWR.t5253 VGND 0.00603f
C46489 VPWR.t986 VGND 0.00433f
C46490 VPWR.t4268 VGND 0.00433f
C46491 VPWR.t5958 VGND 0.00433f
C46492 VPWR.t4551 VGND 0.00431f
C46493 VPWR.t7116 VGND 0.00433f
C46494 VPWR.t872 VGND 0.00433f
C46495 VPWR.t162 VGND 0.01339f
C46496 VPWR.t1563 VGND 0.01652f
C46497 VPWR.t1597 VGND 0.0173f
C46498 VPWR.t1595 VGND 0.03271f
C46499 VPWR.t3821 VGND 0.03338f
C46500 VPWR.t161 VGND 0.05001f
C46501 VPWR.t5747 VGND 0.03181f
C46502 VPWR.t5011 VGND 0.01808f
C46503 VPWR.t5250 VGND 0.0451f
C46504 VPWR.t1455 VGND 0.03192f
C46505 VPWR.t2064 VGND 0.03885f
C46506 VPWR.t5248 VGND 0.05001f
C46507 VPWR.t1503 VGND 0.02277f
C46508 VPWR.t5252 VGND 0.05001f
C46509 VPWR.t985 VGND 0.04744f
C46510 VPWR.t4267 VGND 0.04521f
C46511 VPWR.t5957 VGND 0.0173f
C46512 VPWR.t4550 VGND 0.0298f
C46513 VPWR.t7115 VGND 0.02612f
C46514 VPWR.t215 VGND 0.05001f
C46515 VPWR.t871 VGND 0.08319f
C46516 VPWR.t1556 VGND 0.00433f
C46517 VPWR.t4275 VGND 0.00433f
C46518 VPWR.t573 VGND 0.00433f
C46519 VPWR.t5760 VGND 0.00433f
C46520 VPWR.t2442 VGND 0.00433f
C46521 VPWR.t2191 VGND 0.00433f
C46522 VPWR.t593 VGND 0.00433f
C46523 VPWR.t3715 VGND 0.00433f
C46524 VPWR.t2147 VGND 0.00433f
C46525 VPWR.t2106 VGND 0.00433f
C46526 VPWR.t1483 VGND 0.00433f
C46527 VPWR.t816 VGND 0.00433f
C46528 VPWR.t4572 VGND 0.00433f
C46529 VPWR.t4120 VGND 0.00433f
C46530 VPWR.t5302 VGND 0.00433f
C46531 VPWR.t3800 VGND 0.00433f
C46532 VPWR.t3394 VGND 0.00433f
C46533 VPWR.t1555 VGND 0.05001f
C46534 VPWR.t4274 VGND 0.0173f
C46535 VPWR.t572 VGND 0.04521f
C46536 VPWR.t5759 VGND 0.05001f
C46537 VPWR.t2441 VGND 0.05001f
C46538 VPWR.t2190 VGND 0.05001f
C46539 VPWR.t592 VGND 0.05001f
C46540 VPWR.t3714 VGND 0.05001f
C46541 VPWR.t2146 VGND 0.05001f
C46542 VPWR.t2105 VGND 0.05001f
C46543 VPWR.t1482 VGND 0.05001f
C46544 VPWR.t815 VGND 0.05001f
C46545 VPWR.t4571 VGND 0.05001f
C46546 VPWR.t4119 VGND 0.05001f
C46547 VPWR.t5301 VGND 0.05001f
C46548 VPWR.t3799 VGND 0.0298f
C46549 VPWR.t3393 VGND 0.04122f
C46550 VPWR.t5638 VGND 0.00433f
C46551 VPWR.t652 VGND 0.00433f
C46552 VPWR.t3668 VGND 0.00433f
C46553 VPWR.t418 VGND 0.00433f
C46554 VPWR.t5038 VGND 0.00433f
C46555 VPWR.t3697 VGND 0.00433f
C46556 VPWR.t4765 VGND 0.00433f
C46557 VPWR.t4854 VGND 0.00433f
C46558 VPWR.t2906 VGND 0.00433f
C46559 VPWR.t4164 VGND 0.00433f
C46560 VPWR.t3994 VGND 0.00433f
C46561 VPWR.t1935 VGND 0.00433f
C46562 VPWR.t2041 VGND 0.00433f
C46563 VPWR.t767 VGND 0.00433f
C46564 VPWR.t2305 VGND 0.00433f
C46565 VPWR.t931 VGND 0.00433f
C46566 VPWR.t651 VGND 0.08271f
C46567 VPWR.t417 VGND 0.10001f
C46568 VPWR.t3696 VGND 0.10001f
C46569 VPWR.t4764 VGND 0.10001f
C46570 VPWR.t2905 VGND 0.10001f
C46571 VPWR.t1934 VGND 0.10001f
C46572 VPWR.t766 VGND 0.10001f
C46573 VPWR.t930 VGND 0.06731f
C46574 VPWR.n2751 VGND 0.02233f
C46575 VPWR.n2752 VGND 0.02171f
C46576 VPWR.n2753 VGND 0.02171f
C46577 VPWR.n2754 VGND 0.01577f
C46578 VPWR.n2755 VGND 0.0207f
C46579 VPWR.n2756 VGND 0.02171f
C46580 VPWR.n2757 VGND 0.02171f
C46581 VPWR.n2758 VGND 0.01568f
C46582 VPWR.n2759 VGND 0.01165f
C46583 VPWR.n2760 VGND 0.01144f
C46584 VPWR.n2761 VGND 0.00986f
C46585 VPWR.n2762 VGND 0.13412f
C46586 VPWR.n2763 VGND 0.00656f
C46587 VPWR.n2764 VGND 0.01011f
C46588 VPWR.n2765 VGND 0.01085f
C46589 VPWR.n2766 VGND 0.01085f
C46590 VPWR.n2767 VGND 0.01085f
C46591 VPWR.n2768 VGND 0.01085f
C46592 VPWR.n2769 VGND 0.01085f
C46593 VPWR.n2770 VGND 0.01085f
C46594 VPWR.n2771 VGND 0.01085f
C46595 VPWR.n2772 VGND 0.01085f
C46596 VPWR.n2773 VGND 0.01085f
C46597 VPWR.n2774 VGND 0.01085f
C46598 VPWR.n2775 VGND 0.01085f
C46599 VPWR.n2776 VGND 0.01023f
C46600 VPWR.n2777 VGND 0.00544f
C46601 VPWR.n2778 VGND 0.00758f
C46602 VPWR.n2779 VGND 0.01189f
C46603 VPWR.n2780 VGND 0.01082f
C46604 VPWR.n2781 VGND 0.008f
C46605 VPWR.n2782 VGND 0.01015f
C46606 VPWR.n2783 VGND 0.00627f
C46607 VPWR.n2784 VGND 0.00834f
C46608 VPWR.n2785 VGND 0.0076f
C46609 VPWR.n2786 VGND 0.01209f
C46610 VPWR.n2787 VGND 0.01104f
C46611 VPWR.n2788 VGND 0.01038f
C46612 VPWR.n2789 VGND 0.00784f
C46613 VPWR.n2790 VGND 0.01104f
C46614 VPWR.n2791 VGND 0.0178f
C46615 VPWR.n2792 VGND 0.01209f
C46616 VPWR.n2793 VGND 0.00775f
C46617 VPWR.n2794 VGND 0.00912f
C46618 VPWR.n2795 VGND 0.03941f
C46619 VPWR.n2796 VGND 0.01044f
C46620 VPWR.n2797 VGND 0.00737f
C46621 VPWR.n2798 VGND 0.00766f
C46622 VPWR.n2799 VGND 0.00611f
C46623 VPWR.n2800 VGND 0.01085f
C46624 VPWR.n2801 VGND 0.01044f
C46625 VPWR.n2802 VGND 0.01085f
C46626 VPWR.n2803 VGND 0.01408f
C46627 VPWR.n2804 VGND 0.02171f
C46628 VPWR.n2805 VGND 0.01588f
C46629 VPWR.n2806 VGND 0.02059f
C46630 VPWR.n2807 VGND 0.01568f
C46631 VPWR.n2808 VGND 0.01165f
C46632 VPWR.n2809 VGND 0.01144f
C46633 VPWR.n2810 VGND 0.01085f
C46634 VPWR.n2811 VGND 0.01085f
C46635 VPWR.n2812 VGND 0.01085f
C46636 VPWR.n2813 VGND 0.01085f
C46637 VPWR.n2814 VGND 0.01085f
C46638 VPWR.n2815 VGND 0.01085f
C46639 VPWR.n2816 VGND 0.01085f
C46640 VPWR.n2817 VGND 0.01085f
C46641 VPWR.n2818 VGND 0.01085f
C46642 VPWR.n2819 VGND 0.01085f
C46643 VPWR.n2820 VGND 0.01085f
C46644 VPWR.n2821 VGND 0.01085f
C46645 VPWR.n2822 VGND 0.01085f
C46646 VPWR.n2823 VGND 0.01023f
C46647 VPWR.n2824 VGND 0.00544f
C46648 VPWR.n2825 VGND 0.00758f
C46649 VPWR.n2826 VGND 0.01189f
C46650 VPWR.n2827 VGND 0.01014f
C46651 VPWR.n2828 VGND 0.01004f
C46652 VPWR.n2829 VGND 0.13412f
C46653 VPWR.n2830 VGND 0.13412f
C46654 VPWR.n2831 VGND 0.01186f
C46655 VPWR.n2832 VGND 0.01165f
C46656 VPWR.n2833 VGND 0.00679f
C46657 VPWR.n2834 VGND 0.00462f
C46658 VPWR.n2835 VGND 0.00821f
C46659 VPWR.n2836 VGND 0.01104f
C46660 VPWR.n2837 VGND 0.01209f
C46661 VPWR.n2838 VGND 0.0076f
C46662 VPWR.n2839 VGND 0.00834f
C46663 VPWR.n2840 VGND 0.00974f
C46664 VPWR.n2841 VGND 0.00676f
C46665 VPWR.n2842 VGND 0.01116f
C46666 VPWR.n2843 VGND 0.00977f
C46667 VPWR.n2844 VGND 0.00901f
C46668 VPWR.n2845 VGND 0.01174f
C46669 VPWR.n2846 VGND 0.00665f
C46670 VPWR.t2516 VGND 0.00433f
C46671 VPWR.t4790 VGND 0.00433f
C46672 VPWR.t6650 VGND 0.00116f
C46673 VPWR.t6461 VGND 0.00116f
C46674 VPWR.n2847 VGND 0.00236f
C46675 VPWR.t4172 VGND 0.00427f
C46676 VPWR.t3897 VGND 0.00255f
C46677 VPWR.t3207 VGND 0.00107f
C46678 VPWR.n2848 VGND 0.00292f
C46679 VPWR.n2849 VGND 0.00115f
C46680 VPWR.n2850 VGND 0.00115f
C46681 VPWR.t333 VGND 0.00107f
C46682 VPWR.n2851 VGND 0.00292f
C46683 VPWR.n2852 VGND 0.01584f
C46684 VPWR.n2853 VGND 0.01848f
C46685 VPWR.n2854 VGND 0.01848f
C46686 VPWR.n2855 VGND 0.01584f
C46687 VPWR.n2856 VGND 0.00858f
C46688 VPWR.n2857 VGND 0.00963f
C46689 VPWR.n2858 VGND 0.0035f
C46690 VPWR.n2859 VGND 0.01303f
C46691 VPWR.n2860 VGND 0.01189f
C46692 VPWR.n2861 VGND 0.05372f
C46693 VPWR.t2515 VGND 0.05481f
C46694 VPWR.t6649 VGND 0.0202f
C46695 VPWR.t4171 VGND 0.02277f
C46696 VPWR.t6460 VGND 0.03885f
C46697 VPWR.t3206 VGND 0.04822f
C46698 VPWR.t3896 VGND 0.02768f
C46699 VPWR.t4173 VGND 0.01596f
C46700 VPWR.t325 VGND 0.02289f
C46701 VPWR.t5974 VGND 0.01529f
C46702 VPWR.n2863 VGND 0.03744f
C46703 VPWR.t7047 VGND 0.00826f
C46704 VPWR.t6462 VGND 0.01775f
C46705 VPWR.t2694 VGND 0.03215f
C46706 VPWR.t56 VGND 0.02411f
C46707 VPWR.t6015 VGND 0.02411f
C46708 VPWR.t5095 VGND 0.03215f
C46709 VPWR.t7046 VGND 0.01775f
C46710 VPWR.t6463 VGND 0.00826f
C46711 VPWR.t3898 VGND 0.01533f
C46712 VPWR.t3852 VGND 0.02286f
C46713 VPWR.n2865 VGND 0.03744f
C46714 VPWR.t586 VGND 0.01596f
C46715 VPWR.t5975 VGND 0.02768f
C46716 VPWR.t332 VGND 0.04822f
C46717 VPWR.t7044 VGND 0.03885f
C46718 VPWR.t584 VGND 0.02277f
C46719 VPWR.t6661 VGND 0.0202f
C46720 VPWR.t588 VGND 0.0202f
C46721 VPWR.n2866 VGND 0.03865f
C46722 VPWR.n2867 VGND 0.00145f
C46723 VPWR.t5044 VGND 0.00431f
C46724 VPWR.t6393 VGND 0.00196f
C46725 VPWR.t6030 VGND 0.00157f
C46726 VPWR.n2868 VGND 0.00539f
C46727 VPWR.t5564 VGND 0.00196f
C46728 VPWR.t899 VGND 0.00157f
C46729 VPWR.n2869 VGND 0.00539f
C46730 VPWR.n2870 VGND 0.00145f
C46731 VPWR.t6961 VGND 0.00425f
C46732 VPWR.t5570 VGND 0.0019f
C46733 VPWR.t6265 VGND 0.00427f
C46734 VPWR.t1797 VGND 0.00107f
C46735 VPWR.n2871 VGND 0.00292f
C46736 VPWR.t6421 VGND 0.00156f
C46737 VPWR.n2872 VGND 0.00505f
C46738 VPWR.t5566 VGND 0.00374f
C46739 VPWR.n2873 VGND 0.00115f
C46740 VPWR.t210 VGND 0.01172f
C46741 VPWR.t6826 VGND 0.02411f
C46742 VPWR.t3395 VGND 0.02366f
C46743 VPWR.t3724 VGND 0.02277f
C46744 VPWR.t6392 VGND 0.02277f
C46745 VPWR.t5043 VGND 0.01485f
C46746 VPWR.t6029 VGND 0.03516f
C46747 VPWR.t898 VGND 0.03516f
C46748 VPWR.t5571 VGND 0.01485f
C46749 VPWR.t5563 VGND 0.02277f
C46750 VPWR.t6428 VGND 0.02277f
C46751 VPWR.t6955 VGND 0.0259f
C46752 VPWR.t6426 VGND 0.02456f
C46753 VPWR.t6960 VGND 0.01172f
C46754 VPWR.t6264 VGND 0.0154f
C46755 VPWR.t5569 VGND 0.03405f
C46756 VPWR.t1796 VGND 0.02277f
C46757 VPWR.t6420 VGND 0.02768f
C46758 VPWR.t6262 VGND 0.02902f
C46759 VPWR.t2035 VGND 0.01741f
C46760 VPWR.t1846 VGND 0.02389f
C46761 VPWR.t6941 VGND 0.01839f
C46762 VPWR.t5565 VGND 0.07909f
C46763 VPWR.t4383 VGND 0.04309f
C46764 VPWR.n2874 VGND 0.02783f
C46765 VPWR.t5704 VGND 0.00427f
C46766 VPWR.t1848 VGND 0.00255f
C46767 VPWR.t1332 VGND 0.00107f
C46768 VPWR.n2875 VGND 0.00292f
C46769 VPWR.t6944 VGND 0.00116f
C46770 VPWR.t6656 VGND 0.00116f
C46771 VPWR.n2876 VGND 0.00236f
C46772 VPWR.t2343 VGND 0.00433f
C46773 VPWR.n2877 VGND 0.00115f
C46774 VPWR.t686 VGND 0.00433f
C46775 VPWR.t5277 VGND 0.00433f
C46776 VPWR.t1329 VGND 0.00255f
C46777 VPWR.t4303 VGND 0.00433f
C46778 VPWR.t92 VGND 0.00116f
C46779 VPWR.t6646 VGND 0.00116f
C46780 VPWR.n2878 VGND 0.00236f
C46781 VPWR.t563 VGND 0.00433f
C46782 VPWR.t4046 VGND 0.00433f
C46783 VPWR.t1833 VGND 0.01764f
C46784 VPWR.t6942 VGND 0.02478f
C46785 VPWR.t5703 VGND 0.02147f
C46786 VPWR.t6310 VGND 0.01772f
C46787 VPWR.n2879 VGND 0.03945f
C46788 VPWR.t1847 VGND 0.02534f
C46789 VPWR.t1331 VGND 0.03706f
C46790 VPWR.t5701 VGND 0.03885f
C46791 VPWR.t6943 VGND 0.01741f
C46792 VPWR.t1330 VGND 0.02277f
C46793 VPWR.t6655 VGND 0.03047f
C46794 VPWR.t93 VGND 0.0125f
C46795 VPWR.t1694 VGND 0.03271f
C46796 VPWR.t2342 VGND 0.02411f
C46797 VPWR.t2134 VGND 0.0173f
C46798 VPWR.t90 VGND 0.0211f
C46799 VPWR.t685 VGND 0.02143f
C46800 VPWR.t638 VGND 0.01775f
C46801 VPWR.n2880 VGND 0.03945f
C46802 VPWR.t1328 VGND 0.0336f
C46803 VPWR.t5276 VGND 0.04822f
C46804 VPWR.t91 VGND 0.05001f
C46805 VPWR.t4302 VGND 0.02277f
C46806 VPWR.t6645 VGND 0.0173f
C46807 VPWR.t562 VGND 0.025f
C46808 VPWR.t4045 VGND 0.04122f
C46809 VPWR.t2942 VGND 0.00433f
C46810 VPWR.t5778 VGND 0.00433f
C46811 VPWR.t3733 VGND 0.00433f
C46812 VPWR.t2792 VGND 0.00433f
C46813 VPWR.t4713 VGND 0.00433f
C46814 VPWR.t7088 VGND 0.00433f
C46815 VPWR.t5579 VGND 0.00433f
C46816 VPWR.t1254 VGND 0.00433f
C46817 VPWR.t5354 VGND 0.00433f
C46818 VPWR.t4444 VGND 0.00433f
C46819 VPWR.t3512 VGND 0.00433f
C46820 VPWR.t5871 VGND 0.00433f
C46821 VPWR.t5744 VGND 0.00433f
C46822 VPWR.t2964 VGND 0.00433f
C46823 VPWR.t1082 VGND 0.00433f
C46824 VPWR.t1471 VGND 0.00433f
C46825 VPWR.t2941 VGND 0.08271f
C46826 VPWR.t2791 VGND 0.10001f
C46827 VPWR.t4712 VGND 0.10001f
C46828 VPWR.t1253 VGND 0.10001f
C46829 VPWR.t4443 VGND 0.10001f
C46830 VPWR.t3511 VGND 0.10001f
C46831 VPWR.t2963 VGND 0.10001f
C46832 VPWR.t1081 VGND 0.06731f
C46833 VPWR.n2881 VGND 0.02233f
C46834 VPWR.n2882 VGND 0.02171f
C46835 VPWR.n2883 VGND 0.02171f
C46836 VPWR.n2884 VGND 0.01577f
C46837 VPWR.n2885 VGND 0.0207f
C46838 VPWR.n2886 VGND 0.02171f
C46839 VPWR.n2887 VGND 0.02171f
C46840 VPWR.n2888 VGND 0.01673f
C46841 VPWR.n2889 VGND 0.00893f
C46842 VPWR.n2890 VGND 0.00665f
C46843 VPWR.n2891 VGND 0.01005f
C46844 VPWR.n2892 VGND 0.00387f
C46845 VPWR.n2893 VGND 0.00627f
C46846 VPWR.n2894 VGND 0.00902f
C46847 VPWR.n2895 VGND 0.01302f
C46848 VPWR.n2896 VGND 0.01532f
C46849 VPWR.n2897 VGND 0.00775f
C46850 VPWR.n2898 VGND 0.00823f
C46851 VPWR.n2899 VGND 0.00803f
C46852 VPWR.n2900 VGND 0.00828f
C46853 VPWR.n2901 VGND 0.00858f
C46854 VPWR.n2902 VGND 0.01558f
C46855 VPWR.n2903 VGND 0.01623f
C46856 VPWR.n2904 VGND 0.00753f
C46857 VPWR.n2905 VGND 0.0174f
C46858 VPWR.n2906 VGND 0.01491f
C46859 VPWR.n2907 VGND 0.00902f
C46860 VPWR.n2908 VGND 0.00945f
C46861 VPWR.n2909 VGND 0.0029f
C46862 VPWR.n2910 VGND 0.01039f
C46863 VPWR.n2911 VGND 0.00811f
C46864 VPWR.n2912 VGND 0.01136f
C46865 VPWR.n2913 VGND 0.00932f
C46866 VPWR.n2914 VGND 0.00711f
C46867 VPWR.n2915 VGND 0.00723f
C46868 VPWR.n2916 VGND 0.01165f
C46869 VPWR.n2917 VGND 0.01119f
C46870 VPWR.n2918 VGND 0.0035f
C46871 VPWR.n2919 VGND 0.00458f
C46872 VPWR.n2920 VGND 0.00997f
C46873 VPWR.n2921 VGND 0.13412f
C46874 VPWR.n2922 VGND 0.13412f
C46875 VPWR.n2923 VGND 0.00794f
C46876 VPWR.n2924 VGND 0.00849f
C46877 VPWR.n2925 VGND 0.00947f
C46878 VPWR.n2926 VGND 0.00965f
C46879 VPWR.n2927 VGND 0.01131f
C46880 VPWR.n2928 VGND 0.00629f
C46881 VPWR.n2929 VGND 0.01092f
C46882 VPWR.n2930 VGND 0.01214f
C46883 VPWR.n2931 VGND 0.01824f
C46884 VPWR.n2932 VGND 0.01476f
C46885 VPWR.n2933 VGND 0.00513f
C46886 VPWR.n2934 VGND 0.00702f
C46887 VPWR.n2935 VGND 0.00752f
C46888 VPWR.n2936 VGND 0.00616f
C46889 VPWR.n2937 VGND 0.01147f
C46890 VPWR.n2938 VGND 0.00738f
C46891 VPWR.n2939 VGND 0.01015f
C46892 VPWR.n2940 VGND 0.00622f
C46893 VPWR.n2941 VGND 0.00532f
C46894 VPWR.n2942 VGND 0.00525f
C46895 VPWR.t5447 VGND 0.00431f
C46896 VPWR.t1752 VGND 0.00427f
C46897 VPWR.t4048 VGND 0.00107f
C46898 VPWR.n2943 VGND 0.00292f
C46899 VPWR.t2703 VGND 0.00431f
C46900 VPWR.n2944 VGND 0.00115f
C46901 VPWR.n2945 VGND 0.01099f
C46902 VPWR.n2946 VGND 0.01235f
C46903 VPWR.n2947 VGND 0.00912f
C46904 VPWR.n2948 VGND 0.011f
C46905 VPWR.n2949 VGND 0.00657f
C46906 VPWR.n2950 VGND 0.01165f
C46907 VPWR.n2951 VGND 0.02392f
C46908 VPWR.t5446 VGND 0.02712f
C46909 VPWR.t6395 VGND 0.03125f
C46910 VPWR.t1751 VGND 0.025f
C46911 VPWR.t216 VGND 0.03885f
C46912 VPWR.t4047 VGND 0.04789f
C46913 VPWR.t1749 VGND 0.0154f
C46914 VPWR.t2900 VGND 0.01395f
C46915 VPWR.t2702 VGND 0.03181f
C46916 VPWR.t48 VGND 0.02277f
C46917 VPWR.t1185 VGND 0.02579f
C46918 VPWR.t219 VGND 0.03259f
C46919 VPWR.t4012 VGND 0.0317f
C46920 VPWR.t4014 VGND 0.02779f
C46921 VPWR.t49 VGND 0.0211f
C46922 VPWR.n2952 VGND 0.02438f
C46923 VPWR.t2898 VGND 0.0202f
C46924 VPWR.n2953 VGND 0.02615f
C46925 VPWR.t2899 VGND 0.00255f
C46926 VPWR.t1977 VGND 0.00433f
C46927 VPWR.t51 VGND 0.00116f
C46928 VPWR.t6658 VGND 0.00116f
C46929 VPWR.n2954 VGND 0.00236f
C46930 VPWR.t6134 VGND 0.00433f
C46931 VPWR.t50 VGND 0.03271f
C46932 VPWR.t1976 VGND 0.02277f
C46933 VPWR.t6657 VGND 0.0298f
C46934 VPWR.t6133 VGND 0.06143f
C46935 VPWR.t4617 VGND 0.00433f
C46936 VPWR.t3865 VGND 0.00433f
C46937 VPWR.t3010 VGND 0.00433f
C46938 VPWR.t2721 VGND 0.00433f
C46939 VPWR.t2985 VGND 0.00433f
C46940 VPWR.t6359 VGND 0.00433f
C46941 VPWR.t5682 VGND 0.00433f
C46942 VPWR.t85 VGND 0.00433f
C46943 VPWR.t2328 VGND 0.00433f
C46944 VPWR.t4023 VGND 0.00433f
C46945 VPWR.t2296 VGND 0.00433f
C46946 VPWR.t2345 VGND 0.00433f
C46947 VPWR.t4501 VGND 0.00433f
C46948 VPWR.t4616 VGND 0.05001f
C46949 VPWR.t3864 VGND 0.05001f
C46950 VPWR.t3009 VGND 0.05001f
C46951 VPWR.t2720 VGND 0.05001f
C46952 VPWR.t2984 VGND 0.05001f
C46953 VPWR.t6358 VGND 0.05001f
C46954 VPWR.t5681 VGND 0.05001f
C46955 VPWR.t84 VGND 0.05001f
C46956 VPWR.t2327 VGND 0.05001f
C46957 VPWR.t4022 VGND 0.05001f
C46958 VPWR.t2295 VGND 0.05001f
C46959 VPWR.t2344 VGND 0.0298f
C46960 VPWR.t4500 VGND 0.02065f
C46961 VPWR.n2955 VGND 0.05167f
C46962 VPWR.t4887 VGND 0.00433f
C46963 VPWR.t4886 VGND 0.03929f
C46964 VPWR.n2956 VGND 0.03832f
C46965 VPWR.t567 VGND 0.00433f
C46966 VPWR.t6300 VGND 0.00433f
C46967 VPWR.t4517 VGND 0.00433f
C46968 VPWR.t3245 VGND 0.00433f
C46969 VPWR.t3686 VGND 0.00433f
C46970 VPWR.t6235 VGND 0.00433f
C46971 VPWR.t5948 VGND 0.00433f
C46972 VPWR.t3741 VGND 0.00433f
C46973 VPWR.t566 VGND 0.05247f
C46974 VPWR.t6299 VGND 0.05996f
C46975 VPWR.t4516 VGND 0.05996f
C46976 VPWR.t3244 VGND 0.05996f
C46977 VPWR.t3685 VGND 0.05996f
C46978 VPWR.t6234 VGND 0.05996f
C46979 VPWR.t5947 VGND 0.05996f
C46980 VPWR.t3740 VGND 0.04035f
C46981 VPWR.n2957 VGND 0.03832f
C46982 VPWR.t1500 VGND 0.00433f
C46983 VPWR.t3747 VGND 0.00433f
C46984 VPWR.t1893 VGND 0.00433f
C46985 VPWR.t3845 VGND 0.00433f
C46986 VPWR.t5373 VGND 0.00433f
C46987 VPWR.t6183 VGND 0.00433f
C46988 VPWR.t5055 VGND 0.00433f
C46989 VPWR.t1025 VGND 0.00433f
C46990 VPWR.t1499 VGND 0.05247f
C46991 VPWR.t3746 VGND 0.05996f
C46992 VPWR.t1892 VGND 0.05996f
C46993 VPWR.t3844 VGND 0.05996f
C46994 VPWR.t5372 VGND 0.05996f
C46995 VPWR.t6182 VGND 0.05996f
C46996 VPWR.t5054 VGND 0.05996f
C46997 VPWR.t1024 VGND 0.04035f
C46998 VPWR.n2958 VGND 0.03832f
C46999 VPWR.t4587 VGND 0.00433f
C47000 VPWR.t1809 VGND 0.00433f
C47001 VPWR.t2884 VGND 0.00433f
C47002 VPWR.t1074 VGND 0.00433f
C47003 VPWR.t1818 VGND 0.00433f
C47004 VPWR.t2470 VGND 0.00433f
C47005 VPWR.t1006 VGND 0.00433f
C47006 VPWR.t865 VGND 0.00433f
C47007 VPWR.t4586 VGND 0.05247f
C47008 VPWR.t1808 VGND 0.05996f
C47009 VPWR.t2883 VGND 0.05996f
C47010 VPWR.t1073 VGND 0.05996f
C47011 VPWR.t1817 VGND 0.05996f
C47012 VPWR.t2469 VGND 0.05996f
C47013 VPWR.t1005 VGND 0.05996f
C47014 VPWR.t864 VGND 0.04035f
C47015 VPWR.n2959 VGND 0.03832f
C47016 VPWR.t3528 VGND 0.00433f
C47017 VPWR.t3688 VGND 0.00433f
C47018 VPWR.t2130 VGND 0.00433f
C47019 VPWR.t4339 VGND 0.00433f
C47020 VPWR.t2309 VGND 0.00433f
C47021 VPWR.t4277 VGND 0.00433f
C47022 VPWR.t1088 VGND 0.00433f
C47023 VPWR.t3927 VGND 0.00433f
C47024 VPWR.t3527 VGND 0.05247f
C47025 VPWR.t3687 VGND 0.05996f
C47026 VPWR.t2129 VGND 0.05996f
C47027 VPWR.t4338 VGND 0.05996f
C47028 VPWR.t2308 VGND 0.05996f
C47029 VPWR.t4276 VGND 0.05996f
C47030 VPWR.t1087 VGND 0.05996f
C47031 VPWR.t3926 VGND 0.04035f
C47032 VPWR.n2960 VGND 0.01842f
C47033 VPWR.n2961 VGND 0.0178f
C47034 VPWR.n2962 VGND 0.0178f
C47035 VPWR.n2963 VGND 0.01186f
C47036 VPWR.n2964 VGND 0.01679f
C47037 VPWR.n2965 VGND 0.0178f
C47038 VPWR.n2966 VGND 0.0178f
C47039 VPWR.n2967 VGND 0.01371f
C47040 VPWR.n2968 VGND 0.01189f
C47041 VPWR.n2969 VGND 0.01839f
C47042 VPWR.n2970 VGND 0.01364f
C47043 VPWR.n2971 VGND 0.01177f
C47044 VPWR.n2972 VGND 0.01501f
C47045 VPWR.n2973 VGND 0.01186f
C47046 VPWR.n2974 VGND 0.01679f
C47047 VPWR.n2975 VGND 0.0178f
C47048 VPWR.n2976 VGND 0.0178f
C47049 VPWR.n2977 VGND 0.01371f
C47050 VPWR.n2978 VGND 0.01189f
C47051 VPWR.n2979 VGND 0.01839f
C47052 VPWR.n2980 VGND 0.0178f
C47053 VPWR.n2981 VGND 0.0178f
C47054 VPWR.n2982 VGND 0.01186f
C47055 VPWR.n2983 VGND 0.01679f
C47056 VPWR.n2984 VGND 0.0178f
C47057 VPWR.n2985 VGND 0.0178f
C47058 VPWR.n2986 VGND 0.01371f
C47059 VPWR.n2987 VGND 0.01189f
C47060 VPWR.n2988 VGND 0.01839f
C47061 VPWR.n2989 VGND 0.01609f
C47062 VPWR.n2990 VGND 0.01177f
C47063 VPWR.n2991 VGND 0.01256f
C47064 VPWR.n2992 VGND 0.01186f
C47065 VPWR.n2993 VGND 0.01679f
C47066 VPWR.n2994 VGND 0.0178f
C47067 VPWR.n2995 VGND 0.0178f
C47068 VPWR.n2996 VGND 0.01371f
C47069 VPWR.n2997 VGND 0.01189f
C47070 VPWR.n2998 VGND 0.01597f
C47071 VPWR.n2999 VGND 0.0133f
C47072 VPWR.n3000 VGND 0.01147f
C47073 VPWR.n3001 VGND 0.01085f
C47074 VPWR.n3002 VGND 0.01085f
C47075 VPWR.n3003 VGND 0.01085f
C47076 VPWR.n3004 VGND 0.00665f
C47077 VPWR.n3005 VGND 0.00985f
C47078 VPWR.n3006 VGND 0.01085f
C47079 VPWR.n3007 VGND 0.01013f
C47080 VPWR.n3008 VGND 0.00985f
C47081 VPWR.n3009 VGND 0.01085f
C47082 VPWR.n3010 VGND 0.01085f
C47083 VPWR.n3011 VGND 0.01085f
C47084 VPWR.n3012 VGND 0.0085f
C47085 VPWR.n3013 VGND 0.01189f
C47086 VPWR.n3014 VGND 0.00995f
C47087 VPWR.n3015 VGND 0.00561f
C47088 VPWR.n3016 VGND 0.00885f
C47089 VPWR.n3017 VGND 0.00581f
C47090 VPWR.n3018 VGND 0.01058f
C47091 VPWR.n3019 VGND 0.00701f
C47092 VPWR.n3020 VGND 0.00679f
C47093 VPWR.n3021 VGND 0.13412f
C47094 VPWR.n3022 VGND 0.13412f
C47095 VPWR.n3023 VGND 0.01289f
C47096 VPWR.n3024 VGND 0.01222f
C47097 VPWR.n3025 VGND 0.00834f
C47098 VPWR.n3026 VGND 0.01189f
C47099 VPWR.n3027 VGND 0.00912f
C47100 VPWR.n3028 VGND 0.01067f
C47101 VPWR.n3029 VGND 0.01013f
C47102 VPWR.n3030 VGND 0.00992f
C47103 VPWR.n3031 VGND 0.00387f
C47104 VPWR.n3032 VGND 0.00588f
C47105 VPWR.n3033 VGND 0.008f
C47106 VPWR.n3034 VGND 0.0085f
C47107 VPWR.n3035 VGND 0.01085f
C47108 VPWR.n3036 VGND 0.01085f
C47109 VPWR.n3037 VGND 0.01085f
C47110 VPWR.n3038 VGND 0.00974f
C47111 VPWR.n3039 VGND 0.01023f
C47112 VPWR.n3040 VGND 0.01085f
C47113 VPWR.n3041 VGND 0.01085f
C47114 VPWR.n3042 VGND 0.01144f
C47115 VPWR.t4648 VGND 0.00433f
C47116 VPWR.t2877 VGND 0.00433f
C47117 VPWR.t5562 VGND 0.00433f
C47118 VPWR.t1371 VGND 0.00433f
C47119 VPWR.t2939 VGND 0.00433f
C47120 VPWR.t4035 VGND 0.00433f
C47121 VPWR.t3615 VGND 0.00433f
C47122 VPWR.t6188 VGND 0.00433f
C47123 VPWR.t4711 VGND 0.00433f
C47124 VPWR.t2215 VGND 0.00433f
C47125 VPWR.t3459 VGND 0.00433f
C47126 VPWR.t3044 VGND 0.00433f
C47127 VPWR.n3043 VGND 0.01085f
C47128 VPWR.n3044 VGND 0.01085f
C47129 VPWR.n3045 VGND 0.01085f
C47130 VPWR.n3046 VGND 0.01085f
C47131 VPWR.n3047 VGND 0.01085f
C47132 VPWR.n3048 VGND 0.01085f
C47133 VPWR.n3049 VGND 0.01085f
C47134 VPWR.n3050 VGND 0.01085f
C47135 VPWR.n3051 VGND 0.01085f
C47136 VPWR.n3052 VGND 0.01023f
C47137 VPWR.n3053 VGND 0.00544f
C47138 VPWR.n3054 VGND 0.00758f
C47139 VPWR.n3055 VGND 0.01189f
C47140 VPWR.t2136 VGND 0.06143f
C47141 VPWR.t4647 VGND 0.05001f
C47142 VPWR.t2876 VGND 0.0173f
C47143 VPWR.t5561 VGND 0.04521f
C47144 VPWR.t1370 VGND 0.05001f
C47145 VPWR.t2938 VGND 0.05001f
C47146 VPWR.t4034 VGND 0.05001f
C47147 VPWR.t3614 VGND 0.05001f
C47148 VPWR.t6187 VGND 0.05001f
C47149 VPWR.t4710 VGND 0.05001f
C47150 VPWR.t2214 VGND 0.05001f
C47151 VPWR.t3458 VGND 0.05001f
C47152 VPWR.t3043 VGND 0.05001f
C47153 VPWR.t5644 VGND 0.05001f
C47154 VPWR.t4950 VGND 0.05001f
C47155 VPWR.t5953 VGND 0.05001f
C47156 VPWR.t3122 VGND 0.0298f
C47157 VPWR.t2025 VGND 0.06143f
C47158 VPWR.t2222 VGND 0.00433f
C47159 VPWR.t4826 VGND 0.00433f
C47160 VPWR.t1891 VGND 0.00433f
C47161 VPWR.t5336 VGND 0.00433f
C47162 VPWR.t4333 VGND 0.00433f
C47163 VPWR.t3510 VGND 0.00433f
C47164 VPWR.t2252 VGND 0.00433f
C47165 VPWR.t2444 VGND 0.00433f
C47166 VPWR.t4425 VGND 0.00433f
C47167 VPWR.t2724 VGND 0.00433f
C47168 VPWR.t4180 VGND 0.00433f
C47169 VPWR.t1648 VGND 0.00433f
C47170 VPWR.t4728 VGND 0.00433f
C47171 VPWR.t2820 VGND 0.00433f
C47172 VPWR.t1799 VGND 0.00433f
C47173 VPWR.t5436 VGND 0.00433f
C47174 VPWR.t3211 VGND 0.00433f
C47175 VPWR.t2221 VGND 0.05001f
C47176 VPWR.t4825 VGND 0.0173f
C47177 VPWR.t1890 VGND 0.04521f
C47178 VPWR.t5335 VGND 0.05001f
C47179 VPWR.t4332 VGND 0.05001f
C47180 VPWR.t3509 VGND 0.05001f
C47181 VPWR.t2251 VGND 0.05001f
C47182 VPWR.t2443 VGND 0.05001f
C47183 VPWR.t4424 VGND 0.05001f
C47184 VPWR.t2723 VGND 0.05001f
C47185 VPWR.t4179 VGND 0.05001f
C47186 VPWR.t1647 VGND 0.05001f
C47187 VPWR.t4727 VGND 0.05001f
C47188 VPWR.t2819 VGND 0.05001f
C47189 VPWR.t1798 VGND 0.05001f
C47190 VPWR.t5435 VGND 0.0298f
C47191 VPWR.t3210 VGND 0.06143f
C47192 VPWR.t1716 VGND 0.00433f
C47193 VPWR.t2675 VGND 0.00433f
C47194 VPWR.t5946 VGND 0.00433f
C47195 VPWR.t3557 VGND 0.00433f
C47196 VPWR.t4200 VGND 0.00433f
C47197 VPWR.t2550 VGND 0.00433f
C47198 VPWR.t4901 VGND 0.00433f
C47199 VPWR.t3918 VGND 0.00433f
C47200 VPWR.t2014 VGND 0.00433f
C47201 VPWR.t5732 VGND 0.00433f
C47202 VPWR.t5751 VGND 0.00433f
C47203 VPWR.t1004 VGND 0.00433f
C47204 VPWR.t4633 VGND 0.00433f
C47205 VPWR.t4597 VGND 0.00433f
C47206 VPWR.t599 VGND 0.00433f
C47207 VPWR.t3964 VGND 0.00433f
C47208 VPWR.t2376 VGND 0.00433f
C47209 VPWR.t1715 VGND 0.05001f
C47210 VPWR.t2674 VGND 0.0173f
C47211 VPWR.t5945 VGND 0.04521f
C47212 VPWR.t3556 VGND 0.05001f
C47213 VPWR.t4199 VGND 0.05001f
C47214 VPWR.t2549 VGND 0.05001f
C47215 VPWR.t4900 VGND 0.05001f
C47216 VPWR.t3917 VGND 0.05001f
C47217 VPWR.t2013 VGND 0.05001f
C47218 VPWR.t5731 VGND 0.05001f
C47219 VPWR.t5750 VGND 0.05001f
C47220 VPWR.t1003 VGND 0.05001f
C47221 VPWR.t4632 VGND 0.05001f
C47222 VPWR.t4596 VGND 0.05001f
C47223 VPWR.t598 VGND 0.05001f
C47224 VPWR.t3963 VGND 0.0298f
C47225 VPWR.t2375 VGND 0.04122f
C47226 VPWR.t3562 VGND 0.00433f
C47227 VPWR.t382 VGND 0.00433f
C47228 VPWR.t1697 VGND 0.00433f
C47229 VPWR.t6100 VGND 0.00433f
C47230 VPWR.t2490 VGND 0.00433f
C47231 VPWR.t3030 VGND 0.00433f
C47232 VPWR.t4749 VGND 0.00433f
C47233 VPWR.t894 VGND 0.00433f
C47234 VPWR.t3359 VGND 0.00433f
C47235 VPWR.t2983 VGND 0.00433f
C47236 VPWR.t6137 VGND 0.00433f
C47237 VPWR.t5547 VGND 0.00433f
C47238 VPWR.t2468 VGND 0.00433f
C47239 VPWR.t339 VGND 0.00433f
C47240 VPWR.t2384 VGND 0.00433f
C47241 VPWR.t1658 VGND 0.00433f
C47242 VPWR.t381 VGND 0.08271f
C47243 VPWR.t1696 VGND 0.10001f
C47244 VPWR.t2489 VGND 0.10001f
C47245 VPWR.t893 VGND 0.10001f
C47246 VPWR.t2982 VGND 0.10001f
C47247 VPWR.t5546 VGND 0.10001f
C47248 VPWR.t338 VGND 0.10001f
C47249 VPWR.t1657 VGND 0.06731f
C47250 VPWR.n3056 VGND 0.02233f
C47251 VPWR.n3057 VGND 0.02171f
C47252 VPWR.n3058 VGND 0.02171f
C47253 VPWR.n3059 VGND 0.01577f
C47254 VPWR.n3060 VGND 0.0207f
C47255 VPWR.n3061 VGND 0.02171f
C47256 VPWR.n3062 VGND 0.02171f
C47257 VPWR.n3063 VGND 0.01568f
C47258 VPWR.n3064 VGND 0.01165f
C47259 VPWR.n3065 VGND 0.01144f
C47260 VPWR.n3066 VGND 0.01085f
C47261 VPWR.n3067 VGND 0.01085f
C47262 VPWR.n3068 VGND 0.01017f
C47263 VPWR.n3069 VGND 0.00656f
C47264 VPWR.n3070 VGND 0.0098f
C47265 VPWR.n3071 VGND 0.01085f
C47266 VPWR.n3072 VGND 0.01085f
C47267 VPWR.n3073 VGND 0.01085f
C47268 VPWR.n3074 VGND 0.01085f
C47269 VPWR.n3075 VGND 0.01085f
C47270 VPWR.n3076 VGND 0.01085f
C47271 VPWR.n3077 VGND 0.01085f
C47272 VPWR.n3078 VGND 0.01085f
C47273 VPWR.n3079 VGND 0.01085f
C47274 VPWR.n3080 VGND 0.01023f
C47275 VPWR.n3081 VGND 0.00544f
C47276 VPWR.n3082 VGND 0.00758f
C47277 VPWR.n3083 VGND 0.01189f
C47278 VPWR.n3084 VGND 0.01144f
C47279 VPWR.n3085 VGND 0.01085f
C47280 VPWR.n3086 VGND 0.01085f
C47281 VPWR.n3087 VGND 0.01085f
C47282 VPWR.n3088 VGND 0.01085f
C47283 VPWR.n3089 VGND 0.01085f
C47284 VPWR.n3090 VGND 0.01085f
C47285 VPWR.n3091 VGND 0.01085f
C47286 VPWR.n3092 VGND 0.01085f
C47287 VPWR.n3093 VGND 0.01085f
C47288 VPWR.n3094 VGND 0.01085f
C47289 VPWR.n3095 VGND 0.01085f
C47290 VPWR.n3096 VGND 0.01085f
C47291 VPWR.n3097 VGND 0.01085f
C47292 VPWR.n3098 VGND 0.01023f
C47293 VPWR.n3099 VGND 0.00544f
C47294 VPWR.n3100 VGND 0.00758f
C47295 VPWR.n3101 VGND 0.01189f
C47296 VPWR.n3102 VGND 0.01144f
C47297 VPWR.n3103 VGND 0.01085f
C47298 VPWR.n3104 VGND 0.01085f
C47299 VPWR.n3105 VGND 0.00915f
C47300 VPWR.n3106 VGND 0.00656f
C47301 VPWR.n3107 VGND 0.13412f
C47302 VPWR.n3108 VGND 0.13412f
C47303 VPWR.n3109 VGND 0.00656f
C47304 VPWR.n3110 VGND 0.00803f
C47305 VPWR.n3111 VGND 0.00676f
C47306 VPWR.n3112 VGND 0.01085f
C47307 VPWR.n3113 VGND 0.01144f
C47308 VPWR.n3114 VGND 0.01189f
C47309 VPWR.n3115 VGND 0.0085f
C47310 VPWR.n3116 VGND 0.00627f
C47311 VPWR.n3117 VGND 0.01023f
C47312 VPWR.n3118 VGND 0.01085f
C47313 VPWR.n3119 VGND 0.01085f
C47314 VPWR.n3120 VGND 0.01085f
C47315 VPWR.n3121 VGND 0.01085f
C47316 VPWR.n3122 VGND 0.01085f
C47317 VPWR.n3123 VGND 0.00985f
C47318 VPWR.n3124 VGND 0.01013f
C47319 VPWR.n3125 VGND 0.01085f
C47320 VPWR.n3126 VGND 0.01085f
C47321 VPWR.n3127 VGND 0.01085f
C47322 VPWR.n3128 VGND 0.01085f
C47323 VPWR.n3129 VGND 0.01085f
C47324 VPWR.n3130 VGND 0.01085f
C47325 VPWR.n3131 VGND 0.01144f
C47326 VPWR.t2532 VGND 0.00433f
C47327 VPWR.t3997 VGND 0.00433f
C47328 VPWR.t1756 VGND 0.00433f
C47329 VPWR.t5415 VGND 0.00433f
C47330 VPWR.t722 VGND 0.00433f
C47331 VPWR.t1396 VGND 0.00433f
C47332 VPWR.t710 VGND 0.00433f
C47333 VPWR.t1961 VGND 0.00433f
C47334 VPWR.t1506 VGND 0.00433f
C47335 VPWR.t702 VGND 0.00433f
C47336 VPWR.t1828 VGND 0.00433f
C47337 VPWR.t3922 VGND 0.00433f
C47338 VPWR.n3132 VGND 0.01085f
C47339 VPWR.n3133 VGND 0.01085f
C47340 VPWR.n3134 VGND 0.01085f
C47341 VPWR.n3135 VGND 0.01085f
C47342 VPWR.n3136 VGND 0.01085f
C47343 VPWR.n3137 VGND 0.01085f
C47344 VPWR.n3138 VGND 0.01085f
C47345 VPWR.n3139 VGND 0.01085f
C47346 VPWR.n3140 VGND 0.01085f
C47347 VPWR.n3141 VGND 0.01023f
C47348 VPWR.n3142 VGND 0.00544f
C47349 VPWR.n3143 VGND 0.00758f
C47350 VPWR.n3144 VGND 0.01189f
C47351 VPWR.t5099 VGND 0.06143f
C47352 VPWR.t2531 VGND 0.05001f
C47353 VPWR.t3996 VGND 0.0173f
C47354 VPWR.t1755 VGND 0.04521f
C47355 VPWR.t5414 VGND 0.05001f
C47356 VPWR.t721 VGND 0.05001f
C47357 VPWR.t1395 VGND 0.05001f
C47358 VPWR.t709 VGND 0.05001f
C47359 VPWR.t1960 VGND 0.05001f
C47360 VPWR.t1505 VGND 0.05001f
C47361 VPWR.t701 VGND 0.05001f
C47362 VPWR.t1827 VGND 0.05001f
C47363 VPWR.t3921 VGND 0.05001f
C47364 VPWR.t4943 VGND 0.05001f
C47365 VPWR.t1605 VGND 0.05001f
C47366 VPWR.t2097 VGND 0.05001f
C47367 VPWR.t5264 VGND 0.0298f
C47368 VPWR.t5833 VGND 0.04122f
C47369 VPWR.t2492 VGND 0.00433f
C47370 VPWR.t4591 VGND 0.00433f
C47371 VPWR.t1902 VGND 0.00433f
C47372 VPWR.t2965 VGND 0.00433f
C47373 VPWR.t416 VGND 0.00433f
C47374 VPWR.t2836 VGND 0.00433f
C47375 VPWR.t4631 VGND 0.00433f
C47376 VPWR.t1644 VGND 0.00433f
C47377 VPWR.t732 VGND 0.00433f
C47378 VPWR.t2422 VGND 0.00433f
C47379 VPWR.t1736 VGND 0.00433f
C47380 VPWR.t5220 VGND 0.00433f
C47381 VPWR.t3804 VGND 0.00433f
C47382 VPWR.t3813 VGND 0.00433f
C47383 VPWR.t1973 VGND 0.00433f
C47384 VPWR.t5984 VGND 0.00433f
C47385 VPWR.t2491 VGND 0.08271f
C47386 VPWR.t1901 VGND 0.10001f
C47387 VPWR.t415 VGND 0.10001f
C47388 VPWR.t1643 VGND 0.10001f
C47389 VPWR.t731 VGND 0.10001f
C47390 VPWR.t1735 VGND 0.10001f
C47391 VPWR.t3803 VGND 0.10001f
C47392 VPWR.t1972 VGND 0.06731f
C47393 VPWR.n3145 VGND 0.02233f
C47394 VPWR.n3146 VGND 0.02171f
C47395 VPWR.n3147 VGND 0.02171f
C47396 VPWR.n3148 VGND 0.01577f
C47397 VPWR.n3149 VGND 0.0207f
C47398 VPWR.n3150 VGND 0.02171f
C47399 VPWR.n3151 VGND 0.02171f
C47400 VPWR.n3152 VGND 0.01568f
C47401 VPWR.n3153 VGND 0.01165f
C47402 VPWR.n3154 VGND 0.01144f
C47403 VPWR.n3155 VGND 0.01085f
C47404 VPWR.n3156 VGND 0.01085f
C47405 VPWR.n3157 VGND 0.01017f
C47406 VPWR.n3158 VGND 0.00656f
C47407 VPWR.n3159 VGND 0.13412f
C47408 VPWR.n3160 VGND 0.13412f
C47409 VPWR.n3161 VGND 0.00656f
C47410 VPWR.n3162 VGND 0.0098f
C47411 VPWR.n3163 VGND 0.01085f
C47412 VPWR.n3164 VGND 0.01085f
C47413 VPWR.n3165 VGND 0.01085f
C47414 VPWR.n3166 VGND 0.01085f
C47415 VPWR.n3167 VGND 0.01085f
C47416 VPWR.n3168 VGND 0.01085f
C47417 VPWR.n3169 VGND 0.01085f
C47418 VPWR.n3170 VGND 0.01085f
C47419 VPWR.n3171 VGND 0.01085f
C47420 VPWR.n3172 VGND 0.01023f
C47421 VPWR.n3173 VGND 0.00544f
C47422 VPWR.n3174 VGND 0.00758f
C47423 VPWR.n3175 VGND 0.01189f
C47424 VPWR.n3176 VGND 0.01144f
C47425 VPWR.n3177 VGND 0.01023f
C47426 VPWR.n3178 VGND 0.00974f
C47427 VPWR.n3179 VGND 0.01085f
C47428 VPWR.n3180 VGND 0.00661f
C47429 VPWR.n3181 VGND 0.01014f
C47430 VPWR.n3182 VGND 0.00865f
C47431 VPWR.n3183 VGND 0.00964f
C47432 VPWR.n3184 VGND 0.01129f
C47433 VPWR.n3185 VGND 0.01706f
C47434 VPWR.n3186 VGND 0.01011f
C47435 VPWR.n3187 VGND 0.0116f
C47436 VPWR.n3188 VGND 0.01544f
C47437 VPWR.n3189 VGND 0.00695f
C47438 VPWR.n3190 VGND 0.00512f
C47439 VPWR.n3191 VGND 0.0112f
C47440 VPWR.n3192 VGND 0.00799f
C47441 VPWR.n3193 VGND 0.01325f
C47442 VPWR.n3194 VGND 0.0039f
C47443 VPWR.n3195 VGND 0.00712f
C47444 VPWR.n3196 VGND 0.00713f
C47445 VPWR.n3197 VGND 0.01038f
C47446 VPWR.n3198 VGND 0.00856f
C47447 VPWR.n3199 VGND 0.00899f
C47448 VPWR.n3200 VGND 0.00724f
C47449 VPWR.n3201 VGND 0.01524f
C47450 VPWR.n3202 VGND 0.00819f
C47451 VPWR.n3203 VGND 0.00884f
C47452 VPWR.n3204 VGND 0.00499f
C47453 VPWR.n3205 VGND 0.01139f
C47454 VPWR.n3206 VGND 0.00837f
C47455 VPWR.n3207 VGND 0.01433f
C47456 VPWR.n3208 VGND 0.00868f
C47457 VPWR.n3209 VGND 0.01263f
C47458 VPWR.n3210 VGND 0.01042f
C47459 VPWR.n3211 VGND 0.00772f
C47460 VPWR.n3212 VGND 0.00648f
C47461 VPWR.n3213 VGND 0.00963f
C47462 VPWR.n3214 VGND 0.01447f
C47463 VPWR.n3215 VGND 0.01414f
C47464 VPWR.n3216 VGND 0.00899f
C47465 VPWR.n3217 VGND 0.00836f
C47466 VPWR.n3218 VGND 0.01165f
C47467 VPWR.n3219 VGND 0.01213f
C47468 VPWR.n3220 VGND 0.00338f
C47469 VPWR.n3221 VGND 0.00979f
C47470 VPWR.n3222 VGND 0.13412f
C47471 VPWR.n3223 VGND 0.13412f
C47472 VPWR.n3224 VGND 0.00935f
C47473 VPWR.n3225 VGND 0.00727f
C47474 VPWR.n3226 VGND 0.01045f
C47475 VPWR.n3227 VGND 0.00618f
C47476 VPWR.n3228 VGND 0.01195f
C47477 VPWR.n3229 VGND 0.00512f
C47478 VPWR.n3230 VGND 0.00823f
C47479 VPWR.n3231 VGND 0.00611f
C47480 VPWR.n3232 VGND 0.00861f
C47481 VPWR.n3233 VGND 0.00789f
C47482 VPWR.n3234 VGND 0.00765f
C47483 VPWR.n3235 VGND 0.01197f
C47484 VPWR.n3236 VGND 0.008f
C47485 VPWR.n3237 VGND 0.0088f
C47486 VPWR.n3238 VGND 0.00823f
C47487 VPWR.n3239 VGND 0.0077f
C47488 VPWR.n3240 VGND 0.00604f
C47489 VPWR.n3241 VGND 0.00571f
C47490 VPWR.n3242 VGND 0.01062f
C47491 VPWR.n3243 VGND 0.00692f
C47492 VPWR.t6407 VGND 0.00374f
C47493 VPWR.t982 VGND 0.00431f
C47494 VPWR.t4210 VGND 0.00425f
C47495 VPWR.t168 VGND 0.00132f
C47496 VPWR.t4208 VGND 0.00132f
C47497 VPWR.n3244 VGND 0.00266f
C47498 VPWR.t4212 VGND 0.00132f
C47499 VPWR.t174 VGND 0.00132f
C47500 VPWR.n3245 VGND 0.00266f
C47501 VPWR.t6401 VGND 0.0033f
C47502 VPWR.t1883 VGND 0.00433f
C47503 VPWR.t3335 VGND 0.00433f
C47504 VPWR.t362 VGND 0.00433f
C47505 VPWR.n3246 VGND 0.01634f
C47506 VPWR.n3247 VGND 0.00633f
C47507 VPWR.n3248 VGND 0.00547f
C47508 VPWR.n3249 VGND 0.00626f
C47509 VPWR.n3250 VGND 0.0063f
C47510 VPWR.n3251 VGND 0.00864f
C47511 VPWR.n3252 VGND 0.00873f
C47512 VPWR.n3253 VGND 0.00499f
C47513 VPWR.n3254 VGND 0.01164f
C47514 VPWR.n3255 VGND 0.0314f
C47515 VPWR.t4557 VGND 0.03058f
C47516 VPWR.t6985 VGND 0.03416f
C47517 VPWR.t6510 VGND 0.01172f
C47518 VPWR.t981 VGND 0.0154f
C47519 VPWR.t6406 VGND 0.02534f
C47520 VPWR.t167 VGND 0.03527f
C47521 VPWR.t4209 VGND 0.02277f
C47522 VPWR.t4207 VGND 0.02768f
C47523 VPWR.t172 VGND 0.02277f
C47524 VPWR.t4211 VGND 0.02277f
C47525 VPWR.t6984 VGND 0.02277f
C47526 VPWR.t173 VGND 0.01172f
C47527 VPWR.t6400 VGND 0.03271f
C47528 VPWR.t1882 VGND 0.0461f
C47529 VPWR.t361 VGND 0.08271f
C47530 VPWR.t4994 VGND 0.06731f
C47531 VPWR.t2954 VGND 0.0202f
C47532 VPWR.t948 VGND 0.02612f
C47533 VPWR.t6677 VGND 0.03885f
C47534 VPWR.t3658 VGND 0.04197f
C47535 VPWR.n3256 VGND 0.0314f
C47536 VPWR.t6992 VGND 0.00431f
C47537 VPWR.n3257 VGND 0.00115f
C47538 VPWR.t2420 VGND 0.00433f
C47539 VPWR.t1157 VGND 0.00255f
C47540 VPWR.t6339 VGND 0.00116f
C47541 VPWR.t6485 VGND 0.00116f
C47542 VPWR.n3258 VGND 0.00236f
C47543 VPWR.t5217 VGND 0.00433f
C47544 VPWR.t6095 VGND 0.00433f
C47545 VPWR.t3634 VGND 0.00431f
C47546 VPWR.t4007 VGND 0.00427f
C47547 VPWR.t5836 VGND 0.00107f
C47548 VPWR.n3259 VGND 0.00292f
C47549 VPWR.t2301 VGND 0.01733f
C47550 VPWR.t946 VGND 0.0173f
C47551 VPWR.t1155 VGND 0.025f
C47552 VPWR.t6340 VGND 0.0154f
C47553 VPWR.t6991 VGND 0.03181f
C47554 VPWR.t5357 VGND 0.02277f
C47555 VPWR.t3255 VGND 0.02411f
C47556 VPWR.t3045 VGND 0.025f
C47557 VPWR.t6681 VGND 0.01652f
C47558 VPWR.t6337 VGND 0.01898f
C47559 VPWR.n3261 VGND 0.05115f
C47560 VPWR.t1156 VGND 0.03271f
C47561 VPWR.t2419 VGND 0.04744f
C47562 VPWR.t6338 VGND 0.02355f
C47563 VPWR.t6484 VGND 0.03192f
C47564 VPWR.t5216 VGND 0.01395f
C47565 VPWR.t6094 VGND 0.01395f
C47566 VPWR.t3633 VGND 0.0173f
C47567 VPWR.t3228 VGND 0.03561f
C47568 VPWR.t4006 VGND 0.025f
C47569 VPWR.t6671 VGND 0.03885f
C47570 VPWR.t5835 VGND 0.04789f
C47571 VPWR.t4004 VGND 0.0202f
C47572 VPWR.n3262 VGND 0.02113f
C47573 VPWR.n3263 VGND 0.00115f
C47574 VPWR.t4522 VGND 0.00425f
C47575 VPWR.t3629 VGND 0.00433f
C47576 VPWR.t4817 VGND 0.00255f
C47577 VPWR.t2796 VGND 0.00433f
C47578 VPWR.t7007 VGND 0.00116f
C47579 VPWR.t6473 VGND 0.00116f
C47580 VPWR.n3264 VGND 0.00236f
C47581 VPWR.t343 VGND 0.00433f
C47582 VPWR.t3193 VGND 0.00433f
C47583 VPWR.t404 VGND 0.00426f
C47584 VPWR.t5238 VGND 0.00433f
C47585 VPWR.t402 VGND 0.00164f
C47586 VPWR.t406 VGND 0.00164f
C47587 VPWR.n3265 VGND 0.00329f
C47588 VPWR.t6261 VGND 0.00433f
C47589 VPWR.t400 VGND 0.00224f
C47590 VPWR.t1338 VGND 0.00156f
C47591 VPWR.n3266 VGND 0.00428f
C47592 VPWR.t866 VGND 0.01733f
C47593 VPWR.t4818 VGND 0.0173f
C47594 VPWR.t7005 VGND 0.01172f
C47595 VPWR.t3636 VGND 0.02355f
C47596 VPWR.t6856 VGND 0.03259f
C47597 VPWR.t1411 VGND 0.02768f
C47598 VPWR.t4521 VGND 0.02411f
C47599 VPWR.t5985 VGND 0.02277f
C47600 VPWR.t7004 VGND 0.02478f
C47601 VPWR.n3268 VGND 0.02491f
C47602 VPWR.t3628 VGND 0.03743f
C47603 VPWR.t4816 VGND 0.0173f
C47604 VPWR.t2795 VGND 0.03829f
C47605 VPWR.t7006 VGND 0.02835f
C47606 VPWR.t6472 VGND 0.03672f
C47607 VPWR.t342 VGND 0.0125f
C47608 VPWR.t3192 VGND 0.03516f
C47609 VPWR.t403 VGND 0.0173f
C47610 VPWR.t401 VGND 0.03271f
C47611 VPWR.t5237 VGND 0.02277f
C47612 VPWR.t405 VGND 0.04219f
C47613 VPWR.t399 VGND 0.03505f
C47614 VPWR.t6260 VGND 0.02512f
C47615 VPWR.t1337 VGND 0.0202f
C47616 VPWR.n3269 VGND 0.02649f
C47617 VPWR.t1340 VGND 0.00127f
C47618 VPWR.n3270 VGND 0.00342f
C47619 VPWR.t4903 VGND 0.00433f
C47620 VPWR.t2175 VGND 0.00433f
C47621 VPWR.n3271 VGND 0.00115f
C47622 VPWR.t2232 VGND 0.00433f
C47623 VPWR.t2623 VGND 0.00433f
C47624 VPWR.t5616 VGND 0.00255f
C47625 VPWR.t2418 VGND 0.00433f
C47626 VPWR.t6384 VGND 0.00116f
C47627 VPWR.t6467 VGND 0.00116f
C47628 VPWR.n3272 VGND 0.00236f
C47629 VPWR.t5215 VGND 0.00433f
C47630 VPWR.t2467 VGND 0.00433f
C47631 VPWR.t3514 VGND 0.00433f
C47632 VPWR.t1937 VGND 0.00433f
C47633 VPWR.t5680 VGND 0.00433f
C47634 VPWR.t1023 VGND 0.01775f
C47635 VPWR.t1339 VGND 0.0173f
C47636 VPWR.t407 VGND 0.03204f
C47637 VPWR.t5617 VGND 0.01808f
C47638 VPWR.t4902 VGND 0.03181f
C47639 VPWR.t6385 VGND 0.05001f
C47640 VPWR.t2174 VGND 0.03338f
C47641 VPWR.t950 VGND 0.03862f
C47642 VPWR.t6101 VGND 0.0355f
C47643 VPWR.t2231 VGND 0.01652f
C47644 VPWR.t6382 VGND 0.01339f
C47645 VPWR.n3273 VGND 0.03208f
C47646 VPWR.t2622 VGND 0.0374f
C47647 VPWR.t5615 VGND 0.05001f
C47648 VPWR.t2417 VGND 0.04822f
C47649 VPWR.t6383 VGND 0.02835f
C47650 VPWR.t6466 VGND 0.03672f
C47651 VPWR.t5214 VGND 0.025f
C47652 VPWR.t2466 VGND 0.08271f
C47653 VPWR.t1936 VGND 0.06731f
C47654 VPWR.n3274 VGND 0.0165f
C47655 VPWR.n3275 VGND 0.01634f
C47656 VPWR.n3276 VGND 0.01014f
C47657 VPWR.n3277 VGND 0.00735f
C47658 VPWR.n3278 VGND 0.00963f
C47659 VPWR.n3279 VGND 0.00913f
C47660 VPWR.n3280 VGND 0.0165f
C47661 VPWR.n3281 VGND 0.01185f
C47662 VPWR.n3282 VGND 0.01011f
C47663 VPWR.n3283 VGND 0.01681f
C47664 VPWR.n3284 VGND 0.01282f
C47665 VPWR.n3285 VGND 0.00465f
C47666 VPWR.n3286 VGND 0.0112f
C47667 VPWR.n3287 VGND 0.00957f
C47668 VPWR.n3288 VGND 0.00825f
C47669 VPWR.n3289 VGND 0.007f
C47670 VPWR.n3290 VGND 0.00782f
C47671 VPWR.n3291 VGND 0.00892f
C47672 VPWR.n3292 VGND 0.00697f
C47673 VPWR.n3293 VGND 0.00823f
C47674 VPWR.n3294 VGND 0.00827f
C47675 VPWR.n3295 VGND 0.00735f
C47676 VPWR.n3296 VGND 0.00992f
C47677 VPWR.n3297 VGND 0.00778f
C47678 VPWR.n3298 VGND 0.00823f
C47679 VPWR.n3299 VGND 0.00946f
C47680 VPWR.n3300 VGND 0.01011f
C47681 VPWR.n3301 VGND 0.01165f
C47682 VPWR.n3302 VGND 0.00555f
C47683 VPWR.n3303 VGND 0.01245f
C47684 VPWR.n3304 VGND 0.01139f
C47685 VPWR.n3305 VGND 0.00692f
C47686 VPWR.n3306 VGND 0.00999f
C47687 VPWR.n3307 VGND 0.00673f
C47688 VPWR.n3308 VGND 0.00554f
C47689 VPWR.n3309 VGND 0.00704f
C47690 VPWR.n3310 VGND 0.01099f
C47691 VPWR.n3311 VGND 0.01235f
C47692 VPWR.n3312 VGND 0.01165f
C47693 VPWR.n3313 VGND 0.00893f
C47694 VPWR.n3314 VGND 0.00926f
C47695 VPWR.n3315 VGND 0.01142f
C47696 VPWR.n3316 VGND 0.01177f
C47697 VPWR.n3317 VGND 0.13412f
C47698 VPWR.n3318 VGND 0.13412f
C47699 VPWR.n3319 VGND 0.00532f
C47700 VPWR.n3320 VGND 0.00977f
C47701 VPWR.n3321 VGND 0.0044f
C47702 VPWR.n3322 VGND 0.00817f
C47703 VPWR.n3323 VGND 0.00888f
C47704 VPWR.n3324 VGND 0.01189f
C47705 VPWR.n3325 VGND 0.00912f
C47706 VPWR.n3326 VGND 0.00767f
C47707 VPWR.n3327 VGND 0.00982f
C47708 VPWR.n3328 VGND 0.00829f
C47709 VPWR.n3329 VGND 0.00917f
C47710 VPWR.n3330 VGND 0.00945f
C47711 VPWR.n3331 VGND 0.00448f
C47712 VPWR.n3332 VGND 0.00951f
C47713 VPWR.n3333 VGND 0.00834f
C47714 VPWR.n3334 VGND 0.0086f
C47715 VPWR.n3335 VGND 0.00836f
C47716 VPWR.n3336 VGND 0.00899f
C47717 VPWR.n3337 VGND 0.01256f
C47718 VPWR.t3412 VGND 0.00255f
C47719 VPWR.t103 VGND 0.00116f
C47720 VPWR.t6477 VGND 0.00116f
C47721 VPWR.n3338 VGND 0.00236f
C47722 VPWR.t1699 VGND 0.00433f
C47723 VPWR.t3638 VGND 0.00516f
C47724 VPWR.t6670 VGND 0.00433f
C47725 VPWR.t6047 VGND 0.00426f
C47726 VPWR.t412 VGND 0.00434f
C47727 VPWR.t5396 VGND 0.00433f
C47728 VPWR.t6041 VGND 0.00164f
C47729 VPWR.t6049 VGND 0.00164f
C47730 VPWR.n3339 VGND 0.00329f
C47731 VPWR.t1600 VGND 0.00433f
C47732 VPWR.t6045 VGND 0.00224f
C47733 VPWR.t3672 VGND 0.00156f
C47734 VPWR.n3340 VGND 0.00428f
C47735 VPWR.t3450 VGND 0.00433f
C47736 VPWR.n3341 VGND 0.00782f
C47737 VPWR.n3342 VGND 0.00786f
C47738 VPWR.n3343 VGND 0.01123f
C47739 VPWR.n3344 VGND 0.00576f
C47740 VPWR.n3345 VGND 0.00974f
C47741 VPWR.n3346 VGND 0.00656f
C47742 VPWR.n3347 VGND 0.00802f
C47743 VPWR.n3348 VGND 0.00873f
C47744 VPWR.n3349 VGND 0.00727f
C47745 VPWR.n3350 VGND 0.00651f
C47746 VPWR.n3351 VGND 0.00483f
C47747 VPWR.n3352 VGND 0.00581f
C47748 VPWR.n3353 VGND 0.01058f
C47749 VPWR.n3354 VGND 0.02615f
C47750 VPWR.t102 VGND 0.02355f
C47751 VPWR.t6476 VGND 0.03192f
C47752 VPWR.t1698 VGND 0.01395f
C47753 VPWR.t3637 VGND 0.01172f
C47754 VPWR.t6669 VGND 0.02277f
C47755 VPWR.t6855 VGND 0.03974f
C47756 VPWR.t411 VGND 0.04554f
C47757 VPWR.t6046 VGND 0.04554f
C47758 VPWR.t6040 VGND 0.03505f
C47759 VPWR.t5395 VGND 0.02277f
C47760 VPWR.t6048 VGND 0.0173f
C47761 VPWR.t6044 VGND 0.03271f
C47762 VPWR.t1599 VGND 0.02679f
C47763 VPWR.t3671 VGND 0.04175f
C47764 VPWR.t3669 VGND 0.03103f
C47765 VPWR.t3449 VGND 0.02556f
C47766 VPWR.t6042 VGND 0.0154f
C47767 VPWR.t2637 VGND 0.01172f
C47768 VPWR.t3221 VGND 0.03181f
C47769 VPWR.t6907 VGND 0.03538f
C47770 VPWR.t2640 VGND 0.025f
C47771 VPWR.n3355 VGND 0.02504f
C47772 VPWR.t3893 VGND 0.00433f
C47773 VPWR.t5545 VGND 0.00433f
C47774 VPWR.t2639 VGND 0.00255f
C47775 VPWR.t6906 VGND 0.00116f
C47776 VPWR.t6495 VGND 0.00116f
C47777 VPWR.n3356 VGND 0.00236f
C47778 VPWR.t2326 VGND 0.00433f
C47779 VPWR.t2178 VGND 0.00433f
C47780 VPWR.t634 VGND 0.00433f
C47781 VPWR.t2873 VGND 0.00433f
C47782 VPWR.t5916 VGND 0.00433f
C47783 VPWR.t2621 VGND 0.00433f
C47784 VPWR.t4755 VGND 0.00433f
C47785 VPWR.t1166 VGND 0.00433f
C47786 VPWR.t4630 VGND 0.00433f
C47787 VPWR.t4178 VGND 0.00433f
C47788 VPWR.t5774 VGND 0.00433f
C47789 VPWR.t3448 VGND 0.02356f
C47790 VPWR.t3892 VGND 0.01563f
C47791 VPWR.t1886 VGND 0.0173f
C47792 VPWR.t6908 VGND 0.0086f
C47793 VPWR.n3358 VGND 0.03945f
C47794 VPWR.t2638 VGND 0.0461f
C47795 VPWR.t5544 VGND 0.04822f
C47796 VPWR.t6905 VGND 0.04085f
C47797 VPWR.t6494 VGND 0.03192f
C47798 VPWR.t2325 VGND 0.01395f
C47799 VPWR.t633 VGND 0.05001f
C47800 VPWR.t2872 VGND 0.08271f
C47801 VPWR.t2620 VGND 0.10001f
C47802 VPWR.t1165 VGND 0.10001f
C47803 VPWR.t4177 VGND 0.06731f
C47804 VPWR.n3359 VGND 0.02233f
C47805 VPWR.n3360 VGND 0.01588f
C47806 VPWR.n3361 VGND 0.02059f
C47807 VPWR.n3362 VGND 0.01577f
C47808 VPWR.n3363 VGND 0.01214f
C47809 VPWR.n3364 VGND 0.00913f
C47810 VPWR.n3365 VGND 0.00865f
C47811 VPWR.n3366 VGND 0.00964f
C47812 VPWR.n3367 VGND 0.01129f
C47813 VPWR.n3368 VGND 0.01282f
C47814 VPWR.n3369 VGND 0.01165f
C47815 VPWR.n3370 VGND 0.00645f
C47816 VPWR.n3371 VGND 0.00994f
C47817 VPWR.n3372 VGND 0.00898f
C47818 VPWR.n3373 VGND 0.13412f
C47819 VPWR.n3374 VGND 0.20174f
C47820 VPWR.n3375 VGND 0.01317f
C47821 VPWR.n3376 VGND 0.01206f
C47822 VPWR.n3377 VGND 0.00648f
C47823 VPWR.n3378 VGND 0.00499f
C47824 VPWR.n3379 VGND 0.01284f
C47825 VPWR.n3380 VGND 0.01077f
C47826 VPWR.n3381 VGND 0.008f
C47827 VPWR.n3382 VGND 0.01129f
C47828 VPWR.n3383 VGND 0.01824f
C47829 VPWR.n3384 VGND 0.00561f
C47830 VPWR.n3385 VGND 0.01189f
C47831 VPWR.n3386 VGND 0.00912f
C47832 VPWR.n3387 VGND 0.01189f
C47833 VPWR.n3388 VGND 0.01762f
C47834 VPWR.n3389 VGND 0.02171f
C47835 VPWR.n3390 VGND 0.02171f
C47836 VPWR.n3391 VGND 0.0207f
C47837 VPWR.n3392 VGND 0.01577f
C47838 VPWR.n3393 VGND 0.02171f
C47839 VPWR.n3394 VGND 0.02171f
C47840 VPWR.n3395 VGND 0.02079f
C47841 VPWR.n3396 VGND 0.00541f
C47842 VPWR.n3397 VGND 0.01189f
C47843 VPWR.n3398 VGND 0.01023f
C47844 VPWR.n3399 VGND 0.00878f
C47845 VPWR.n3400 VGND 0.0083f
C47846 VPWR.n3401 VGND 0.00946f
C47847 VPWR.n3402 VGND 0.01085f
C47848 VPWR.n3403 VGND 0.01085f
C47849 VPWR.n3404 VGND 0.01085f
C47850 VPWR.n3405 VGND 0.01085f
C47851 VPWR.n3406 VGND 0.00985f
C47852 VPWR.n3407 VGND 0.00839f
C47853 VPWR.n3408 VGND 0.01085f
C47854 VPWR.n3409 VGND 0.01085f
C47855 VPWR.n3410 VGND 0.01085f
C47856 VPWR.n3411 VGND 0.01085f
C47857 VPWR.n3412 VGND 0.01085f
C47858 VPWR.n3413 VGND 0.01144f
C47859 VPWR.n3414 VGND 0.01189f
C47860 VPWR.n3415 VGND 0.00735f
C47861 VPWR.n3416 VGND 0.01077f
C47862 VPWR.n3417 VGND 0.0085f
C47863 VPWR.n3418 VGND 0.01085f
C47864 VPWR.n3419 VGND 0.01085f
C47865 VPWR.n3420 VGND 0.01085f
C47866 VPWR.n3421 VGND 0.01085f
C47867 VPWR.n3422 VGND 0.01085f
C47868 VPWR.n3423 VGND 0.01085f
C47869 VPWR.n3424 VGND 0.00985f
C47870 VPWR.n3425 VGND 0.00839f
C47871 VPWR.n3426 VGND 0.01085f
C47872 VPWR.n3427 VGND 0.01085f
C47873 VPWR.n3428 VGND 0.01085f
C47874 VPWR.n3429 VGND 0.01085f
C47875 VPWR.n3430 VGND 0.01085f
C47876 VPWR.n3431 VGND 0.01085f
C47877 VPWR.n3432 VGND 0.01144f
C47878 VPWR.t5765 VGND 0.00433f
C47879 VPWR.t3431 VGND 0.00433f
C47880 VPWR.n3433 VGND 0.01568f
C47881 VPWR.n3434 VGND 0.01097f
C47882 VPWR.n3435 VGND 0.05372f
C47883 VPWR.t3430 VGND 0.08751f
C47884 VPWR.t4285 VGND 0.10001f
C47885 VPWR.t3742 VGND 0.10001f
C47886 VPWR.t1607 VGND 0.10001f
C47887 VPWR.t2663 VGND 0.10001f
C47888 VPWR.t1999 VGND 0.10001f
C47889 VPWR.t2015 VGND 0.10001f
C47890 VPWR.t86 VGND 0.06731f
C47891 VPWR.n3436 VGND 0.02233f
C47892 VPWR.n3437 VGND 0.02171f
C47893 VPWR.n3438 VGND 0.02171f
C47894 VPWR.n3439 VGND 0.01577f
C47895 VPWR.n3440 VGND 0.0207f
C47896 VPWR.n3441 VGND 0.02134f
C47897 VPWR.n3442 VGND 0.01177f
C47898 VPWR.n3443 VGND 0.20174f
C47899 VPWR.t3649 VGND 0.00433f
C47900 VPWR.t3429 VGND 0.00433f
C47901 VPWR.n3444 VGND 0.01513f
C47902 VPWR.t2903 VGND 0.00433f
C47903 VPWR.t2886 VGND 0.00433f
C47904 VPWR.t6198 VGND 0.00433f
C47905 VPWR.t2823 VGND 0.00433f
C47906 VPWR.t2643 VGND 0.00433f
C47907 VPWR.t5178 VGND 0.00433f
C47908 VPWR.t5067 VGND 0.00433f
C47909 VPWR.t3270 VGND 0.00433f
C47910 VPWR.t3824 VGND 0.00433f
C47911 VPWR.t6052 VGND 0.00433f
C47912 VPWR.t698 VGND 0.00433f
C47913 VPWR.t4858 VGND 0.00433f
C47914 VPWR.t1211 VGND 0.00433f
C47915 VPWR.t3979 VGND 0.00433f
C47916 VPWR.t1839 VGND 0.00433f
C47917 VPWR.t3806 VGND 0.00433f
C47918 VPWR.t3978 VGND 0.0298f
C47919 VPWR.t1838 VGND 0.04521f
C47920 VPWR.t3805 VGND 0.025f
C47921 VPWR.n3445 VGND 0.00665f
C47922 VPWR.n3446 VGND 0.00723f
C47923 VPWR.n3447 VGND 0.00912f
C47924 VPWR.n3448 VGND 0.00735f
C47925 VPWR.t485 VGND 0.00433f
C47926 VPWR.t1653 VGND 0.00433f
C47927 VPWR.n3449 VGND 0.01673f
C47928 VPWR.n3450 VGND 0.01165f
C47929 VPWR.t1210 VGND 0.04122f
C47930 VPWR.t484 VGND 0.08271f
C47931 VPWR.t3428 VGND 0.10001f
C47932 VPWR.t2885 VGND 0.10001f
C47933 VPWR.t2822 VGND 0.10001f
C47934 VPWR.t2642 VGND 0.10001f
C47935 VPWR.t3269 VGND 0.10001f
C47936 VPWR.t3823 VGND 0.10001f
C47937 VPWR.t697 VGND 0.06731f
C47938 VPWR.n3451 VGND 0.02233f
C47939 VPWR.n3452 VGND 0.02171f
C47940 VPWR.n3453 VGND 0.02171f
C47941 VPWR.n3454 VGND 0.01577f
C47942 VPWR.n3455 VGND 0.0207f
C47943 VPWR.n3456 VGND 0.02134f
C47944 VPWR.n3457 VGND 0.01177f
C47945 VPWR.n3458 VGND 0.13412f
C47946 VPWR.t3612 VGND 0.00433f
C47947 VPWR.t71 VGND 0.00433f
C47948 VPWR.n3459 VGND 0.01513f
C47949 VPWR.t4549 VGND 0.00433f
C47950 VPWR.t2186 VGND 0.00433f
C47951 VPWR.t3987 VGND 0.00433f
C47952 VPWR.t3029 VGND 0.00433f
C47953 VPWR.t4370 VGND 0.00433f
C47954 VPWR.t5522 VGND 0.00433f
C47955 VPWR.t963 VGND 0.00433f
C47956 VPWR.t3156 VGND 0.00433f
C47957 VPWR.t6195 VGND 0.00433f
C47958 VPWR.t658 VGND 0.00433f
C47959 VPWR.t5459 VGND 0.00433f
C47960 VPWR.t2282 VGND 0.00433f
C47961 VPWR.t5524 VGND 0.00433f
C47962 VPWR.t1998 VGND 0.00433f
C47963 VPWR.t4905 VGND 0.00433f
C47964 VPWR.t1334 VGND 0.00433f
C47965 VPWR.t1997 VGND 0.0298f
C47966 VPWR.t4904 VGND 0.04521f
C47967 VPWR.t1333 VGND 0.025f
C47968 VPWR.n3460 VGND 0.00665f
C47969 VPWR.n3461 VGND 0.00723f
C47970 VPWR.n3462 VGND 0.00912f
C47971 VPWR.n3463 VGND 0.00735f
C47972 VPWR.t3257 VGND 0.00433f
C47973 VPWR.t1444 VGND 0.00433f
C47974 VPWR.n3464 VGND 0.01673f
C47975 VPWR.n3465 VGND 0.01165f
C47976 VPWR.t5523 VGND 0.04122f
C47977 VPWR.t1443 VGND 0.08271f
C47978 VPWR.t70 VGND 0.10001f
C47979 VPWR.t2185 VGND 0.10001f
C47980 VPWR.t3028 VGND 0.10001f
C47981 VPWR.t4369 VGND 0.10001f
C47982 VPWR.t962 VGND 0.10001f
C47983 VPWR.t657 VGND 0.10001f
C47984 VPWR.t2281 VGND 0.06731f
C47985 VPWR.n3466 VGND 0.02233f
C47986 VPWR.n3467 VGND 0.02171f
C47987 VPWR.n3468 VGND 0.02171f
C47988 VPWR.n3469 VGND 0.01577f
C47989 VPWR.n3470 VGND 0.0207f
C47990 VPWR.n3471 VGND 0.02134f
C47991 VPWR.n3472 VGND 0.01177f
C47992 VPWR.n3473 VGND 0.13412f
C47993 VPWR.t1140 VGND 0.00433f
C47994 VPWR.t4554 VGND 0.00433f
C47995 VPWR.n3474 VGND 0.01513f
C47996 VPWR.t3498 VGND 0.00433f
C47997 VPWR.t6357 VGND 0.00433f
C47998 VPWR.t1359 VGND 0.00433f
C47999 VPWR.t5698 VGND 0.00433f
C48000 VPWR.t5676 VGND 0.00433f
C48001 VPWR.t621 VGND 0.00433f
C48002 VPWR.t1398 VGND 0.00433f
C48003 VPWR.t2402 VGND 0.00433f
C48004 VPWR.t4418 VGND 0.00433f
C48005 VPWR.t6229 VGND 0.00433f
C48006 VPWR.t5344 VGND 0.00433f
C48007 VPWR.t1014 VGND 0.00433f
C48008 VPWR.t2388 VGND 0.00433f
C48009 VPWR.t430 VGND 0.00433f
C48010 VPWR.t4386 VGND 0.00433f
C48011 VPWR.t7130 VGND 0.00433f
C48012 VPWR.t429 VGND 0.0298f
C48013 VPWR.t4385 VGND 0.04521f
C48014 VPWR.t7129 VGND 0.025f
C48015 VPWR.n3475 VGND 0.00665f
C48016 VPWR.n3476 VGND 0.00723f
C48017 VPWR.n3477 VGND 0.00912f
C48018 VPWR.n3478 VGND 0.00735f
C48019 VPWR.t558 VGND 0.00433f
C48020 VPWR.t4977 VGND 0.00433f
C48021 VPWR.n3479 VGND 0.01673f
C48022 VPWR.n3480 VGND 0.01165f
C48023 VPWR.t2387 VGND 0.04122f
C48024 VPWR.t557 VGND 0.08271f
C48025 VPWR.t1139 VGND 0.10001f
C48026 VPWR.t3497 VGND 0.10001f
C48027 VPWR.t1358 VGND 0.10001f
C48028 VPWR.t620 VGND 0.10001f
C48029 VPWR.t1397 VGND 0.10001f
C48030 VPWR.t4417 VGND 0.10001f
C48031 VPWR.t1013 VGND 0.06731f
C48032 VPWR.n3481 VGND 0.02233f
C48033 VPWR.n3482 VGND 0.02171f
C48034 VPWR.n3483 VGND 0.02171f
C48035 VPWR.n3484 VGND 0.01577f
C48036 VPWR.n3485 VGND 0.0207f
C48037 VPWR.n3486 VGND 0.02134f
C48038 VPWR.n3487 VGND 0.01177f
C48039 VPWR.n3488 VGND 0.13412f
C48040 VPWR.t5197 VGND 0.00433f
C48041 VPWR.t7082 VGND 0.00433f
C48042 VPWR.n3489 VGND 0.01513f
C48043 VPWR.t422 VGND 0.00433f
C48044 VPWR.t2741 VGND 0.00433f
C48045 VPWR.t3558 VGND 0.00433f
C48046 VPWR.t3100 VGND 0.00433f
C48047 VPWR.t4910 VGND 0.00433f
C48048 VPWR.t3966 VGND 0.00433f
C48049 VPWR.t2670 VGND 0.00433f
C48050 VPWR.t3861 VGND 0.00433f
C48051 VPWR.t3491 VGND 0.00433f
C48052 VPWR.t426 VGND 0.00433f
C48053 VPWR.t1900 VGND 0.00433f
C48054 VPWR.t2821 VGND 0.00433f
C48055 VPWR.t2112 VGND 0.00433f
C48056 VPWR.t3287 VGND 0.00433f
C48057 VPWR.t4628 VGND 0.00433f
C48058 VPWR.t4703 VGND 0.00433f
C48059 VPWR.t3286 VGND 0.0298f
C48060 VPWR.t4627 VGND 0.04521f
C48061 VPWR.t4702 VGND 0.025f
C48062 VPWR.n3490 VGND 0.00665f
C48063 VPWR.n3491 VGND 0.00723f
C48064 VPWR.n3492 VGND 0.00912f
C48065 VPWR.n3493 VGND 0.00735f
C48066 VPWR.t5879 VGND 0.00433f
C48067 VPWR.t1446 VGND 0.00433f
C48068 VPWR.n3494 VGND 0.01673f
C48069 VPWR.n3495 VGND 0.01165f
C48070 VPWR.t2111 VGND 0.04122f
C48071 VPWR.t1445 VGND 0.08271f
C48072 VPWR.t5196 VGND 0.10001f
C48073 VPWR.t421 VGND 0.10001f
C48074 VPWR.t3099 VGND 0.10001f
C48075 VPWR.t3965 VGND 0.10001f
C48076 VPWR.t2669 VGND 0.10001f
C48077 VPWR.t425 VGND 0.10001f
C48078 VPWR.t1899 VGND 0.06731f
C48079 VPWR.n3496 VGND 0.02233f
C48080 VPWR.n3497 VGND 0.02171f
C48081 VPWR.n3498 VGND 0.02171f
C48082 VPWR.n3499 VGND 0.01577f
C48083 VPWR.n3500 VGND 0.0207f
C48084 VPWR.n3501 VGND 0.02134f
C48085 VPWR.n3502 VGND 0.01177f
C48086 VPWR.n3503 VGND 0.13412f
C48087 VPWR.t3090 VGND 0.00433f
C48088 VPWR.t4780 VGND 0.00433f
C48089 VPWR.n3504 VGND 0.01513f
C48090 VPWR.t4030 VGND 0.00433f
C48091 VPWR.t3820 VGND 0.00433f
C48092 VPWR.t1299 VGND 0.00433f
C48093 VPWR.t2316 VGND 0.00433f
C48094 VPWR.t5109 VGND 0.00433f
C48095 VPWR.t642 VGND 0.00433f
C48096 VPWR.t4629 VGND 0.00433f
C48097 VPWR.t3289 VGND 0.00433f
C48098 VPWR.t4761 VGND 0.00433f
C48099 VPWR.t6070 VGND 0.00433f
C48100 VPWR.t3986 VGND 0.00433f
C48101 VPWR.t329 VGND 0.00433f
C48102 VPWR.t2672 VGND 0.00433f
C48103 VPWR.t1836 VGND 0.00433f
C48104 VPWR.t4493 VGND 0.00433f
C48105 VPWR.t1523 VGND 0.00433f
C48106 VPWR.t1835 VGND 0.0298f
C48107 VPWR.t4492 VGND 0.04521f
C48108 VPWR.t1522 VGND 0.025f
C48109 VPWR.n3505 VGND 0.00665f
C48110 VPWR.n3506 VGND 0.00723f
C48111 VPWR.n3507 VGND 0.00912f
C48112 VPWR.n3508 VGND 0.00735f
C48113 VPWR.t2008 VGND 0.00433f
C48114 VPWR.t6152 VGND 0.00433f
C48115 VPWR.n3509 VGND 0.01673f
C48116 VPWR.n3510 VGND 0.01165f
C48117 VPWR.t2671 VGND 0.04122f
C48118 VPWR.t2007 VGND 0.08271f
C48119 VPWR.t3089 VGND 0.10001f
C48120 VPWR.t3819 VGND 0.10001f
C48121 VPWR.t1298 VGND 0.10001f
C48122 VPWR.t641 VGND 0.10001f
C48123 VPWR.t3288 VGND 0.10001f
C48124 VPWR.t4760 VGND 0.10001f
C48125 VPWR.t328 VGND 0.06731f
C48126 VPWR.n3511 VGND 0.02233f
C48127 VPWR.n3512 VGND 0.02171f
C48128 VPWR.n3513 VGND 0.02171f
C48129 VPWR.n3514 VGND 0.01577f
C48130 VPWR.n3515 VGND 0.0207f
C48131 VPWR.n3516 VGND 0.02134f
C48132 VPWR.n3517 VGND 0.01177f
C48133 VPWR.n3518 VGND 0.13412f
C48134 VPWR.t3034 VGND 0.00433f
C48135 VPWR.t4293 VGND 0.00433f
C48136 VPWR.n3519 VGND 0.01513f
C48137 VPWR.t5640 VGND 0.00433f
C48138 VPWR.t7080 VGND 0.00433f
C48139 VPWR.t4261 VGND 0.00433f
C48140 VPWR.t6433 VGND 0.00433f
C48141 VPWR.t317 VGND 0.00433f
C48142 VPWR.t559 VGND 0.00433f
C48143 VPWR.t5560 VGND 0.00433f
C48144 VPWR.t1142 VGND 0.00433f
C48145 VPWR.t2298 VGND 0.00433f
C48146 VPWR.t5091 VGND 0.00433f
C48147 VPWR.t3995 VGND 0.00433f
C48148 VPWR.t3541 VGND 0.00433f
C48149 VPWR.t2788 VGND 0.00433f
C48150 VPWR.t1136 VGND 0.00433f
C48151 VPWR.t4114 VGND 0.00433f
C48152 VPWR.t7074 VGND 0.00433f
C48153 VPWR.t1135 VGND 0.0298f
C48154 VPWR.t4113 VGND 0.04521f
C48155 VPWR.t7073 VGND 0.025f
C48156 VPWR.n3520 VGND 0.00665f
C48157 VPWR.n3521 VGND 0.00723f
C48158 VPWR.n3522 VGND 0.00912f
C48159 VPWR.n3523 VGND 0.00735f
C48160 VPWR.t3212 VGND 0.00433f
C48161 VPWR.t2339 VGND 0.00433f
C48162 VPWR.n3524 VGND 0.01673f
C48163 VPWR.n3525 VGND 0.01165f
C48164 VPWR.t2787 VGND 0.04122f
C48165 VPWR.t2338 VGND 0.08271f
C48166 VPWR.t3033 VGND 0.10001f
C48167 VPWR.t5639 VGND 0.10001f
C48168 VPWR.t4260 VGND 0.10001f
C48169 VPWR.t316 VGND 0.10001f
C48170 VPWR.t1141 VGND 0.10001f
C48171 VPWR.t2297 VGND 0.10001f
C48172 VPWR.t3540 VGND 0.06731f
C48173 VPWR.n3526 VGND 0.02233f
C48174 VPWR.n3527 VGND 0.02171f
C48175 VPWR.n3528 VGND 0.02171f
C48176 VPWR.n3529 VGND 0.01577f
C48177 VPWR.n3530 VGND 0.0207f
C48178 VPWR.n3531 VGND 0.02134f
C48179 VPWR.n3532 VGND 0.01177f
C48180 VPWR.n3533 VGND 0.13412f
C48181 VPWR.t5799 VGND 0.00433f
C48182 VPWR.t6028 VGND 0.00433f
C48183 VPWR.n3534 VGND 0.01513f
C48184 VPWR.t5390 VGND 0.00433f
C48185 VPWR.t1814 VGND 0.00433f
C48186 VPWR.t3233 VGND 0.00433f
C48187 VPWR.t366 VGND 0.00433f
C48188 VPWR.t4003 VGND 0.00433f
C48189 VPWR.t2514 VGND 0.00433f
C48190 VPWR.t2897 VGND 0.00433f
C48191 VPWR.t2986 VGND 0.00433f
C48192 VPWR.t2848 VGND 0.00433f
C48193 VPWR.t1394 VGND 0.00433f
C48194 VPWR.t624 VGND 0.00433f
C48195 VPWR.t69 VGND 0.00433f
C48196 VPWR.t2330 VGND 0.00433f
C48197 VPWR.t3651 VGND 0.00433f
C48198 VPWR.t2666 VGND 0.00433f
C48199 VPWR.t4420 VGND 0.00433f
C48200 VPWR.t3650 VGND 0.0298f
C48201 VPWR.t2665 VGND 0.04521f
C48202 VPWR.t4419 VGND 0.025f
C48203 VPWR.n3535 VGND 0.00665f
C48204 VPWR.n3536 VGND 0.00723f
C48205 VPWR.n3537 VGND 0.00912f
C48206 VPWR.n3538 VGND 0.00735f
C48207 VPWR.t1076 VGND 0.00433f
C48208 VPWR.t3405 VGND 0.00433f
C48209 VPWR.n3539 VGND 0.01673f
C48210 VPWR.n3540 VGND 0.01165f
C48211 VPWR.t2329 VGND 0.04122f
C48212 VPWR.t1075 VGND 0.08271f
C48213 VPWR.t5798 VGND 0.10001f
C48214 VPWR.t1813 VGND 0.10001f
C48215 VPWR.t365 VGND 0.10001f
C48216 VPWR.t2513 VGND 0.10001f
C48217 VPWR.t2896 VGND 0.10001f
C48218 VPWR.t1393 VGND 0.10001f
C48219 VPWR.t68 VGND 0.06731f
C48220 VPWR.n3541 VGND 0.02233f
C48221 VPWR.n3542 VGND 0.02171f
C48222 VPWR.n3543 VGND 0.02171f
C48223 VPWR.n3544 VGND 0.01577f
C48224 VPWR.n3545 VGND 0.0207f
C48225 VPWR.n3546 VGND 0.02134f
C48226 VPWR.n3547 VGND 0.01177f
C48227 VPWR.n3548 VGND 0.13412f
C48228 VPWR.t5243 VGND 0.00433f
C48229 VPWR.t7087 VGND 0.00433f
C48230 VPWR.n3549 VGND 0.01513f
C48231 VPWR.t4348 VGND 0.00433f
C48232 VPWR.t2180 VGND 0.00433f
C48233 VPWR.t4408 VGND 0.00433f
C48234 VPWR.t3167 VGND 0.00433f
C48235 VPWR.t6309 VGND 0.00433f
C48236 VPWR.t5712 VGND 0.00433f
C48237 VPWR.t6096 VGND 0.00433f
C48238 VPWR.t2962 VGND 0.00433f
C48239 VPWR.t5743 VGND 0.00433f
C48240 VPWR.t2414 VGND 0.00433f
C48241 VPWR.t1062 VGND 0.00433f
C48242 VPWR.t4068 VGND 0.00433f
C48243 VPWR.t4973 VGND 0.00433f
C48244 VPWR.t2850 VGND 0.00433f
C48245 VPWR.t1746 VGND 0.00433f
C48246 VPWR.t2189 VGND 0.00433f
C48247 VPWR.t2849 VGND 0.0298f
C48248 VPWR.t1745 VGND 0.04521f
C48249 VPWR.t2188 VGND 0.025f
C48250 VPWR.n3550 VGND 0.00665f
C48251 VPWR.n3551 VGND 0.00723f
C48252 VPWR.n3552 VGND 0.00912f
C48253 VPWR.n3553 VGND 0.00735f
C48254 VPWR.t2303 VGND 0.00433f
C48255 VPWR.t927 VGND 0.00433f
C48256 VPWR.n3554 VGND 0.01673f
C48257 VPWR.n3555 VGND 0.01165f
C48258 VPWR.t4972 VGND 0.04122f
C48259 VPWR.t926 VGND 0.08271f
C48260 VPWR.t5242 VGND 0.10001f
C48261 VPWR.t2179 VGND 0.10001f
C48262 VPWR.t3166 VGND 0.10001f
C48263 VPWR.t5711 VGND 0.10001f
C48264 VPWR.t2961 VGND 0.10001f
C48265 VPWR.t2413 VGND 0.10001f
C48266 VPWR.t1061 VGND 0.06731f
C48267 VPWR.n3556 VGND 0.02233f
C48268 VPWR.n3557 VGND 0.02171f
C48269 VPWR.n3558 VGND 0.02171f
C48270 VPWR.n3559 VGND 0.01577f
C48271 VPWR.n3560 VGND 0.0207f
C48272 VPWR.n3561 VGND 0.02134f
C48273 VPWR.n3562 VGND 0.01177f
C48274 VPWR.n3563 VGND 0.13412f
C48275 VPWR.t1971 VGND 0.00433f
C48276 VPWR.t3693 VGND 0.00433f
C48277 VPWR.n3564 VGND 0.01513f
C48278 VPWR.t4588 VGND 0.00433f
C48279 VPWR.t874 VGND 0.00433f
C48280 VPWR.t1568 VGND 0.00433f
C48281 VPWR.t2302 VGND 0.00433f
C48282 VPWR.t4246 VGND 0.00433f
C48283 VPWR.t1086 VGND 0.00433f
C48284 VPWR.t2040 VGND 0.00433f
C48285 VPWR.t5371 VGND 0.00433f
C48286 VPWR.t1242 VGND 0.00433f
C48287 VPWR.t5733 VGND 0.00433f
C48288 VPWR.t4194 VGND 0.00433f
C48289 VPWR.t3341 VGND 0.00433f
C48290 VPWR.t1734 VGND 0.00433f
C48291 VPWR.t5370 VGND 0.00433f
C48292 VPWR.t2617 VGND 0.00433f
C48293 VPWR.t517 VGND 0.00433f
C48294 VPWR.t5369 VGND 0.0298f
C48295 VPWR.t2616 VGND 0.04521f
C48296 VPWR.t516 VGND 0.025f
C48297 VPWR.n3565 VGND 0.00665f
C48298 VPWR.n3566 VGND 0.00723f
C48299 VPWR.n3567 VGND 0.00912f
C48300 VPWR.n3568 VGND 0.00735f
C48301 VPWR.t2118 VGND 0.00433f
C48302 VPWR.t6232 VGND 0.00433f
C48303 VPWR.n3569 VGND 0.01673f
C48304 VPWR.n3570 VGND 0.01165f
C48305 VPWR.t1733 VGND 0.04122f
C48306 VPWR.t2117 VGND 0.08271f
C48307 VPWR.t1970 VGND 0.10001f
C48308 VPWR.t873 VGND 0.10001f
C48309 VPWR.t1567 VGND 0.10001f
C48310 VPWR.t1085 VGND 0.10001f
C48311 VPWR.t2039 VGND 0.10001f
C48312 VPWR.t1241 VGND 0.10001f
C48313 VPWR.t3340 VGND 0.06731f
C48314 VPWR.n3571 VGND 0.02233f
C48315 VPWR.n3572 VGND 0.02171f
C48316 VPWR.n3573 VGND 0.02171f
C48317 VPWR.n3574 VGND 0.01577f
C48318 VPWR.n3575 VGND 0.0207f
C48319 VPWR.n3576 VGND 0.02134f
C48320 VPWR.n3577 VGND 0.01177f
C48321 VPWR.n3578 VGND 0.13412f
C48322 VPWR.t3982 VGND 0.00433f
C48323 VPWR.t802 VGND 0.00433f
C48324 VPWR.n3579 VGND 0.01513f
C48325 VPWR.t3757 VGND 0.00433f
C48326 VPWR.t5789 VGND 0.00433f
C48327 VPWR.t3909 VGND 0.00433f
C48328 VPWR.t4660 VGND 0.00433f
C48329 VPWR.t694 VGND 0.00433f
C48330 VPWR.t1931 VGND 0.00433f
C48331 VPWR.t4317 VGND 0.00433f
C48332 VPWR.t1291 VGND 0.00433f
C48333 VPWR.t2217 VGND 0.00433f
C48334 VPWR.t3863 VGND 0.00433f
C48335 VPWR.t4773 VGND 0.00433f
C48336 VPWR.t2110 VGND 0.00433f
C48337 VPWR.t2743 VGND 0.00433f
C48338 VPWR.t5290 VGND 0.00433f
C48339 VPWR.t3465 VGND 0.00433f
C48340 VPWR.t5467 VGND 0.00433f
C48341 VPWR.t5289 VGND 0.0298f
C48342 VPWR.t3464 VGND 0.04521f
C48343 VPWR.t5466 VGND 0.025f
C48344 VPWR.n3580 VGND 0.00665f
C48345 VPWR.n3581 VGND 0.00723f
C48346 VPWR.n3582 VGND 0.00912f
C48347 VPWR.n3583 VGND 0.00735f
C48348 VPWR.t3053 VGND 0.00433f
C48349 VPWR.t5207 VGND 0.00433f
C48350 VPWR.n3584 VGND 0.01673f
C48351 VPWR.n3585 VGND 0.01165f
C48352 VPWR.t2742 VGND 0.04122f
C48353 VPWR.t3052 VGND 0.08271f
C48354 VPWR.t801 VGND 0.10001f
C48355 VPWR.t3756 VGND 0.10001f
C48356 VPWR.t3908 VGND 0.10001f
C48357 VPWR.t693 VGND 0.10001f
C48358 VPWR.t1290 VGND 0.10001f
C48359 VPWR.t2216 VGND 0.10001f
C48360 VPWR.t2109 VGND 0.06731f
C48361 VPWR.n3586 VGND 0.02233f
C48362 VPWR.n3587 VGND 0.02171f
C48363 VPWR.n3588 VGND 0.02171f
C48364 VPWR.n3589 VGND 0.01577f
C48365 VPWR.n3590 VGND 0.0207f
C48366 VPWR.n3591 VGND 0.02134f
C48367 VPWR.n3592 VGND 0.01177f
C48368 VPWR.n3593 VGND 0.13412f
C48369 VPWR.t3923 VGND 0.00433f
C48370 VPWR.t2866 VGND 0.00433f
C48371 VPWR.n3594 VGND 0.01513f
C48372 VPWR.t5053 VGND 0.00433f
C48373 VPWR.t2391 VGND 0.00433f
C48374 VPWR.t3078 VGND 0.00433f
C48375 VPWR.t3048 VGND 0.00433f
C48376 VPWR.t3862 VGND 0.00433f
C48377 VPWR.t55 VGND 0.00433f
C48378 VPWR.t2699 VGND 0.00433f
C48379 VPWR.t3106 VGND 0.00433f
C48380 VPWR.t1858 VGND 0.00433f
C48381 VPWR.t5278 VGND 0.00433f
C48382 VPWR.t4584 VGND 0.00433f
C48383 VPWR.t5419 VGND 0.00433f
C48384 VPWR.t7102 VGND 0.00433f
C48385 VPWR.t6068 VGND 0.00433f
C48386 VPWR.t1784 VGND 0.00433f
C48387 VPWR.t1624 VGND 0.00433f
C48388 VPWR.t6067 VGND 0.0298f
C48389 VPWR.t1783 VGND 0.04521f
C48390 VPWR.t1623 VGND 0.025f
C48391 VPWR.n3595 VGND 0.00665f
C48392 VPWR.n3596 VGND 0.00723f
C48393 VPWR.n3597 VGND 0.00912f
C48394 VPWR.n3598 VGND 0.00735f
C48395 VPWR.t2234 VGND 0.00433f
C48396 VPWR.t6212 VGND 0.00433f
C48397 VPWR.n3599 VGND 0.01673f
C48398 VPWR.n3600 VGND 0.01165f
C48399 VPWR.t7101 VGND 0.04122f
C48400 VPWR.t2233 VGND 0.08271f
C48401 VPWR.t2865 VGND 0.10001f
C48402 VPWR.t2390 VGND 0.10001f
C48403 VPWR.t3047 VGND 0.10001f
C48404 VPWR.t54 VGND 0.10001f
C48405 VPWR.t2698 VGND 0.10001f
C48406 VPWR.t1857 VGND 0.10001f
C48407 VPWR.t4583 VGND 0.06731f
C48408 VPWR.n3601 VGND 0.02233f
C48409 VPWR.n3602 VGND 0.02171f
C48410 VPWR.n3603 VGND 0.02171f
C48411 VPWR.n3604 VGND 0.01577f
C48412 VPWR.n3605 VGND 0.0207f
C48413 VPWR.n3606 VGND 0.02134f
C48414 VPWR.n3607 VGND 0.01177f
C48415 VPWR.n3608 VGND 0.13412f
C48416 VPWR.t3201 VGND 0.00433f
C48417 VPWR.t1027 VGND 0.00433f
C48418 VPWR.n3609 VGND 0.01513f
C48419 VPWR.t3368 VGND 0.00433f
C48420 VPWR.t1988 VGND 0.00433f
C48421 VPWR.t3956 VGND 0.00433f
C48422 VPWR.t6351 VGND 0.00433f
C48423 VPWR.t1353 VGND 0.00433f
C48424 VPWR.t4642 VGND 0.00433f
C48425 VPWR.t1801 VGND 0.00433f
C48426 VPWR.t4787 VGND 0.00433f
C48427 VPWR.t2003 VGND 0.00433f
C48428 VPWR.t1898 VGND 0.00433f
C48429 VPWR.t4520 VGND 0.00433f
C48430 VPWR.t3595 VGND 0.00433f
C48431 VPWR.t2786 VGND 0.00433f
C48432 VPWR.t4786 VGND 0.00433f
C48433 VPWR.t3261 VGND 0.00433f
C48434 VPWR.t1307 VGND 0.00433f
C48435 VPWR.t4785 VGND 0.0298f
C48436 VPWR.t3260 VGND 0.04521f
C48437 VPWR.t1306 VGND 0.025f
C48438 VPWR.n3610 VGND 0.00665f
C48439 VPWR.n3611 VGND 0.00723f
C48440 VPWR.n3612 VGND 0.00912f
C48441 VPWR.n3613 VGND 0.00735f
C48442 VPWR.t4161 VGND 0.00433f
C48443 VPWR.t2944 VGND 0.00433f
C48444 VPWR.n3614 VGND 0.01673f
C48445 VPWR.n3615 VGND 0.01165f
C48446 VPWR.t2785 VGND 0.04122f
C48447 VPWR.t2943 VGND 0.08271f
C48448 VPWR.t1026 VGND 0.10001f
C48449 VPWR.t1987 VGND 0.10001f
C48450 VPWR.t3955 VGND 0.10001f
C48451 VPWR.t1352 VGND 0.10001f
C48452 VPWR.t1800 VGND 0.10001f
C48453 VPWR.t1897 VGND 0.10001f
C48454 VPWR.t3594 VGND 0.06731f
C48455 VPWR.n3616 VGND 0.02233f
C48456 VPWR.n3617 VGND 0.02171f
C48457 VPWR.n3618 VGND 0.02171f
C48458 VPWR.n3619 VGND 0.01577f
C48459 VPWR.n3620 VGND 0.0207f
C48460 VPWR.n3621 VGND 0.02134f
C48461 VPWR.n3622 VGND 0.01177f
C48462 VPWR.n3623 VGND 0.13412f
C48463 VPWR.t3407 VGND 0.00433f
C48464 VPWR.t6345 VGND 0.00433f
C48465 VPWR.n3624 VGND 0.01513f
C48466 VPWR.t648 VGND 0.00433f
C48467 VPWR.t2389 VGND 0.00433f
C48468 VPWR.t2726 VGND 0.00433f
C48469 VPWR.t4233 VGND 0.00433f
C48470 VPWR.t4001 VGND 0.00433f
C48471 VPWR.t4081 VGND 0.00433f
C48472 VPWR.t3488 VGND 0.00433f
C48473 VPWR.t1982 VGND 0.00433f
C48474 VPWR.t4355 VGND 0.00433f
C48475 VPWR.t2565 VGND 0.00433f
C48476 VPWR.t5788 VGND 0.00433f
C48477 VPWR.t4884 VGND 0.00433f
C48478 VPWR.t3925 VGND 0.00433f
C48479 VPWR.t4116 VGND 0.00433f
C48480 VPWR.t2406 VGND 0.00433f
C48481 VPWR.t3216 VGND 0.00433f
C48482 VPWR.t4115 VGND 0.0298f
C48483 VPWR.t2405 VGND 0.04521f
C48484 VPWR.t3215 VGND 0.025f
C48485 VPWR.n3625 VGND 0.00665f
C48486 VPWR.n3626 VGND 0.00723f
C48487 VPWR.n3627 VGND 0.00912f
C48488 VPWR.n3628 VGND 0.00735f
C48489 VPWR.t5076 VGND 0.00433f
C48490 VPWR.t3189 VGND 0.00433f
C48491 VPWR.n3629 VGND 0.01673f
C48492 VPWR.n3630 VGND 0.01165f
C48493 VPWR.t3924 VGND 0.04122f
C48494 VPWR.t3188 VGND 0.08271f
C48495 VPWR.t3406 VGND 0.10001f
C48496 VPWR.t647 VGND 0.10001f
C48497 VPWR.t2725 VGND 0.10001f
C48498 VPWR.t4000 VGND 0.10001f
C48499 VPWR.t1981 VGND 0.10001f
C48500 VPWR.t2564 VGND 0.10001f
C48501 VPWR.t4883 VGND 0.06731f
C48502 VPWR.n3631 VGND 0.02233f
C48503 VPWR.n3632 VGND 0.02171f
C48504 VPWR.n3633 VGND 0.02171f
C48505 VPWR.n3634 VGND 0.01577f
C48506 VPWR.n3635 VGND 0.0207f
C48507 VPWR.n3636 VGND 0.02134f
C48508 VPWR.n3637 VGND 0.01177f
C48509 VPWR.n3638 VGND 0.13412f
C48510 VPWR.t5865 VGND 0.00433f
C48511 VPWR.t4245 VGND 0.00433f
C48512 VPWR.n3639 VGND 0.01513f
C48513 VPWR.t4150 VGND 0.00433f
C48514 VPWR.t374 VGND 0.00433f
C48515 VPWR.t6355 VGND 0.00433f
C48516 VPWR.t5346 VGND 0.00433f
C48517 VPWR.t792 VGND 0.00433f
C48518 VPWR.t4533 VGND 0.00433f
C48519 VPWR.t659 VGND 0.00433f
C48520 VPWR.t3 VGND 0.00433f
C48521 VPWR.t6455 VGND 0.00433f
C48522 VPWR.t6115 VGND 0.00433f
C48523 VPWR.t483 VGND 0.00433f
C48524 VPWR.t4585 VGND 0.00433f
C48525 VPWR.t81 VGND 0.00433f
C48526 VPWR.t5314 VGND 0.00433f
C48527 VPWR.t6076 VGND 0.00433f
C48528 VPWR.t3604 VGND 0.00433f
C48529 VPWR.t5313 VGND 0.0298f
C48530 VPWR.t6075 VGND 0.04521f
C48531 VPWR.t3603 VGND 0.025f
C48532 VPWR.n3640 VGND 0.00665f
C48533 VPWR.n3641 VGND 0.00723f
C48534 VPWR.n3642 VGND 0.00912f
C48535 VPWR.n3643 VGND 0.00735f
C48536 VPWR.t1920 VGND 0.00433f
C48537 VPWR.t743 VGND 0.00433f
C48538 VPWR.n3644 VGND 0.01673f
C48539 VPWR.n3645 VGND 0.01165f
C48540 VPWR.t80 VGND 0.04122f
C48541 VPWR.t742 VGND 0.08271f
C48542 VPWR.t4244 VGND 0.10001f
C48543 VPWR.t373 VGND 0.10001f
C48544 VPWR.t5345 VGND 0.10001f
C48545 VPWR.t791 VGND 0.10001f
C48546 VPWR.t2 VGND 0.10001f
C48547 VPWR.t6114 VGND 0.10001f
C48548 VPWR.t482 VGND 0.06731f
C48549 VPWR.n3646 VGND 0.02233f
C48550 VPWR.n3647 VGND 0.02171f
C48551 VPWR.n3648 VGND 0.02171f
C48552 VPWR.n3649 VGND 0.01577f
C48553 VPWR.n3650 VGND 0.0207f
C48554 VPWR.n3651 VGND 0.02134f
C48555 VPWR.n3652 VGND 0.01177f
C48556 VPWR.n3653 VGND 0.13412f
C48557 VPWR.t6019 VGND 0.00433f
C48558 VPWR.t1189 VGND 0.00433f
C48559 VPWR.n3654 VGND 0.01513f
C48560 VPWR.t2755 VGND 0.00433f
C48561 VPWR.t6816 VGND 0.00433f
C48562 VPWR.t2187 VGND 0.00433f
C48563 VPWR.t781 VGND 0.00433f
C48564 VPWR.t3901 VGND 0.00433f
C48565 VPWR.t3105 VGND 0.00433f
C48566 VPWR.t747 VGND 0.00433f
C48567 VPWR.t2244 VGND 0.00433f
C48568 VPWR.t4548 VGND 0.00433f
C48569 VPWR.t3745 VGND 0.00433f
C48570 VPWR.t3639 VGND 0.00433f
C48571 VPWR.t2611 VGND 0.00433f
C48572 VPWR.t3723 VGND 0.00433f
C48573 VPWR.t3721 VGND 0.00433f
C48574 VPWR.t5534 VGND 0.00433f
C48575 VPWR.t4218 VGND 0.00433f
C48576 VPWR.t3720 VGND 0.0298f
C48577 VPWR.t5533 VGND 0.04521f
C48578 VPWR.t4217 VGND 0.025f
C48579 VPWR.n3655 VGND 0.00665f
C48580 VPWR.n3656 VGND 0.00723f
C48581 VPWR.n3657 VGND 0.00912f
C48582 VPWR.n3658 VGND 0.00735f
C48583 VPWR.t2583 VGND 0.00433f
C48584 VPWR.t3445 VGND 0.00433f
C48585 VPWR.n3659 VGND 0.01673f
C48586 VPWR.n3660 VGND 0.01165f
C48587 VPWR.t3722 VGND 0.04122f
C48588 VPWR.t2582 VGND 0.08271f
C48589 VPWR.t1188 VGND 0.10001f
C48590 VPWR.t2754 VGND 0.10001f
C48591 VPWR.t780 VGND 0.10001f
C48592 VPWR.t3104 VGND 0.10001f
C48593 VPWR.t746 VGND 0.10001f
C48594 VPWR.t3744 VGND 0.10001f
C48595 VPWR.t2610 VGND 0.06731f
C48596 VPWR.n3661 VGND 0.02233f
C48597 VPWR.n3662 VGND 0.02171f
C48598 VPWR.n3663 VGND 0.02171f
C48599 VPWR.n3664 VGND 0.01577f
C48600 VPWR.n3665 VGND 0.0207f
C48601 VPWR.n3666 VGND 0.02134f
C48602 VPWR.n3667 VGND 0.01177f
C48603 VPWR.n3668 VGND 0.13412f
C48604 VPWR.t6207 VGND 0.00433f
C48605 VPWR.t5465 VGND 0.00433f
C48606 VPWR.n3669 VGND 0.01513f
C48607 VPWR.t5898 VGND 0.00433f
C48608 VPWR.t4168 VGND 0.00433f
C48609 VPWR.t3040 VGND 0.00433f
C48610 VPWR.t4366 VGND 0.00433f
C48611 VPWR.t1915 VGND 0.00433f
C48612 VPWR.t384 VGND 0.00433f
C48613 VPWR.t1363 VGND 0.00433f
C48614 VPWR.t3453 VGND 0.00433f
C48615 VPWR.t2907 VGND 0.00433f
C48616 VPWR.t1460 VGND 0.00433f
C48617 VPWR.t6021 VGND 0.00433f
C48618 VPWR.t1758 VGND 0.00433f
C48619 VPWR.t4347 VGND 0.00433f
C48620 VPWR.t2169 VGND 0.00433f
C48621 VPWR.t5551 VGND 0.00433f
C48622 VPWR.t3838 VGND 0.00433f
C48623 VPWR.t2168 VGND 0.0298f
C48624 VPWR.t5550 VGND 0.04521f
C48625 VPWR.t3837 VGND 0.025f
C48626 VPWR.n3670 VGND 0.00665f
C48627 VPWR.n3671 VGND 0.00723f
C48628 VPWR.n3672 VGND 0.00912f
C48629 VPWR.n3673 VGND 0.00735f
C48630 VPWR.t3442 VGND 0.00433f
C48631 VPWR.t1378 VGND 0.00433f
C48632 VPWR.n3674 VGND 0.01673f
C48633 VPWR.n3675 VGND 0.01165f
C48634 VPWR.t4346 VGND 0.04122f
C48635 VPWR.t1377 VGND 0.08271f
C48636 VPWR.t5464 VGND 0.10001f
C48637 VPWR.t4167 VGND 0.10001f
C48638 VPWR.t3039 VGND 0.10001f
C48639 VPWR.t383 VGND 0.10001f
C48640 VPWR.t1362 VGND 0.10001f
C48641 VPWR.t1459 VGND 0.10001f
C48642 VPWR.t1757 VGND 0.06731f
C48643 VPWR.n3676 VGND 0.02233f
C48644 VPWR.n3677 VGND 0.02171f
C48645 VPWR.n3678 VGND 0.02171f
C48646 VPWR.n3679 VGND 0.01577f
C48647 VPWR.n3680 VGND 0.0207f
C48648 VPWR.n3681 VGND 0.02134f
C48649 VPWR.n3682 VGND 0.01177f
C48650 VPWR.n3683 VGND 0.13412f
C48651 VPWR.t5094 VGND 0.00433f
C48652 VPWR.t3111 VGND 0.00433f
C48653 VPWR.n3684 VGND 0.01513f
C48654 VPWR.t3440 VGND 0.00433f
C48655 VPWR.t1244 VGND 0.00433f
C48656 VPWR.t4659 VGND 0.00433f
C48657 VPWR.t1297 VGND 0.00433f
C48658 VPWR.t1540 VGND 0.00433f
C48659 VPWR.t2904 VGND 0.00433f
C48660 VPWR.t1656 VGND 0.00433f
C48661 VPWR.t965 VGND 0.00433f
C48662 VPWR.t3178 VGND 0.00433f
C48663 VPWR.t530 VGND 0.00433f
C48664 VPWR.t4287 VGND 0.00433f
C48665 VPWR.t3077 VGND 0.00433f
C48666 VPWR.t4374 VGND 0.0202f
C48667 VPWR.t4375 VGND 0.00433f
C48668 VPWR.t3343 VGND 0.00433f
C48669 VPWR.t5288 VGND 0.00433f
C48670 VPWR.t5296 VGND 0.00433f
C48671 VPWR.t3342 VGND 0.04231f
C48672 VPWR.t5287 VGND 0.05001f
C48673 VPWR.t5295 VGND 0.03271f
C48674 VPWR.t6111 VGND 0.01775f
C48675 VPWR.n3685 VGND 0.05167f
C48676 VPWR.t6112 VGND 0.00433f
C48677 VPWR.t5864 VGND 0.00433f
C48678 VPWR.t4733 VGND 0.00433f
C48679 VPWR.t2631 VGND 0.00433f
C48680 VPWR.t6185 VGND 0.00433f
C48681 VPWR.t5502 VGND 0.00433f
C48682 VPWR.t954 VGND 0.05247f
C48683 VPWR.t1821 VGND 0.05996f
C48684 VPWR.t5378 VGND 0.05996f
C48685 VPWR.t2987 VGND 0.05996f
C48686 VPWR.t856 VGND 0.05996f
C48687 VPWR.t1434 VGND 0.05996f
C48688 VPWR.t4776 VGND 0.05996f
C48689 VPWR.t1091 VGND 0.04035f
C48690 VPWR.t5863 VGND 0.0589f
C48691 VPWR.t4732 VGND 0.05996f
C48692 VPWR.t2630 VGND 0.05996f
C48693 VPWR.t6184 VGND 0.05996f
C48694 VPWR.t5501 VGND 0.05247f
C48695 VPWR.n3686 VGND 0.03832f
C48696 VPWR.t1092 VGND 0.00433f
C48697 VPWR.t4777 VGND 0.00433f
C48698 VPWR.t1435 VGND 0.00433f
C48699 VPWR.t857 VGND 0.00433f
C48700 VPWR.t2988 VGND 0.00433f
C48701 VPWR.t5379 VGND 0.00433f
C48702 VPWR.n3687 VGND 0.0178f
C48703 VPWR.n3688 VGND 0.01679f
C48704 VPWR.n3689 VGND 0.01186f
C48705 VPWR.n3690 VGND 0.0178f
C48706 VPWR.n3691 VGND 0.0178f
C48707 VPWR.n3692 VGND 0.01839f
C48708 VPWR.n3693 VGND 0.01189f
C48709 VPWR.n3694 VGND 0.01371f
C48710 VPWR.n3695 VGND 0.0178f
C48711 VPWR.n3696 VGND 0.0178f
C48712 VPWR.n3697 VGND 0.01679f
C48713 VPWR.n3698 VGND 0.01186f
C48714 VPWR.n3699 VGND 0.01315f
C48715 VPWR.n3700 VGND 0.01107f
C48716 VPWR.n3701 VGND 0.00665f
C48717 VPWR.n3702 VGND 0.01008f
C48718 VPWR.n3703 VGND 0.00974f
C48719 VPWR.n3704 VGND 0.00909f
C48720 VPWR.t4131 VGND 0.00433f
C48721 VPWR.t4294 VGND 0.00433f
C48722 VPWR.n3705 VGND 0.01762f
C48723 VPWR.n3706 VGND 0.01189f
C48724 VPWR.n3707 VGND 0.02102f
C48725 VPWR.t4130 VGND 0.08271f
C48726 VPWR.t3110 VGND 0.10001f
C48727 VPWR.t1243 VGND 0.10001f
C48728 VPWR.t1296 VGND 0.10001f
C48729 VPWR.t1539 VGND 0.10001f
C48730 VPWR.t964 VGND 0.10001f
C48731 VPWR.t529 VGND 0.10001f
C48732 VPWR.t3076 VGND 0.06731f
C48733 VPWR.n3708 VGND 0.02233f
C48734 VPWR.n3709 VGND 0.02171f
C48735 VPWR.n3710 VGND 0.02171f
C48736 VPWR.n3711 VGND 0.01577f
C48737 VPWR.n3712 VGND 0.0207f
C48738 VPWR.n3713 VGND 0.02134f
C48739 VPWR.n3714 VGND 0.01177f
C48740 VPWR.n3715 VGND 0.13412f
C48741 VPWR.n3716 VGND 0.10419f
C48742 VPWR.n3717 VGND 0.01177f
C48743 VPWR.n3718 VGND 0.01513f
C48744 VPWR.n3719 VGND 0.01568f
C48745 VPWR.n3720 VGND 0.01097f
C48746 VPWR.n3721 VGND 0.01144f
C48747 VPWR.n3722 VGND 0.01085f
C48748 VPWR.n3723 VGND 0.01085f
C48749 VPWR.n3724 VGND 0.01085f
C48750 VPWR.n3725 VGND 0.01085f
C48751 VPWR.n3726 VGND 0.01085f
C48752 VPWR.n3727 VGND 0.01085f
C48753 VPWR.n3728 VGND 0.00839f
C48754 VPWR.n3729 VGND 0.00985f
C48755 VPWR.n3730 VGND 0.01085f
C48756 VPWR.n3731 VGND 0.01085f
C48757 VPWR.n3732 VGND 0.01085f
C48758 VPWR.n3733 VGND 0.01085f
C48759 VPWR.n3734 VGND 0.01085f
C48760 VPWR.n3735 VGND 0.01085f
C48761 VPWR.n3736 VGND 0.0085f
C48762 VPWR.n3737 VGND 0.01077f
C48763 VPWR.n3738 VGND 0.00735f
C48764 VPWR.n3739 VGND 0.01189f
C48765 VPWR.n3740 VGND 0.01144f
C48766 VPWR.n3741 VGND 0.01085f
C48767 VPWR.n3742 VGND 0.01085f
C48768 VPWR.n3743 VGND 0.01085f
C48769 VPWR.n3744 VGND 0.01085f
C48770 VPWR.n3745 VGND 0.01085f
C48771 VPWR.n3746 VGND 0.00839f
C48772 VPWR.n3747 VGND 0.00985f
C48773 VPWR.n3748 VGND 0.01085f
C48774 VPWR.n3749 VGND 0.01085f
C48775 VPWR.n3750 VGND 0.01085f
C48776 VPWR.n3751 VGND 0.01085f
C48777 VPWR.n3752 VGND 0.00946f
C48778 VPWR.n3753 VGND 0.0083f
C48779 VPWR.n3754 VGND 0.10419f
C48780 VPWR.n3755 VGND 1.17131f
C48781 VPWR.n3756 VGND 0.01177f
C48782 VPWR.n3757 VGND 0.01163f
C48783 VPWR.n3758 VGND 0.01189f
C48784 VPWR.n3759 VGND 0.01839f
C48785 VPWR.n3760 VGND 0.0178f
C48786 VPWR.n3761 VGND 0.0178f
C48787 VPWR.n3762 VGND 0.01186f
C48788 VPWR.n3763 VGND 0.01679f
C48789 VPWR.n3764 VGND 0.0178f
C48790 VPWR.n3765 VGND 0.0178f
C48791 VPWR.n3766 VGND 0.01371f
C48792 VPWR.n3767 VGND 0.01189f
C48793 VPWR.n3768 VGND 0.01839f
C48794 VPWR.n3769 VGND 0.0178f
C48795 VPWR.n3770 VGND 0.0178f
C48796 VPWR.n3771 VGND 0.01186f
C48797 VPWR.n3772 VGND 0.01679f
C48798 VPWR.n3773 VGND 0.0178f
C48799 VPWR.n3774 VGND 0.01538f
C48800 VPWR.n3775 VGND 0.01177f
C48801 VPWR.n3776 VGND 0.78236f
C48802 VPWR.n3777 VGND 0.10419f
C48803 VPWR.n3778 VGND 0.01177f
C48804 VPWR.n3779 VGND 0.01309f
C48805 VPWR.n3780 VGND 0.01189f
C48806 VPWR.n3781 VGND 0.00889f
C48807 VPWR.n3782 VGND 0.00994f
C48808 VPWR.n3783 VGND 0.01085f
C48809 VPWR.n3784 VGND 0.01085f
C48810 VPWR.n3785 VGND 0.01085f
C48811 VPWR.n3786 VGND 0.01085f
C48812 VPWR.n3787 VGND 0.01085f
C48813 VPWR.n3788 VGND 0.00839f
C48814 VPWR.n3789 VGND 0.00985f
C48815 VPWR.n3790 VGND 0.01085f
C48816 VPWR.n3791 VGND 0.01085f
C48817 VPWR.n3792 VGND 0.01085f
C48818 VPWR.n3793 VGND 0.01085f
C48819 VPWR.n3794 VGND 0.01085f
C48820 VPWR.n3795 VGND 0.01085f
C48821 VPWR.n3796 VGND 0.01023f
C48822 VPWR.n3797 VGND 0.01189f
C48823 VPWR.n3798 VGND 0.00909f
C48824 VPWR.n3799 VGND 0.01303f
C48825 VPWR.n3800 VGND 0.01189f
C48826 VPWR.n3801 VGND 0.01144f
C48827 VPWR.n3802 VGND 0.01085f
C48828 VPWR.n3803 VGND 0.01085f
C48829 VPWR.n3804 VGND 0.01085f
C48830 VPWR.n3805 VGND 0.00839f
C48831 VPWR.n3806 VGND 0.00985f
C48832 VPWR.n3807 VGND 0.01085f
C48833 VPWR.n3808 VGND 0.01085f
C48834 VPWR.n3809 VGND 0.01085f
C48835 VPWR.n3810 VGND 0.01085f
C48836 VPWR.n3811 VGND 0.01085f
C48837 VPWR.n3812 VGND 0.01085f
C48838 VPWR.n3813 VGND 0.00741f
C48839 VPWR.n3814 VGND 0.00768f
C48840 VPWR.n3815 VGND 0.10419f
C48841 VPWR.n3816 VGND 0.78236f
C48842 VPWR.n3817 VGND 0.00768f
C48843 VPWR.n3818 VGND 0.01186f
C48844 VPWR.n3819 VGND 0.01839f
C48845 VPWR.n3820 VGND 0.0178f
C48846 VPWR.n3821 VGND 0.0178f
C48847 VPWR.n3822 VGND 0.01186f
C48848 VPWR.n3823 VGND 0.01679f
C48849 VPWR.n3824 VGND 0.0178f
C48850 VPWR.n3825 VGND 0.0178f
C48851 VPWR.n3826 VGND 0.01371f
C48852 VPWR.n3827 VGND 0.01189f
C48853 VPWR.n3828 VGND 0.01839f
C48854 VPWR.n3829 VGND 0.0178f
C48855 VPWR.n3830 VGND 0.0178f
C48856 VPWR.n3831 VGND 0.01186f
C48857 VPWR.n3832 VGND 0.01679f
C48858 VPWR.n3833 VGND 0.0178f
C48859 VPWR.n3834 VGND 0.0178f
C48860 VPWR.n3835 VGND 0.01333f
C48861 VPWR.n3836 VGND 0.00768f
C48862 VPWR.n3837 VGND 0.58789f
C48863 VPWR.n3838 VGND 0.10419f
C48864 VPWR.n3839 VGND 0.00768f
C48865 VPWR.n3840 VGND 0.00941f
.ends

