tt_um_algofoogle_vgaringosc_parax simulation

.include /home/anton/ttsetup@ttgf0p2/pdk/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/anton/ttsetup@ttgf0p2/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/anton/ttsetup@ttgf0p2/pdk/gf180mcuD/libs.tech/ngspice/smbb000149.ngspice typical
.include /home/anton/ttsetup@ttgf0p2/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/spice/gf180mcu_fd_sc_mcu7t5v0.spice

* This the SPICE netlist PEX (extraction from my design's GDS layout, including parasitics)
* which was generated with: make pex
* NOTE: That Make target assumes you have already generated the GDS using LibreLane,
* and that the source GDS therefore comes from runs/wokwi/final/gds/.
.include "tt_um_algofoogle_vgaringosc.from_gds.sim.spice"

* gf180mcuD uses 3.3V core logic:
.param vcc=3.3
vcc vcc 0 {vcc}

* Instantiate the tt_um_algofoogle_vgaringosc_parax DUT` (i.e. the circuit presenting my design)...
*NOTE: Port ordering matches how it was extracted by Magic:
xtt
+ 0
+ vcc
+ clk
+ ena
+ rst_n
+ ui_in[0]
+ ui_in[1]
+ ui_in[2]
+ ui_in[3]
+ ui_in[4]
+ ui_in[5]
+ ui_in[6]
+ ui_in[7]
+ uio_in[0]
+ uio_in[1]
+ uio_in[2]
+ uio_in[3]
+ uio_in[4]
+ uio_in[5]
+ uio_in[6]
+ uio_in[7]
+ uio_oe[0]
+ uio_oe[1]
+ uio_oe[2]
+ uio_oe[3]
+ uio_oe[4]
+ uio_oe[5]
+ uio_oe[6]
+ uio_oe[7]
+ uio_out[0]
+ uio_out[1]
+ uio_out[2]
+ uio_out[3]
+ uio_out[4]
+ uio_out[5]
+ uio_out[6]
+ uio_out[7]
+ uo_out[0]
+ uo_out[1]
+ uo_out[2]
+ uo_out[3]
+ uo_out[4]
+ uo_out[5]
+ uo_out[6]
+ uo_out[7]
+ tt_um_algofoogle_vgaringosc_parax

* Configure the inputs for this design...
VinEna    ena GND dc {vcc}
Vin0 ui_in[0] GND dc 0.0    ; clksel[0] ...Select a ring oscillator tapped at 'chain 10'...
Vin1 ui_in[1] GND dc {vcc}  ; clksel[1] ...
Vin2 ui_in[2] GND dc 0.0    ; clksel[2] ...
Vin3 ui_in[3] GND dc {vcc}  ; clksel[3] ...TAP10 ~= 75MHz?
Vin4 ui_in[4] GND dc 0.0    ; altclk ...not used unless clksel[3:0]==1
Vin5 ui_in[5] GND dc 0.0    ; mode[0] ...
Vin6 ui_in[6] GND dc 0.0    ; mode[1] ...(not used yet)
Vin7 ui_in[7] GND dc 0.0    ; vga_mode: 0=regular 640x480 59.94Hz

* Pulse generators...
*       net     ref fn     init   alt  dly  rise  fall  dut  period
* 25MHz system clock:
Vclk    clk     GND PULSE   0.0 {vcc}   0n    1n    1n  20n  40n
* reset signal (asserted for 80ns, starting 10ns into the simulation):
Vreset  rst_n   GND PULSE {vcc}   0.0  10n    1n    1n  80n  34m

*** Some options for speeding things up (at the cost of accuracy):
* * 1G-ohm shunt from all nodes to GND:
* .option rshunt = 1e9
* .options method=trap xmu=0.495
* .options reltol=2e-3 abstol=1e-11 vntol=1e-5 ; 0.2%, 10pA, 10uV -- Defaults: 1e-3 (0.1%), 1e-12 (1pA), 1e-6 (1uV).

.control
    save
    + vcc
    + i(vcc)
    + ena
    + clk
    + rst_n
    + "ui_in[0]"
    + "ui_in[1]"
    + "ui_in[2]"
    + "ui_in[3]"
    + "ui_in[4]"
    + "ui_in[5]"
    + "ui_in[6]"
    + "ui_in[7]"
    + "uio_in[0]"
    + "uio_in[1]"
    + "uio_in[2]"
    + "uio_in[3]"
    + "uio_in[4]"
    + "uio_in[5]"
    + "uio_in[6]"
    + "uio_in[7]"
    + "uio_oe[0]"
    + "uio_oe[1]"
    + "uio_oe[2]"
    + "uio_oe[3]"
    + "uio_oe[4]"
    + "uio_oe[5]"
    + "uio_oe[6]"
    + "uio_oe[7]"
    + "uio_out[0]"
    + "uio_out[1]"
    + "uio_out[2]"
    + "uio_out[3]"
    + "uio_out[4]"
    + "uio_out[5]"
    + "uio_out[6]"
    + "uio_out[7]"
    + "uo_out[0]"
    + "uo_out[1]"
    + "uo_out[2]"
    + "uo_out[3]"
    + "uo_out[4]"
    + "uo_out[5]"
    + "uo_out[6]"
    + "uo_out[7]"

    tran 8n 8193u 0 8n UIC ; 8192u is about 256 lines.

    * Write all the 'save' vectors (above) to a RAW file:
    write sim_out/full_spice_sim.raw

    * Save a snapshot of the simulation, so that hopefully we could resume it later:
    snsave sim_out/full_spice_sim.snap

    * Set up some colours for charting:
    set  color0=black           ; Background.
    set  color1=rgb:44/44/44    ; Text/grid.
    set  color2=rgb:77/00/77    ; (Dark magenta)
    set  color3=rgb:77/77/00    ; (Dark yellow)
    set  color4=rgb:ff/00/00    ; (Red)
    set  color5=rgb:00/ff/00    ; (Green)
    set  color6=rgb:00/00/ff    ; (Blue)
    set  color7=rgb:99/00/00    ; (Red, DARK)
    set  color8=rgb:00/99/00    ; (Green, DARK)
    set  color9=rgb:00/00/99    ; (Blue, DARK)
    set color10=rgb:cc/cc/00    ; (Mid yellow)
    set color11=rgb:cc/00/cc    ; (Mid magenta)

    * Plot the key signals w e care about:
    plot ena/4.4+0 clk/4.4+1 rst_n/4.4+2 "uio_out[4]"/4.4+3 "uio_out[5]"/4.4+4 "uio_out[6]"/4.4+5 "uio_out[7]"/4.4+6 "uo_out[7]"/4.4+7 "uo_out[3]"/4.4+8

.endc
.end
