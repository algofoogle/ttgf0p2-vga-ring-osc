`default_nettype none
//`timescale 1ns / 1ps

// See: https://gf180mcu-pdk.readthedocs.io/en/latest/digital/standard_cells/gf180mcu_fd_sc_mcu7t5v0/cells/inv/gf180mcu_fd_sc_mcu7t5v0__inv_1.html
`define PDK_INVERTER_CELL   gf180mcu_fd_sc_mcu7t5v0__inv_2
//NOTE: If you change this cell, the port names may need to be altered in any instances.

// This is to manage lint checking to not report about unconnected power pins.
// Thanks https://github.com/dlmiles/ttgf0p2-ringosc-5inv/blob/main/src/project.v
`ifdef USE_POWER_PINS
`define LINT_OFF_PINMISSING_POWER_PINS /* verilator lint_off PINMISSING */
`define LINT_ON_PINMISSING_POWER_PINS /* verilator lint_on PINMISSING */
`else
`define LINT_OFF_PINMISSING_POWER_PINS /* */
`define LINT_ON_PINMISSING_POWER_PINS /* */
`endif


module inverter_cell (
    input   wire a,
    output  wire y
);

    `LINT_OFF_PINMISSING_POWER_PINS
    (* keep_hierarchy *) `PDK_INVERTER_CELL pdkinv_notouch_ (
        .I  (a),
        .ZN (y)
    );
    `LINT_ON_PINMISSING_POWER_PINS

endmodule


// A chain of inverters (not a ring, itself)
module inv_chain #(
    parameter N = 10 // SHOULD BE EVEN.
) (
    input a,
    output y
);

    wire [N-1:0] ins;
    wire [N-1:0] outs;
    assign ins[0] = a;
    assign ins[N-1:1] = outs[N-2:0];
    assign y = outs[N-1];
    (* keep_hierarchy *) inverter_cell inv_array [N-1:0] ( .a(ins), .y(outs) );

endmodule


// A ring where the point of loopback is selectable:
module tapped_ring #(
    //NOTE: These parameters must be even-numbered since
    // there is a final baked-in inverter that makes the ring odd.
    //NOTE: These are deltas, i.e. each in turn is added to those before it.
    parameter TAP00 = 2,   // => 3      => 820
    parameter TAP01 = 2,   // => 5      => 492
    parameter TAP02 = 2,   // => 7      => 351
    parameter TAP03 = 2,   // => 9      => 273
    parameter TAP04 = 4,   // => 13     => 189
    parameter TAP05 = 4,   // => 17     => 145
    parameter TAP06 = 4,   // => 21     => 117
    parameter TAP07 = 4,   // => 25     => 98
    parameter TAP08 = 8,   // => 33     => 75
    parameter TAP09 = 8,   // => 41     => 60 MHz
    parameter TAP10 = 8,   // => 49     => 50
    parameter TAP11 = 16,  // => 65     => 38
    parameter TAP12 = 32,  // => 97     => ?
    parameter TAP13 = 64,  // => 161    => ?
    // Spares (not normally used by this design):
    parameter TAP14 = 2,   // => 163    => ?
    parameter TAP15 = 2    // => 165    => ?
) (
    input ena,
    input [3:0] tap,
    output y
);
    wire ring_head;
    wire [15:0] chain;

    assign y = ena && chain[tap];

    (* keep_hierarchy *) inverter_cell         head ( .a(y),         .y(ring_head) ); // If all the counts below are even, this makes it odd.
    (* keep_hierarchy *) inv_chain #(.N(TAP00)) c00 ( .a(ring_head), .y(chain[ 0]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP01)) c01 ( .a(chain[ 0]), .y(chain[ 1]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP02)) c02 ( .a(chain[ 1]), .y(chain[ 2]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP03)) c03 ( .a(chain[ 2]), .y(chain[ 3]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP04)) c04 ( .a(chain[ 3]), .y(chain[ 4]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP05)) c05 ( .a(chain[ 4]), .y(chain[ 5]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP06)) c06 ( .a(chain[ 5]), .y(chain[ 6]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP07)) c07 ( .a(chain[ 6]), .y(chain[ 7]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP08)) c08 ( .a(chain[ 7]), .y(chain[ 8]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP09)) c09 ( .a(chain[ 8]), .y(chain[ 9]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP10)) c10 ( .a(chain[ 9]), .y(chain[10]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP11)) c11 ( .a(chain[10]), .y(chain[11]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP12)) c12 ( .a(chain[11]), .y(chain[12]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP13)) c13 ( .a(chain[12]), .y(chain[13]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP14)) c14 ( .a(chain[13]), .y(chain[14]) );
    (* keep_hierarchy *) inv_chain #(.N(TAP15)) c15 ( .a(chain[14]), .y(chain[15]) );
endmodule

// Just a short, fixed ring: by default, 5 instances of inv_1:
module ringosc_inv1 #(
    parameter N = 5 // Must be odd-numbered!
) (
    input ena,
    output y
);
    wire [N-1:0] ins;
    wire [N-1:0] outs;
    assign ins[N-1:1] = outs[N-2:0];
    assign ins[0] = outs[N-1] & ena; // ena==0 will break the loop (stop the oscillator ring, hence flush it out too).
    assign y = ins[0];
    (* keep_hierarchy *) gf180mcu_fd_sc_mcu7t5v0__inv_1 inv_array_notouch_ [N-1:0] (.I(ins), .ZN(outs));
endmodule

// Another short, fixed ring: by default, 5 instances of inv_4:
module ringosc_inv4 #(
    parameter N = 5 // Must be odd-numbered!
) (
    input ena,
    output y
);
    wire [N-1:0] ins;
    wire [N-1:0] outs;
    assign ins[N-1:1] = outs[N-2:0];
    assign ins[0] = outs[N-1] & ena; // ena==0 will break the loop (stop the oscillator ring, hence flush it out too).
    assign y = ins[0];
    (* keep_hierarchy *) gf180mcu_fd_sc_mcu7t5v0__inv_4 inv_array_notouch_ [N-1:0] (.I(ins), .ZN(outs));
endmodule
